magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 4790 1094
<< pwell >>
rect -86 -86 4790 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 716 215 836 333
rect 940 215 1060 333
rect 1164 215 1284 333
rect 1353 215 1473 333
rect 1577 215 1697 333
rect 1761 215 1881 333
rect 1993 215 2113 333
rect 2217 215 2337 333
rect 2849 215 2969 333
rect 3017 215 3137 333
rect 3285 69 3405 333
rect 3509 69 3629 333
rect 3733 69 3853 333
rect 3957 69 4077 333
rect 4181 69 4301 333
rect 4405 69 4525 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 736 593 836 793
rect 989 593 1089 793
rect 1193 593 1293 793
rect 1373 593 1473 793
rect 1577 593 1677 793
rect 1781 593 1881 793
rect 2217 573 2317 773
rect 2485 573 2585 773
rect 2833 573 2933 773
rect 3037 573 3137 773
rect 3285 573 3385 939
rect 3489 573 3589 939
rect 3693 573 3793 939
rect 3897 573 3997 939
rect 4101 573 4201 939
rect 4305 573 4405 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 468 274 497 320
rect 543 274 556 320
rect 468 175 556 274
rect 628 274 716 333
rect 628 228 641 274
rect 687 228 716 274
rect 628 215 716 228
rect 836 320 940 333
rect 836 274 865 320
rect 911 274 940 320
rect 836 215 940 274
rect 1060 320 1164 333
rect 1060 274 1089 320
rect 1135 274 1164 320
rect 1060 215 1164 274
rect 1284 215 1353 333
rect 1473 274 1577 333
rect 1473 228 1502 274
rect 1548 228 1577 274
rect 1473 215 1577 228
rect 1697 215 1761 333
rect 1881 320 1993 333
rect 1881 274 1910 320
rect 1956 274 1993 320
rect 1881 215 1993 274
rect 2113 274 2217 333
rect 2113 228 2142 274
rect 2188 228 2217 274
rect 2113 215 2217 228
rect 2337 320 2425 333
rect 2337 274 2366 320
rect 2412 274 2425 320
rect 2337 215 2425 274
rect 2761 320 2849 333
rect 2761 274 2774 320
rect 2820 274 2849 320
rect 2761 215 2849 274
rect 2969 215 3017 333
rect 3137 215 3285 333
rect 3197 128 3285 215
rect 3197 82 3210 128
rect 3256 82 3285 128
rect 3197 69 3285 82
rect 3405 320 3509 333
rect 3405 180 3434 320
rect 3480 180 3509 320
rect 3405 69 3509 180
rect 3629 222 3733 333
rect 3629 82 3658 222
rect 3704 82 3733 222
rect 3629 69 3733 82
rect 3853 320 3957 333
rect 3853 180 3882 320
rect 3928 180 3957 320
rect 3853 69 3957 180
rect 4077 222 4181 333
rect 4077 82 4106 222
rect 4152 82 4181 222
rect 4077 69 4181 82
rect 4301 320 4405 333
rect 4301 180 4330 320
rect 4376 180 4405 320
rect 4301 69 4405 180
rect 4525 222 4613 333
rect 4525 82 4554 222
rect 4600 82 4613 222
rect 4525 69 4613 82
<< mvpdiff >>
rect 56 739 144 849
rect 56 599 69 739
rect 115 599 144 739
rect 56 573 144 599
rect 244 836 348 849
rect 244 696 273 836
rect 319 696 348 836
rect 244 573 348 696
rect 448 726 536 849
rect 1941 823 2013 836
rect 1941 793 1954 823
rect 448 586 477 726
rect 523 586 536 726
rect 648 780 736 793
rect 648 734 661 780
rect 707 734 736 780
rect 648 593 736 734
rect 836 746 989 793
rect 836 606 865 746
rect 911 606 989 746
rect 836 593 989 606
rect 1089 746 1193 793
rect 1089 606 1118 746
rect 1164 606 1193 746
rect 1089 593 1193 606
rect 1293 593 1373 793
rect 1473 780 1577 793
rect 1473 734 1502 780
rect 1548 734 1577 780
rect 1473 593 1577 734
rect 1677 652 1781 793
rect 1677 606 1706 652
rect 1752 606 1781 652
rect 1677 593 1781 606
rect 1881 777 1954 793
rect 2000 777 2013 823
rect 1881 593 2013 777
rect 3205 773 3285 939
rect 2129 632 2217 773
rect 448 573 536 586
rect 2129 586 2142 632
rect 2188 586 2217 632
rect 2129 573 2217 586
rect 2317 726 2485 773
rect 2317 586 2346 726
rect 2392 586 2485 726
rect 2317 573 2485 586
rect 2585 632 2673 773
rect 2585 586 2614 632
rect 2660 586 2673 632
rect 2585 573 2673 586
rect 2745 760 2833 773
rect 2745 714 2758 760
rect 2804 714 2833 760
rect 2745 573 2833 714
rect 2933 726 3037 773
rect 2933 586 2962 726
rect 3008 586 3037 726
rect 2933 573 3037 586
rect 3137 760 3285 773
rect 3137 620 3166 760
rect 3212 620 3285 760
rect 3137 573 3285 620
rect 3385 726 3489 939
rect 3385 586 3414 726
rect 3460 586 3489 726
rect 3385 573 3489 586
rect 3589 926 3693 939
rect 3589 786 3618 926
rect 3664 786 3693 926
rect 3589 573 3693 786
rect 3793 726 3897 939
rect 3793 586 3822 726
rect 3868 586 3897 726
rect 3793 573 3897 586
rect 3997 926 4101 939
rect 3997 786 4026 926
rect 4072 786 4101 926
rect 3997 573 4101 786
rect 4201 726 4305 939
rect 4201 586 4230 726
rect 4276 586 4305 726
rect 4201 573 4305 586
rect 4405 926 4493 939
rect 4405 786 4434 926
rect 4480 786 4493 926
rect 4405 573 4493 786
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 641 228 687 274
rect 865 274 911 320
rect 1089 274 1135 320
rect 1502 228 1548 274
rect 1910 274 1956 320
rect 2142 228 2188 274
rect 2366 274 2412 320
rect 2774 274 2820 320
rect 3210 82 3256 128
rect 3434 180 3480 320
rect 3658 82 3704 222
rect 3882 180 3928 320
rect 4106 82 4152 222
rect 4330 180 4376 320
rect 4554 82 4600 222
<< mvpdiffc >>
rect 69 599 115 739
rect 273 696 319 836
rect 477 586 523 726
rect 661 734 707 780
rect 865 606 911 746
rect 1118 606 1164 746
rect 1502 734 1548 780
rect 1706 606 1752 652
rect 1954 777 2000 823
rect 2142 586 2188 632
rect 2346 586 2392 726
rect 2614 586 2660 632
rect 2758 714 2804 760
rect 2962 586 3008 726
rect 3166 620 3212 760
rect 3414 586 3460 726
rect 3618 786 3664 926
rect 3822 586 3868 726
rect 4026 786 4072 926
rect 4230 586 4276 726
rect 4434 786 4480 926
<< polysilicon >>
rect 348 933 1293 973
rect 144 849 244 893
rect 348 849 448 933
rect 989 872 1089 885
rect 736 793 836 837
rect 989 826 1002 872
rect 1048 826 1089 872
rect 989 793 1089 826
rect 1193 872 1293 933
rect 1193 826 1234 872
rect 1280 826 1293 872
rect 1781 913 2933 953
rect 3285 939 3385 983
rect 3489 939 3589 983
rect 3693 939 3793 983
rect 3897 939 3997 983
rect 4101 939 4201 983
rect 4305 939 4405 983
rect 1193 793 1293 826
rect 1373 793 1473 837
rect 1577 793 1677 837
rect 1781 793 1881 913
rect 2217 852 2317 865
rect 2217 806 2230 852
rect 2276 806 2317 852
rect 2217 773 2317 806
rect 2485 773 2585 817
rect 2833 773 2933 913
rect 3037 773 3137 817
rect 144 494 244 573
rect 144 448 157 494
rect 203 448 244 494
rect 144 377 244 448
rect 124 333 244 377
rect 348 425 448 573
rect 348 379 372 425
rect 418 379 448 425
rect 348 377 448 379
rect 736 512 836 593
rect 736 466 749 512
rect 795 466 836 512
rect 989 533 1089 593
rect 1193 549 1293 593
rect 1373 560 1473 593
rect 989 493 1147 533
rect 736 377 836 466
rect 1107 433 1147 493
rect 1373 514 1414 560
rect 1460 514 1473 560
rect 1107 412 1284 433
rect 1107 393 1211 412
rect 348 333 468 377
rect 716 333 836 377
rect 940 333 1060 377
rect 1164 366 1211 393
rect 1257 366 1284 412
rect 1373 377 1473 514
rect 1164 333 1284 366
rect 1353 333 1473 377
rect 1577 468 1677 593
rect 1577 422 1590 468
rect 1636 422 1677 468
rect 1577 377 1677 422
rect 1781 377 1881 593
rect 2217 377 2317 573
rect 1577 333 1697 377
rect 1761 333 1881 377
rect 1993 333 2113 377
rect 2217 333 2337 377
rect 124 131 244 175
rect 348 115 468 175
rect 716 171 836 215
rect 940 115 1060 215
rect 1164 171 1284 215
rect 1353 171 1473 215
rect 1577 171 1697 215
rect 1761 171 1881 215
rect 1993 182 2113 215
rect 348 75 1060 115
rect 1993 136 2006 182
rect 2052 136 2113 182
rect 2217 171 2337 215
rect 1993 123 2113 136
rect 2485 123 2585 573
rect 2833 490 2933 573
rect 2833 444 2846 490
rect 2892 444 2933 490
rect 2833 393 2933 444
rect 3037 493 3137 573
rect 3037 447 3050 493
rect 3096 447 3137 493
rect 2849 333 2969 393
rect 3037 377 3137 447
rect 3017 333 3137 377
rect 3285 433 3385 573
rect 3489 433 3589 573
rect 3693 529 3793 573
rect 3285 412 3589 433
rect 3285 366 3298 412
rect 3344 393 3589 412
rect 3344 366 3405 393
rect 3285 333 3405 366
rect 3509 377 3589 393
rect 3733 465 3793 529
rect 3897 465 3997 573
rect 4101 465 4201 573
rect 4305 465 4405 573
rect 3733 452 4525 465
rect 3733 406 3746 452
rect 3792 406 3926 452
rect 3972 406 4127 452
rect 4173 406 4525 452
rect 3733 393 4525 406
rect 3509 333 3629 377
rect 3733 333 3853 393
rect 3957 333 4077 393
rect 4181 333 4301 393
rect 4405 333 4525 393
rect 2849 171 2969 215
rect 3017 171 3137 215
rect 1993 83 2585 123
rect 3285 25 3405 69
rect 3509 25 3629 69
rect 3733 25 3853 69
rect 3957 25 4077 69
rect 4181 25 4301 69
rect 4405 25 4525 69
<< polycontact >>
rect 1002 826 1048 872
rect 1234 826 1280 872
rect 2230 806 2276 852
rect 157 448 203 494
rect 372 379 418 425
rect 749 466 795 512
rect 1414 514 1460 560
rect 1211 366 1257 412
rect 1590 422 1636 468
rect 2006 136 2052 182
rect 2846 444 2892 490
rect 3050 447 3096 493
rect 3298 366 3344 412
rect 3746 406 3792 452
rect 3926 406 3972 452
rect 4127 406 4173 452
<< metal1 >>
rect 0 926 4704 1098
rect 0 918 3618 926
rect 273 836 319 918
rect 69 739 115 750
rect 661 780 707 918
rect 273 685 319 696
rect 477 726 523 737
rect 115 599 418 634
rect 69 588 418 599
rect 142 494 314 542
rect 142 448 157 494
rect 203 448 314 494
rect 372 425 418 588
rect 372 337 418 379
rect 49 320 418 337
rect 95 291 418 320
rect 661 723 707 734
rect 753 826 1002 872
rect 1048 826 1059 872
rect 1223 826 1234 872
rect 1280 826 1291 872
rect 753 677 799 826
rect 523 631 799 677
rect 865 746 911 757
rect 523 586 543 631
rect 477 320 543 586
rect 589 512 806 542
rect 589 466 749 512
rect 795 466 806 512
rect 49 263 95 274
rect 477 274 497 320
rect 865 320 911 606
rect 477 263 543 274
rect 641 274 687 285
rect 273 234 319 245
rect 273 90 319 188
rect 865 263 911 274
rect 1089 746 1164 757
rect 1089 606 1118 746
rect 1223 677 1291 826
rect 1502 780 1548 918
rect 1943 823 2011 918
rect 1943 777 1954 823
rect 2000 777 2011 823
rect 2230 852 2276 863
rect 1502 723 1548 734
rect 1594 731 1909 744
rect 2230 731 2276 806
rect 2758 760 2804 918
rect 1594 698 2276 731
rect 1594 677 1640 698
rect 1864 685 2276 698
rect 2346 726 2392 737
rect 1223 631 1640 677
rect 1089 504 1164 606
rect 1695 606 1706 652
rect 1752 606 1763 652
rect 1695 560 1763 606
rect 2131 586 2142 632
rect 2188 586 2199 632
rect 2131 560 2199 586
rect 1403 514 1414 560
rect 1460 514 2199 560
rect 3166 760 3212 918
rect 3664 918 4026 926
rect 3618 775 3664 786
rect 4072 918 4434 926
rect 4026 775 4072 786
rect 4480 918 4704 926
rect 4434 775 4480 786
rect 2758 703 2804 714
rect 2962 726 3008 737
rect 1089 468 1358 504
rect 1089 458 1590 468
rect 1089 320 1135 458
rect 1313 422 1590 458
rect 1636 422 1647 468
rect 1200 366 1211 412
rect 1257 376 1268 412
rect 1257 366 1864 376
rect 1200 330 1864 366
rect 1089 263 1135 274
rect 641 90 687 228
rect 1491 228 1502 274
rect 1548 228 1559 274
rect 1491 90 1559 228
rect 1818 182 1864 330
rect 1910 320 1956 514
rect 2346 423 2392 586
rect 2274 377 2392 423
rect 2614 632 2962 643
rect 2660 597 2962 632
rect 2274 285 2320 377
rect 2614 331 2660 586
rect 3166 609 3212 620
rect 3414 726 3461 737
rect 2962 575 3008 586
rect 3460 586 3461 726
rect 2706 490 2903 542
rect 3414 504 3461 586
rect 3822 726 3868 737
rect 4230 726 4376 737
rect 3868 586 4230 621
rect 4276 586 4376 726
rect 3822 575 4376 586
rect 2706 444 2846 490
rect 2892 444 2903 490
rect 3050 493 3461 504
rect 3096 465 3461 493
rect 3096 458 4184 465
rect 3050 436 3096 447
rect 3415 452 4184 458
rect 3136 366 3298 412
rect 3344 366 3355 412
rect 3415 406 3746 452
rect 3792 406 3926 452
rect 3972 406 4127 452
rect 4173 406 4184 452
rect 1910 263 1956 274
rect 2142 274 2320 285
rect 2188 228 2320 274
rect 2366 320 2820 331
rect 2412 274 2774 320
rect 2366 263 2820 274
rect 2142 217 2320 228
rect 3136 217 3182 366
rect 1818 136 2006 182
rect 2052 136 2063 182
rect 2142 171 3182 217
rect 3415 320 3480 406
rect 4318 331 4376 575
rect 3415 180 3434 320
rect 3881 320 4376 331
rect 3415 169 3480 180
rect 3658 222 3704 233
rect 3199 90 3210 128
rect 0 82 3210 90
rect 3256 90 3267 128
rect 3256 82 3658 90
rect 3881 180 3882 320
rect 3928 279 4330 320
rect 3881 169 3928 180
rect 4106 222 4152 233
rect 3704 82 4106 90
rect 4318 180 4330 279
rect 4318 169 4376 180
rect 4554 222 4600 233
rect 4152 82 4554 90
rect 4600 82 4704 90
rect 0 -90 4704 82
<< labels >>
flabel metal1 s 142 448 314 542 0 FreeSans 200 0 0 0 CLK
port 3 nsew clock input
flabel metal1 s 589 466 806 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4230 621 4376 737 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2706 444 2903 542 0 FreeSans 200 0 0 0 SETN
port 2 nsew default input
flabel metal1 s 0 918 4704 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 641 274 687 285 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 3822 621 3868 737 1 Q
port 4 nsew default output
rlabel metal1 s 3822 575 4376 621 1 Q
port 4 nsew default output
rlabel metal1 s 4318 331 4376 575 1 Q
port 4 nsew default output
rlabel metal1 s 3881 279 4376 331 1 Q
port 4 nsew default output
rlabel metal1 s 4318 169 4376 279 1 Q
port 4 nsew default output
rlabel metal1 s 3881 169 3928 279 1 Q
port 4 nsew default output
rlabel metal1 s 4434 777 4480 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4026 777 4072 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3618 777 3664 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3166 777 3212 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2758 777 2804 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1943 777 2011 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1502 777 1548 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 777 707 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 777 319 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4434 775 4480 777 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 4026 775 4072 777 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3618 775 3664 777 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3166 775 3212 777 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2758 775 2804 777 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1502 775 1548 777 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 775 707 777 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 775 319 777 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3166 723 3212 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2758 723 2804 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1502 723 1548 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 661 723 707 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 723 319 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3166 703 3212 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2758 703 2804 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 703 319 723 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3166 685 3212 703 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 273 685 319 703 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3166 609 3212 685 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1491 245 1559 274 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 641 245 687 274 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1491 233 1559 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 641 233 687 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4554 128 4600 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4106 128 4152 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3658 128 3704 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1491 128 1559 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 641 128 687 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 128 319 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4554 90 4600 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4106 90 4152 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3658 90 3704 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3199 90 3267 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1491 90 1559 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 128 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4704 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4704 1008
string GDS_END 693442
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 683132
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
