magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 770 1486
<< nmos >>
rect 120 209 176 385
rect 324 209 380 452
<< pmos >>
rect 120 1015 176 1191
rect 324 908 380 1191
<< ndiff >>
rect 236 385 324 452
rect 32 371 120 385
rect 32 325 45 371
rect 91 325 120 371
rect 32 209 120 325
rect 176 268 324 385
rect 176 222 249 268
rect 295 222 324 268
rect 176 209 324 222
rect 380 405 468 452
rect 380 359 409 405
rect 455 359 468 405
rect 380 209 468 359
<< pdiff >>
rect 32 1075 120 1191
rect 32 1029 45 1075
rect 91 1029 120 1075
rect 32 1015 120 1029
rect 176 1178 324 1191
rect 176 1132 249 1178
rect 295 1132 324 1178
rect 176 1015 324 1132
rect 236 908 324 1015
rect 380 1071 468 1191
rect 380 925 409 1071
rect 455 925 468 1071
rect 380 908 468 925
<< ndiffc >>
rect 45 325 91 371
rect 249 222 295 268
rect 409 359 455 405
<< pdiffc >>
rect 45 1029 91 1075
rect 249 1132 295 1178
rect 409 925 455 1071
<< psubdiff >>
rect 28 87 656 100
rect 28 41 69 87
rect 615 41 656 87
rect 28 28 656 41
<< nsubdiff >>
rect 28 1359 656 1372
rect 28 1313 69 1359
rect 615 1313 656 1359
rect 28 1300 656 1313
<< psubdiffcont >>
rect 69 41 615 87
<< nsubdiffcont >>
rect 69 1313 615 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 324 1191 380 1235
rect 120 848 176 1015
rect 120 835 202 848
rect 120 789 143 835
rect 189 789 202 835
rect 120 776 202 789
rect 324 716 380 908
rect 32 703 380 716
rect 32 657 45 703
rect 91 657 380 703
rect 32 644 380 657
rect 120 571 202 584
rect 120 525 143 571
rect 189 525 202 571
rect 120 512 202 525
rect 120 385 176 512
rect 324 452 380 644
rect 120 165 176 209
rect 324 165 380 209
<< polycontact >>
rect 143 789 189 835
rect 45 657 91 703
rect 143 525 189 571
<< metal1 >>
rect 0 1359 684 1400
rect 0 1313 69 1359
rect 615 1313 684 1359
rect 0 1178 684 1313
rect 0 1132 249 1178
rect 295 1132 684 1178
rect 42 1075 94 1086
rect 42 1029 45 1075
rect 91 1029 94 1075
rect 42 703 94 1029
rect 42 657 45 703
rect 91 657 94 703
rect 42 371 94 657
rect 42 325 45 371
rect 91 325 94 371
rect 42 314 94 325
rect 140 835 192 1086
rect 140 789 143 835
rect 189 789 192 835
rect 140 571 192 789
rect 140 525 143 571
rect 189 525 192 571
rect 140 314 192 525
rect 406 1071 458 1086
rect 406 925 409 1071
rect 455 925 458 1071
rect 406 405 458 925
rect 406 359 409 405
rect 455 359 458 405
rect 406 314 458 359
rect 0 222 249 268
rect 295 222 684 268
rect 0 87 684 222
rect 0 41 69 87
rect 615 41 684 87
rect 0 0 684 41
<< labels >>
rlabel metal1 s 0 1132 684 1400 4 vdd
port 3 nsew
rlabel metal1 s 0 0 684 268 4 vss
port 5 nsew
rlabel metal1 s 140 314 192 1086 4 i
port 7 nsew
rlabel metal1 s 406 314 458 1086 4 q
port 9 nsew
<< end >>
