magic
tech gf180mcuD
magscale 1 10
timestamp 1751558652
<< nwell >>
rect -86 354 1094 870
<< pwell >>
rect -86 -86 1094 354
<< nmos >>
rect 116 68 172 212
rect 276 68 332 212
rect 436 68 492 212
rect 596 68 652 212
rect 756 68 812 212
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
<< ndiff >>
rect 28 163 116 212
rect 28 117 41 163
rect 87 117 116 163
rect 28 68 116 117
rect 172 127 276 212
rect 172 81 201 127
rect 247 81 276 127
rect 172 68 276 81
rect 332 163 436 212
rect 332 117 361 163
rect 407 117 436 163
rect 332 68 436 117
rect 492 127 596 212
rect 492 81 521 127
rect 567 81 596 127
rect 492 68 596 81
rect 652 163 756 212
rect 652 117 681 163
rect 727 117 756 163
rect 652 68 756 117
rect 812 127 980 212
rect 812 81 841 127
rect 887 81 980 127
rect 812 68 980 81
<< pdiff >>
rect 28 655 116 716
rect 28 573 41 655
rect 87 573 116 655
rect 28 440 116 573
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 667 436 716
rect 332 453 361 667
rect 407 453 436 667
rect 332 440 436 453
rect 492 703 596 716
rect 492 657 521 703
rect 567 657 596 703
rect 492 440 596 657
rect 652 667 756 716
rect 652 453 681 667
rect 727 453 756 667
rect 652 440 756 453
rect 812 703 980 716
rect 812 453 841 703
rect 887 453 980 703
rect 812 440 980 453
<< ndiffc >>
rect 41 117 87 163
rect 201 81 247 127
rect 361 117 407 163
rect 521 81 567 127
rect 681 117 727 163
rect 841 81 887 127
<< pdiffc >>
rect 41 573 87 655
rect 201 657 247 703
rect 361 453 407 667
rect 521 657 567 703
rect 681 453 727 667
rect 841 453 887 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 116 405 172 440
rect 276 406 332 440
rect 74 382 172 405
rect 74 336 89 382
rect 135 336 172 382
rect 74 314 172 336
rect 220 394 332 406
rect 436 401 492 440
rect 596 401 652 440
rect 756 401 812 440
rect 436 394 812 401
rect 220 385 812 394
rect 220 339 233 385
rect 279 347 812 385
rect 279 339 492 347
rect 220 338 492 339
rect 220 315 332 338
rect 116 212 172 314
rect 276 212 332 315
rect 436 212 492 338
rect 596 212 652 347
rect 756 212 812 347
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
<< polycontact >>
rect 89 336 135 382
rect 233 339 279 385
<< metal1 >>
rect 0 724 1008 844
rect 201 703 247 724
rect 41 655 87 676
rect 521 703 567 724
rect 201 646 247 657
rect 361 667 440 678
rect 87 573 266 579
rect 41 533 266 573
rect 41 382 135 457
rect 41 336 89 382
rect 41 314 135 336
rect 220 406 266 533
rect 407 453 440 667
rect 841 703 887 724
rect 521 646 567 657
rect 681 667 760 678
rect 361 408 440 453
rect 727 453 760 667
rect 681 408 760 453
rect 841 428 887 453
rect 220 385 279 406
rect 220 339 233 385
rect 220 315 279 339
rect 361 351 760 408
rect 220 235 266 315
rect 41 189 266 235
rect 41 163 87 189
rect 361 163 440 351
rect 41 106 87 117
rect 201 127 247 138
rect 407 117 440 163
rect 681 163 760 351
rect 361 106 440 117
rect 521 127 567 138
rect 201 60 247 81
rect 727 117 760 163
rect 681 106 760 117
rect 841 127 887 146
rect 521 60 567 81
rect 841 60 887 81
rect 0 -60 1008 60
<< labels >>
flabel metal1 s 0 724 1008 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1008 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 41 314 135 457 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 681 106 760 678 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
flabel metal1 361 106 440 678 0 FreeSans 200 0 0 0 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1008 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
