magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 1226 1486
<< nmos >>
rect 120 209 176 385
rect 280 209 336 385
rect 440 209 496 385
rect 600 209 656 385
rect 760 209 816 385
rect 964 209 1020 452
<< pmos >>
rect 120 1015 176 1191
rect 280 1015 336 1191
rect 440 1015 496 1191
rect 600 1015 656 1191
rect 760 1015 816 1191
rect 964 908 1020 1191
<< ndiff >>
rect 876 385 964 452
rect 32 371 120 385
rect 32 325 45 371
rect 91 325 120 371
rect 32 209 120 325
rect 176 268 280 385
rect 176 222 205 268
rect 251 222 280 268
rect 176 209 280 222
rect 336 209 440 385
rect 496 371 600 385
rect 496 325 525 371
rect 571 325 600 371
rect 496 209 600 325
rect 656 209 760 385
rect 816 268 964 385
rect 816 222 889 268
rect 935 222 964 268
rect 816 209 964 222
rect 1020 405 1108 452
rect 1020 359 1049 405
rect 1095 359 1108 405
rect 1020 209 1108 359
<< pdiff >>
rect 32 1075 120 1191
rect 32 1029 45 1075
rect 91 1029 120 1075
rect 32 1015 120 1029
rect 176 1178 280 1191
rect 176 1132 205 1178
rect 251 1132 280 1178
rect 176 1015 280 1132
rect 336 1015 440 1191
rect 496 1075 600 1191
rect 496 1029 525 1075
rect 571 1029 600 1075
rect 496 1015 600 1029
rect 656 1015 760 1191
rect 816 1178 964 1191
rect 816 1132 889 1178
rect 935 1132 964 1178
rect 816 1015 964 1132
rect 876 908 964 1015
rect 1020 1071 1108 1191
rect 1020 925 1049 1071
rect 1095 925 1108 1071
rect 1020 908 1108 925
<< ndiffc >>
rect 45 325 91 371
rect 205 222 251 268
rect 525 325 571 371
rect 889 222 935 268
rect 1049 359 1095 405
<< pdiffc >>
rect 45 1029 91 1075
rect 205 1132 251 1178
rect 525 1029 571 1075
rect 889 1132 935 1178
rect 1049 925 1095 1071
<< psubdiff >>
rect 28 87 1112 100
rect 28 41 47 87
rect 1093 41 1112 87
rect 28 28 1112 41
<< nsubdiff >>
rect 28 1359 1112 1372
rect 28 1313 47 1359
rect 1093 1313 1112 1359
rect 28 1300 1112 1313
<< psubdiffcont >>
rect 47 41 1093 87
<< nsubdiffcont >>
rect 47 1313 1093 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 600 1191 656 1235
rect 760 1191 816 1235
rect 964 1191 1020 1235
rect 120 716 176 1015
rect 280 848 336 1015
rect 228 835 336 848
rect 228 789 241 835
rect 287 789 336 835
rect 228 776 336 789
rect 440 716 496 1015
rect 600 848 656 1015
rect 544 835 656 848
rect 544 789 557 835
rect 603 789 656 835
rect 544 776 656 789
rect 120 703 656 716
rect 120 657 143 703
rect 189 657 656 703
rect 120 644 656 657
rect 120 385 176 644
rect 228 571 336 584
rect 228 525 241 571
rect 287 525 336 571
rect 228 512 336 525
rect 384 571 496 584
rect 384 525 397 571
rect 443 525 496 571
rect 384 512 496 525
rect 280 385 336 512
rect 440 385 496 512
rect 600 385 656 644
rect 760 584 816 1015
rect 964 716 1020 908
rect 864 703 1020 716
rect 864 657 877 703
rect 923 657 1020 703
rect 864 644 1020 657
rect 704 571 816 584
rect 704 525 717 571
rect 763 525 816 571
rect 704 512 816 525
rect 760 385 816 512
rect 964 452 1020 644
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
rect 600 165 656 209
rect 760 165 816 209
rect 964 165 1020 209
<< polycontact >>
rect 241 789 287 835
rect 557 789 603 835
rect 143 657 189 703
rect 241 525 287 571
rect 397 525 443 571
rect 877 657 923 703
rect 717 525 763 571
<< metal1 >>
rect 0 1359 1140 1400
rect 0 1313 47 1359
rect 1093 1313 1140 1359
rect 0 1178 1140 1313
rect 0 1132 205 1178
rect 251 1132 889 1178
rect 935 1132 1140 1178
rect 42 1075 94 1086
rect 42 1029 45 1075
rect 91 1029 94 1075
rect 42 382 94 1029
rect 140 703 192 1086
rect 140 657 143 703
rect 189 657 192 703
rect 140 428 192 657
rect 238 835 290 1086
rect 525 1075 926 1086
rect 571 1029 926 1075
rect 525 1018 926 1029
rect 238 789 241 835
rect 287 789 290 835
rect 238 571 290 789
rect 238 525 241 571
rect 287 525 290 571
rect 238 428 290 525
rect 394 835 603 846
rect 394 789 557 835
rect 394 778 603 789
rect 394 571 446 778
rect 394 525 397 571
rect 443 525 446 571
rect 394 382 446 525
rect 714 571 766 972
rect 714 525 717 571
rect 763 525 766 571
rect 714 428 766 525
rect 874 703 926 1018
rect 874 657 877 703
rect 923 657 926 703
rect 874 382 926 657
rect 42 371 446 382
rect 42 325 45 371
rect 91 325 446 371
rect 42 314 446 325
rect 525 371 926 382
rect 571 325 926 371
rect 525 314 926 325
rect 1046 1071 1098 1086
rect 1046 925 1049 1071
rect 1095 925 1098 1071
rect 1046 405 1098 925
rect 1046 359 1049 405
rect 1095 359 1098 405
rect 1046 314 1098 359
rect 0 222 205 268
rect 251 222 889 268
rect 935 222 1140 268
rect 0 87 1140 222
rect 0 41 47 87
rect 1093 41 1140 87
rect 0 0 1140 41
<< labels >>
rlabel metal1 s 0 1132 1140 1400 4 vdd
port 3 nsew
rlabel metal1 s 0 0 1140 268 4 vss
port 5 nsew
rlabel metal1 s 140 428 192 1086 4 cmd
port 7 nsew
rlabel metal1 s 238 428 290 1086 4 i0
port 9 nsew
rlabel metal1 s 714 428 766 972 4 i1
port 11 nsew
rlabel metal1 s 1046 314 1098 1086 4 q
port 13 nsew
<< end >>
