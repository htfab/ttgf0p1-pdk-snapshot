magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 352 1318 870
<< pwell >>
rect -86 -86 1318 352
<< metal1 >>
rect 0 724 1232 844
rect 273 632 319 724
rect 24 354 214 430
rect 136 232 214 354
rect 350 356 538 430
rect 350 242 430 356
rect 584 310 648 664
rect 801 317 874 567
rect 920 241 984 573
rect 590 195 984 241
rect 1030 232 1102 460
rect 590 181 636 195
rect 38 60 106 163
rect 430 135 636 181
rect 920 181 984 195
rect 734 60 802 149
rect 920 135 1196 181
rect 0 -60 1232 60
<< obsm1 >>
rect 56 586 126 676
rect 466 586 534 676
rect 56 518 534 586
rect 709 630 1183 676
rect 709 506 755 630
rect 1137 506 1183 630
<< labels >>
rlabel metal1 s 1030 232 1102 460 6 A1
port 1 nsew default input
rlabel metal1 s 801 317 874 567 6 A2
port 2 nsew default input
rlabel metal1 s 350 242 430 356 6 B1
port 3 nsew default input
rlabel metal1 s 350 356 538 430 6 B1
port 3 nsew default input
rlabel metal1 s 136 232 214 354 6 B2
port 4 nsew default input
rlabel metal1 s 24 354 214 430 6 B2
port 4 nsew default input
rlabel metal1 s 584 310 648 664 6 C
port 5 nsew default input
rlabel metal1 s 920 135 1196 181 6 ZN
port 6 nsew default output
rlabel metal1 s 920 181 984 195 6 ZN
port 6 nsew default output
rlabel metal1 s 430 135 636 181 6 ZN
port 6 nsew default output
rlabel metal1 s 590 181 636 195 6 ZN
port 6 nsew default output
rlabel metal1 s 590 195 984 241 6 ZN
port 6 nsew default output
rlabel metal1 s 920 241 984 573 6 ZN
port 6 nsew default output
rlabel metal1 s 273 632 319 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 724 1232 844 6 VDD
port 7 nsew power bidirectional abutment
rlabel nwell s -86 352 1318 870 6 VNW
port 8 nsew power bidirectional
rlabel pwell s -86 -86 1318 352 6 VPW
port 9 nsew ground bidirectional
rlabel metal1 s 0 -60 1232 60 8 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 734 60 802 149 6 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 163 6 VSS
port 10 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1232 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1295882
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1291726
<< end >>
