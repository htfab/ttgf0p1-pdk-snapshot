magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 1454 1486
<< nmos >>
rect 120 209 176 385
rect 280 209 336 385
rect 440 209 496 385
rect 688 209 744 385
rect 848 209 904 385
rect 1008 209 1064 385
<< pmos >>
rect 120 1015 176 1191
rect 280 1015 336 1191
rect 440 1015 496 1191
rect 688 1015 744 1191
rect 848 1015 904 1191
rect 1008 1015 1064 1191
<< ndiff >>
rect 32 371 120 385
rect 32 325 45 371
rect 91 325 120 371
rect 32 209 120 325
rect 176 268 280 385
rect 176 222 205 268
rect 251 222 280 268
rect 176 209 280 222
rect 336 209 440 385
rect 496 371 688 385
rect 496 325 569 371
rect 615 325 688 371
rect 496 209 688 325
rect 744 209 848 385
rect 904 268 1008 385
rect 904 222 933 268
rect 979 222 1008 268
rect 904 209 1008 222
rect 1064 371 1152 385
rect 1064 325 1093 371
rect 1139 325 1152 371
rect 1064 209 1152 325
<< pdiff >>
rect 32 1075 120 1191
rect 32 1029 45 1075
rect 91 1029 120 1075
rect 32 1015 120 1029
rect 176 1178 280 1191
rect 176 1132 205 1178
rect 251 1132 280 1178
rect 176 1015 280 1132
rect 336 1075 440 1191
rect 336 1029 365 1075
rect 411 1029 440 1075
rect 336 1015 440 1029
rect 496 1015 688 1191
rect 744 1075 848 1191
rect 744 1029 773 1075
rect 819 1029 848 1075
rect 744 1015 848 1029
rect 904 1178 1008 1191
rect 904 1132 933 1178
rect 979 1132 1008 1178
rect 904 1015 1008 1132
rect 1064 1075 1152 1191
rect 1064 1029 1093 1075
rect 1139 1029 1152 1075
rect 1064 1015 1152 1029
rect 556 943 628 1015
rect 556 897 569 943
rect 615 897 628 943
rect 556 884 628 897
<< ndiffc >>
rect 45 325 91 371
rect 205 222 251 268
rect 569 325 615 371
rect 933 222 979 268
rect 1093 325 1139 371
<< pdiffc >>
rect 45 1029 91 1075
rect 205 1132 251 1178
rect 365 1029 411 1075
rect 773 1029 819 1075
rect 933 1132 979 1178
rect 1093 1029 1139 1075
rect 569 897 615 943
<< psubdiff >>
rect 28 87 1340 100
rect 28 41 61 87
rect 1307 41 1340 87
rect 28 28 1340 41
<< nsubdiff >>
rect 28 1359 1340 1372
rect 28 1313 61 1359
rect 1307 1313 1340 1359
rect 28 1300 1340 1313
<< psubdiffcont >>
rect 61 41 1307 87
<< nsubdiffcont >>
rect 61 1313 1307 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 688 1191 744 1235
rect 848 1191 904 1235
rect 1008 1191 1064 1235
rect 120 914 176 1015
rect 280 914 336 1015
rect 120 901 336 914
rect 120 855 143 901
rect 189 855 336 901
rect 120 842 336 855
rect 440 782 496 1015
rect 384 769 496 782
rect 384 723 397 769
rect 443 723 496 769
rect 384 710 496 723
rect 688 650 744 1015
rect 848 914 904 1015
rect 1008 914 1064 1015
rect 848 901 1064 914
rect 848 855 965 901
rect 1011 855 1064 901
rect 848 842 1064 855
rect 32 637 744 650
rect 32 591 45 637
rect 91 591 744 637
rect 32 578 744 591
rect 792 637 1152 650
rect 792 591 805 637
rect 851 591 1093 637
rect 1139 591 1152 637
rect 792 578 1152 591
rect 120 505 336 518
rect 120 459 143 505
rect 189 459 336 505
rect 120 446 336 459
rect 384 505 496 518
rect 384 459 397 505
rect 443 459 496 505
rect 384 446 496 459
rect 120 385 176 446
rect 280 385 336 446
rect 440 385 496 446
rect 688 385 744 578
rect 848 385 904 578
rect 952 505 1064 518
rect 952 459 965 505
rect 1011 459 1064 505
rect 952 446 1064 459
rect 1008 385 1064 446
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
rect 688 165 744 209
rect 848 165 904 209
rect 1008 165 1064 209
<< polycontact >>
rect 143 855 189 901
rect 397 723 443 769
rect 965 855 1011 901
rect 45 591 91 637
rect 805 591 851 637
rect 1093 591 1139 637
rect 143 459 189 505
rect 397 459 443 505
rect 965 459 1011 505
<< metal1 >>
rect 0 1359 1368 1400
rect 0 1313 61 1359
rect 1307 1313 1368 1359
rect 0 1178 1368 1313
rect 0 1132 205 1178
rect 251 1132 933 1178
rect 979 1132 1368 1178
rect 42 1075 94 1086
rect 42 1029 45 1075
rect 91 1029 94 1075
rect 42 637 94 1029
rect 42 591 45 637
rect 91 591 94 637
rect 42 371 94 591
rect 42 325 45 371
rect 91 325 94 371
rect 42 314 94 325
rect 140 901 192 1086
rect 365 1075 819 1086
rect 411 1029 773 1075
rect 365 1018 819 1029
rect 140 855 143 901
rect 189 855 192 901
rect 140 505 192 855
rect 140 459 143 505
rect 189 459 192 505
rect 140 314 192 459
rect 238 954 290 972
rect 238 943 615 954
rect 238 897 569 943
rect 238 886 615 897
rect 962 901 1014 1086
rect 238 382 290 886
rect 962 855 965 901
rect 1011 855 1014 901
rect 397 769 854 780
rect 443 723 854 769
rect 397 712 854 723
rect 802 637 854 712
rect 802 591 805 637
rect 851 591 854 637
rect 802 580 854 591
rect 962 516 1014 855
rect 397 505 1014 516
rect 443 459 965 505
rect 1011 459 1014 505
rect 397 448 1014 459
rect 238 371 615 382
rect 238 325 569 371
rect 238 314 615 325
rect 962 314 1014 448
rect 1090 1075 1142 1086
rect 1090 1029 1093 1075
rect 1139 1029 1142 1075
rect 1090 637 1142 1029
rect 1090 591 1093 637
rect 1139 591 1142 637
rect 1090 371 1142 591
rect 1090 325 1093 371
rect 1139 325 1142 371
rect 1090 314 1142 325
rect 0 222 205 268
rect 251 222 933 268
rect 979 222 1368 268
rect 0 87 1368 222
rect 0 41 61 87
rect 1307 41 1368 87
rect 0 0 1368 41
<< labels >>
rlabel metal1 s 0 1132 1368 1400 4 vdd
port 3 nsew
rlabel metal1 s 0 0 1368 268 4 vss
port 5 nsew
rlabel metal1 s 140 314 192 1086 4 i0
port 7 nsew
rlabel metal1 s 238 314 290 972 4 q
port 9 nsew
rlabel metal1 s 962 314 1014 1086 4 i1
port 11 nsew
<< end >>
