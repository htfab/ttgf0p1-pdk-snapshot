magic
tech gf180mcuD
magscale 1 10
timestamp 1753432499
<< nwell >>
rect -86 354 2214 870
<< pwell >>
rect -86 -86 2214 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 756 68 812 268
rect 916 68 972 268
rect 1076 68 1132 268
rect 1236 68 1292 268
rect 1396 68 1452 268
rect 1556 68 1612 268
rect 1716 68 1772 268
rect 1876 68 1932 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
rect 1076 440 1132 716
rect 1236 440 1292 716
rect 1396 440 1452 716
rect 1556 440 1612 716
rect 1716 440 1772 716
rect 1876 440 1932 716
<< ndiff >>
rect 28 127 116 268
rect 28 81 41 127
rect 87 81 116 127
rect 28 68 116 81
rect 172 255 276 268
rect 172 209 201 255
rect 247 209 276 255
rect 172 68 276 209
rect 332 127 436 268
rect 332 81 361 127
rect 407 81 436 127
rect 332 68 436 81
rect 492 255 596 268
rect 492 209 521 255
rect 567 209 596 255
rect 492 68 596 209
rect 652 127 756 268
rect 652 81 681 127
rect 727 81 756 127
rect 652 68 756 81
rect 812 152 916 268
rect 812 106 841 152
rect 887 106 916 152
rect 812 68 916 106
rect 972 255 1076 268
rect 972 209 1001 255
rect 1047 209 1076 255
rect 972 68 1076 209
rect 1132 152 1236 268
rect 1132 106 1161 152
rect 1207 106 1236 152
rect 1132 68 1236 106
rect 1292 255 1396 268
rect 1292 209 1321 255
rect 1367 209 1396 255
rect 1292 68 1396 209
rect 1452 183 1556 268
rect 1452 137 1481 183
rect 1527 137 1556 183
rect 1452 68 1556 137
rect 1612 127 1716 268
rect 1612 81 1641 127
rect 1687 81 1716 127
rect 1612 68 1716 81
rect 1772 192 1876 268
rect 1772 146 1801 192
rect 1847 146 1876 192
rect 1772 68 1876 146
rect 1932 255 2024 268
rect 1932 81 1961 255
rect 2007 81 2024 255
rect 1932 68 2024 81
<< pdiff >>
rect 28 639 116 716
rect 28 593 41 639
rect 87 593 116 639
rect 28 440 116 593
rect 172 499 276 716
rect 172 453 201 499
rect 247 453 276 499
rect 172 440 276 453
rect 332 667 436 716
rect 332 621 361 667
rect 407 621 436 667
rect 332 440 436 621
rect 492 499 596 716
rect 492 453 521 499
rect 567 453 596 499
rect 492 440 596 453
rect 652 667 756 716
rect 652 621 681 667
rect 727 621 756 667
rect 652 440 756 621
rect 812 703 916 716
rect 812 657 841 703
rect 887 657 916 703
rect 812 440 916 657
rect 972 600 1076 716
rect 972 554 1001 600
rect 1047 554 1076 600
rect 972 440 1076 554
rect 1132 703 1236 716
rect 1132 657 1161 703
rect 1207 657 1236 703
rect 1132 440 1236 657
rect 1292 600 1396 716
rect 1292 554 1321 600
rect 1367 554 1396 600
rect 1292 440 1396 554
rect 1452 703 1556 716
rect 1452 657 1481 703
rect 1527 657 1556 703
rect 1452 440 1556 657
rect 1612 600 1716 716
rect 1612 554 1641 600
rect 1687 554 1716 600
rect 1612 440 1716 554
rect 1772 703 1876 716
rect 1772 657 1801 703
rect 1847 657 1876 703
rect 1772 440 1876 657
rect 1932 645 2024 716
rect 1932 599 1961 645
rect 2007 599 2024 645
rect 1932 440 2024 599
<< ndiffc >>
rect 41 81 87 127
rect 201 209 247 255
rect 361 81 407 127
rect 521 209 567 255
rect 681 81 727 127
rect 841 106 887 152
rect 1001 209 1047 255
rect 1161 106 1207 152
rect 1321 209 1367 255
rect 1481 137 1527 183
rect 1641 81 1687 127
rect 1801 146 1847 192
rect 1961 81 2007 255
<< pdiffc >>
rect 41 593 87 639
rect 201 453 247 499
rect 361 621 407 667
rect 521 453 567 499
rect 681 621 727 667
rect 841 657 887 703
rect 1001 554 1047 600
rect 1161 657 1207 703
rect 1321 554 1367 600
rect 1481 657 1527 703
rect 1641 554 1687 600
rect 1801 657 1847 703
rect 1961 599 2007 645
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 1076 716 1132 760
rect 1236 716 1292 760
rect 1396 716 1452 760
rect 1556 716 1612 760
rect 1716 716 1772 760
rect 1876 716 1932 760
rect 116 391 172 440
rect 276 391 332 440
rect 436 391 492 440
rect 596 391 652 440
rect 756 391 812 440
rect 76 378 652 391
rect 76 332 89 378
rect 504 332 652 378
rect 76 318 652 332
rect 713 378 812 391
rect 713 332 733 378
rect 779 332 812 378
rect 713 318 812 332
rect 116 268 172 318
rect 276 268 332 318
rect 436 268 492 318
rect 596 268 652 318
rect 756 268 812 318
rect 916 391 972 440
rect 1076 391 1132 440
rect 1236 391 1292 440
rect 1396 391 1452 440
rect 916 378 1452 391
rect 916 332 929 378
rect 1439 332 1452 378
rect 916 318 1452 332
rect 916 268 972 318
rect 1076 268 1132 318
rect 1236 268 1292 318
rect 1396 268 1452 318
rect 1556 391 1612 440
rect 1716 391 1772 440
rect 1876 391 1932 440
rect 1556 378 1932 391
rect 1556 332 1569 378
rect 1919 332 1932 378
rect 1556 318 1932 332
rect 1556 268 1612 318
rect 1716 268 1772 318
rect 1876 268 1932 318
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
rect 1076 24 1132 68
rect 1236 24 1292 68
rect 1396 24 1452 68
rect 1556 24 1612 68
rect 1716 24 1772 68
rect 1876 24 1932 68
<< polycontact >>
rect 89 332 504 378
rect 733 332 779 378
rect 929 332 1439 378
rect 1569 332 1919 378
<< metal1 >>
rect 0 724 2128 844
rect 841 703 887 724
rect 41 639 361 667
rect 87 621 361 639
rect 407 621 681 667
rect 727 621 738 667
rect 841 646 887 657
rect 1161 703 1207 724
rect 1161 646 1207 657
rect 1481 703 1527 724
rect 1481 646 1527 657
rect 1801 703 1847 724
rect 1801 646 1847 657
rect 41 574 87 593
rect 692 600 738 621
rect 1961 645 2007 660
rect 692 554 1001 600
rect 1047 554 1321 600
rect 1367 554 1641 600
rect 1687 599 1961 600
rect 1687 554 2007 599
rect 187 453 201 499
rect 247 453 521 499
rect 567 453 619 499
rect 76 378 504 391
rect 76 332 89 378
rect 76 318 504 332
rect 550 255 619 453
rect 752 462 1602 508
rect 752 391 798 462
rect 1556 391 1602 462
rect 713 378 798 391
rect 713 332 733 378
rect 779 332 798 378
rect 713 318 798 332
rect 916 378 1452 391
rect 916 332 929 378
rect 1439 332 1452 378
rect 916 318 1452 332
rect 1556 378 1932 391
rect 1556 332 1569 378
rect 1919 332 1932 378
rect 1556 318 1932 332
rect 1961 255 2007 274
rect 161 209 201 255
rect 247 209 521 255
rect 567 209 1001 255
rect 1047 209 1321 255
rect 1367 209 1379 255
rect 1481 198 1847 244
rect 1481 183 1527 198
rect 41 127 87 138
rect 41 60 87 81
rect 361 127 407 138
rect 361 60 407 81
rect 681 127 727 138
rect 820 106 841 152
rect 887 106 1161 152
rect 1207 137 1481 152
rect 1801 192 1847 198
rect 1207 106 1527 137
rect 1641 127 1687 138
rect 1801 131 1847 146
rect 681 60 727 81
rect 1641 60 1687 81
rect 1961 60 2007 81
rect 0 -60 2128 60
<< labels >>
flabel metal1 s 0 724 2128 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 2128 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 550 209 619 499 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 76 318 504 391 0 FreeSans 200 0 0 0 C
port 6 nsew signal input
flabel metal1 1556 318 1932 391 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel metal1 916 318 1452 391 0 FreeSans 200 0 0 0 A
port 8 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 2128 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
