magic
tech gf180mcuD
timestamp 1755069416
<< properties >>
string gencell eFuse_0
string library gf180mcu
string parameter m=1
<< end >>
