magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 770 1486
<< nmos >>
rect 120 209 176 385
rect 280 209 336 385
rect 440 209 496 385
<< pmos >>
rect 120 1015 176 1191
rect 280 1015 336 1191
rect 440 1015 496 1191
<< ndiff >>
rect 32 371 120 385
rect 32 325 45 371
rect 91 325 120 371
rect 32 209 120 325
rect 176 268 280 385
rect 176 222 205 268
rect 251 222 280 268
rect 176 209 280 222
rect 336 371 440 385
rect 336 325 365 371
rect 411 325 440 371
rect 336 209 440 325
rect 496 371 620 385
rect 496 325 561 371
rect 607 325 620 371
rect 496 209 620 325
<< pdiff >>
rect 32 1178 120 1191
rect 32 1132 45 1178
rect 91 1132 120 1178
rect 32 1015 120 1132
rect 176 1015 280 1191
rect 336 1075 440 1191
rect 336 1029 365 1075
rect 411 1029 440 1075
rect 336 1015 440 1029
rect 496 1178 620 1191
rect 496 1132 561 1178
rect 607 1132 620 1178
rect 496 1015 620 1132
<< ndiffc >>
rect 45 325 91 371
rect 205 222 251 268
rect 365 325 411 371
rect 561 325 607 371
<< pdiffc >>
rect 45 1132 91 1178
rect 365 1029 411 1075
rect 561 1132 607 1178
<< psubdiff >>
rect 28 87 656 100
rect 28 41 69 87
rect 615 41 656 87
rect 28 28 656 41
<< nsubdiff >>
rect 28 1359 656 1372
rect 28 1313 69 1359
rect 615 1313 656 1359
rect 28 1300 656 1313
<< psubdiffcont >>
rect 69 41 615 87
<< nsubdiffcont >>
rect 69 1313 615 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 120 716 176 1015
rect 280 716 336 1015
rect 32 703 176 716
rect 32 657 45 703
rect 91 657 176 703
rect 32 644 176 657
rect 224 703 336 716
rect 224 657 237 703
rect 283 657 336 703
rect 224 644 336 657
rect 120 385 176 644
rect 280 385 336 644
rect 440 716 496 1015
rect 440 703 522 716
rect 440 657 463 703
rect 509 657 522 703
rect 440 644 522 657
rect 440 385 496 644
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
<< polycontact >>
rect 45 657 91 703
rect 237 657 283 703
rect 463 657 509 703
<< metal1 >>
rect 0 1359 684 1400
rect 0 1313 69 1359
rect 615 1313 684 1359
rect 0 1178 684 1313
rect 0 1132 45 1178
rect 91 1132 561 1178
rect 607 1132 684 1178
rect 42 703 94 1086
rect 42 657 45 703
rect 91 657 94 703
rect 42 428 94 657
rect 234 703 286 1086
rect 365 1075 610 1086
rect 411 1029 610 1075
rect 365 1018 610 1029
rect 234 657 237 703
rect 283 657 286 703
rect 234 428 286 657
rect 460 703 512 972
rect 460 657 463 703
rect 509 657 512 703
rect 45 371 411 382
rect 91 325 365 371
rect 45 314 411 325
rect 460 314 512 657
rect 558 371 610 1018
rect 558 325 561 371
rect 607 325 610 371
rect 558 314 610 325
rect 0 222 205 268
rect 251 222 684 268
rect 0 87 684 222
rect 0 41 69 87
rect 615 41 684 87
rect 0 0 684 41
<< labels >>
rlabel metal1 s 0 1132 684 1400 4 vdd
port 3 nsew
rlabel metal1 s 0 0 684 268 4 vss
port 5 nsew
rlabel metal1 s 42 428 94 1086 4 i0
port 7 nsew
rlabel metal1 s 234 428 286 1086 4 i1
port 9 nsew
rlabel metal1 s 558 314 610 1086 4 nq
port 11 nsew
rlabel metal1 s 460 314 512 972 4 i2
port 13 nsew
<< end >>
