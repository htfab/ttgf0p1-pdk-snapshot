magic
tech gf180mcuD
timestamp 1755005639
<< properties >>
string GDS_END 335378
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 334606
<< end >>
