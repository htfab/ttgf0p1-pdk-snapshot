magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 998 1486
<< nmos >>
rect 120 209 176 584
rect 280 209 336 584
rect 440 209 496 584
rect 600 209 656 584
<< pmos >>
rect 120 776 176 1191
rect 280 776 336 1191
rect 440 776 496 1191
rect 600 776 656 1191
<< ndiff >>
rect 32 268 120 584
rect 32 222 45 268
rect 91 222 120 268
rect 32 209 120 222
rect 176 209 280 584
rect 336 209 440 584
rect 496 209 600 584
rect 656 571 744 584
rect 656 325 685 571
rect 731 325 744 571
rect 656 209 744 325
<< pdiff >>
rect 32 1178 120 1191
rect 32 1132 45 1178
rect 91 1132 120 1178
rect 32 776 120 1132
rect 176 1055 280 1191
rect 176 809 205 1055
rect 251 809 280 1055
rect 176 776 280 809
rect 336 1178 440 1191
rect 336 1132 365 1178
rect 411 1132 440 1178
rect 336 776 440 1132
rect 496 1055 600 1191
rect 496 809 525 1055
rect 571 809 600 1055
rect 496 776 600 809
rect 656 1178 744 1191
rect 656 1132 685 1178
rect 731 1132 744 1178
rect 656 776 744 1132
<< ndiffc >>
rect 45 222 91 268
rect 685 325 731 571
<< pdiffc >>
rect 45 1132 91 1178
rect 205 809 251 1055
rect 365 1132 411 1178
rect 525 809 571 1055
rect 685 1132 731 1178
<< psubdiff >>
rect 28 87 884 100
rect 28 41 83 87
rect 829 41 884 87
rect 28 28 884 41
<< nsubdiff >>
rect 28 1359 884 1372
rect 28 1313 83 1359
rect 829 1313 884 1359
rect 28 1300 884 1313
<< psubdiffcont >>
rect 83 41 829 87
<< nsubdiffcont >>
rect 83 1313 829 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 600 1191 656 1235
rect 120 716 176 776
rect 280 716 336 776
rect 440 716 496 776
rect 600 716 656 776
rect 32 703 176 716
rect 32 657 45 703
rect 91 657 176 703
rect 32 644 176 657
rect 224 703 336 716
rect 224 657 237 703
rect 283 657 336 703
rect 224 644 336 657
rect 384 703 496 716
rect 384 657 397 703
rect 443 657 496 703
rect 384 644 496 657
rect 544 703 656 716
rect 544 657 557 703
rect 603 657 656 703
rect 544 644 656 657
rect 120 584 176 644
rect 280 584 336 644
rect 440 584 496 644
rect 600 584 656 644
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
rect 600 165 656 209
<< polycontact >>
rect 45 657 91 703
rect 237 657 283 703
rect 397 657 443 703
rect 557 657 603 703
<< metal1 >>
rect 0 1359 912 1400
rect 0 1313 83 1359
rect 829 1313 912 1359
rect 0 1178 912 1313
rect 0 1132 45 1178
rect 91 1132 365 1178
rect 411 1132 685 1178
rect 731 1132 912 1178
rect 42 703 94 1086
rect 205 1055 734 1086
rect 251 809 525 1055
rect 571 809 734 1055
rect 205 798 734 809
rect 42 657 45 703
rect 91 657 94 703
rect 42 314 94 657
rect 234 703 286 752
rect 234 657 237 703
rect 283 657 286 703
rect 234 314 286 657
rect 394 703 446 752
rect 394 657 397 703
rect 443 657 446 703
rect 394 314 446 657
rect 554 703 606 752
rect 554 657 557 703
rect 603 657 606 703
rect 554 314 606 657
rect 682 571 734 798
rect 682 325 685 571
rect 731 325 734 571
rect 682 314 734 325
rect 0 222 45 268
rect 91 222 912 268
rect 0 87 912 222
rect 0 41 83 87
rect 829 41 912 87
rect 0 0 912 41
<< labels >>
rlabel metal1 s 0 0 912 268 4 vss
port 3 nsew
rlabel metal1 s 0 1132 912 1400 4 vdd
port 5 nsew
rlabel metal1 s 42 314 94 1086 4 i0
port 7 nsew
rlabel metal1 s 682 314 734 1086 4 nq
port 9 nsew
rlabel metal1 s 234 314 286 752 4 i1
port 11 nsew
rlabel metal1 s 394 314 446 752 4 i2
port 13 nsew
rlabel metal1 s 554 314 606 752 4 i3
port 15 nsew
<< end >>
