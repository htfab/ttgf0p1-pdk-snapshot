magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< isosubstrate >>
rect 1385 -83 2701 2911
<< nwell >>
rect -83 1213 1045 2911
rect 1385 1213 2701 2911
<< mvnmos >>
rect 286 270 426 870
rect 530 270 670 870
rect 1913 270 2053 870
rect 2157 270 2297 870
<< mvpmos >>
rect 286 1958 426 2558
rect 530 1958 670 2558
rect 1913 1358 2053 2558
rect 2157 1358 2297 2558
<< mvndiff >>
rect 198 857 286 870
rect 198 811 211 857
rect 257 811 286 857
rect 198 752 286 811
rect 198 706 211 752
rect 257 706 286 752
rect 198 647 286 706
rect 198 601 211 647
rect 257 601 286 647
rect 198 541 286 601
rect 198 495 211 541
rect 257 495 286 541
rect 198 435 286 495
rect 198 389 211 435
rect 257 389 286 435
rect 198 329 286 389
rect 198 283 211 329
rect 257 283 286 329
rect 198 270 286 283
rect 426 857 530 870
rect 426 811 455 857
rect 501 811 530 857
rect 426 752 530 811
rect 426 706 455 752
rect 501 706 530 752
rect 426 647 530 706
rect 426 601 455 647
rect 501 601 530 647
rect 426 541 530 601
rect 426 495 455 541
rect 501 495 530 541
rect 426 435 530 495
rect 426 389 455 435
rect 501 389 530 435
rect 426 329 530 389
rect 426 283 455 329
rect 501 283 530 329
rect 426 270 530 283
rect 670 857 758 870
rect 670 811 699 857
rect 745 811 758 857
rect 670 752 758 811
rect 670 706 699 752
rect 745 706 758 752
rect 670 647 758 706
rect 670 601 699 647
rect 745 601 758 647
rect 670 541 758 601
rect 670 495 699 541
rect 745 495 758 541
rect 670 435 758 495
rect 670 389 699 435
rect 745 389 758 435
rect 670 329 758 389
rect 670 283 699 329
rect 745 283 758 329
rect 670 270 758 283
rect 1825 857 1913 870
rect 1825 811 1838 857
rect 1884 811 1913 857
rect 1825 752 1913 811
rect 1825 706 1838 752
rect 1884 706 1913 752
rect 1825 647 1913 706
rect 1825 601 1838 647
rect 1884 601 1913 647
rect 1825 541 1913 601
rect 1825 495 1838 541
rect 1884 495 1913 541
rect 1825 435 1913 495
rect 1825 389 1838 435
rect 1884 389 1913 435
rect 1825 329 1913 389
rect 1825 283 1838 329
rect 1884 283 1913 329
rect 1825 270 1913 283
rect 2053 857 2157 870
rect 2053 811 2082 857
rect 2128 811 2157 857
rect 2053 752 2157 811
rect 2053 706 2082 752
rect 2128 706 2157 752
rect 2053 647 2157 706
rect 2053 601 2082 647
rect 2128 601 2157 647
rect 2053 541 2157 601
rect 2053 495 2082 541
rect 2128 495 2157 541
rect 2053 435 2157 495
rect 2053 389 2082 435
rect 2128 389 2157 435
rect 2053 329 2157 389
rect 2053 283 2082 329
rect 2128 283 2157 329
rect 2053 270 2157 283
rect 2297 857 2385 870
rect 2297 811 2326 857
rect 2372 811 2385 857
rect 2297 752 2385 811
rect 2297 706 2326 752
rect 2372 706 2385 752
rect 2297 647 2385 706
rect 2297 601 2326 647
rect 2372 601 2385 647
rect 2297 541 2385 601
rect 2297 495 2326 541
rect 2372 495 2385 541
rect 2297 435 2385 495
rect 2297 389 2326 435
rect 2372 389 2385 435
rect 2297 329 2385 389
rect 2297 283 2326 329
rect 2372 283 2385 329
rect 2297 270 2385 283
<< mvpdiff >>
rect 198 2545 286 2558
rect 198 2499 211 2545
rect 257 2499 286 2545
rect 198 2440 286 2499
rect 198 2394 211 2440
rect 257 2394 286 2440
rect 198 2335 286 2394
rect 198 2289 211 2335
rect 257 2289 286 2335
rect 198 2229 286 2289
rect 198 2183 211 2229
rect 257 2183 286 2229
rect 198 2123 286 2183
rect 198 2077 211 2123
rect 257 2077 286 2123
rect 198 2017 286 2077
rect 198 1971 211 2017
rect 257 1971 286 2017
rect 198 1958 286 1971
rect 426 2545 530 2558
rect 426 2499 455 2545
rect 501 2499 530 2545
rect 426 2440 530 2499
rect 426 2394 455 2440
rect 501 2394 530 2440
rect 426 2335 530 2394
rect 426 2289 455 2335
rect 501 2289 530 2335
rect 426 2229 530 2289
rect 426 2183 455 2229
rect 501 2183 530 2229
rect 426 2123 530 2183
rect 426 2077 455 2123
rect 501 2077 530 2123
rect 426 2017 530 2077
rect 426 1971 455 2017
rect 501 1971 530 2017
rect 426 1958 530 1971
rect 670 2545 758 2558
rect 670 2499 699 2545
rect 745 2499 758 2545
rect 670 2440 758 2499
rect 670 2394 699 2440
rect 745 2394 758 2440
rect 670 2335 758 2394
rect 670 2289 699 2335
rect 745 2289 758 2335
rect 670 2229 758 2289
rect 670 2183 699 2229
rect 745 2183 758 2229
rect 670 2123 758 2183
rect 670 2077 699 2123
rect 745 2077 758 2123
rect 670 2017 758 2077
rect 670 1971 699 2017
rect 745 1971 758 2017
rect 670 1958 758 1971
rect 1825 2545 1913 2558
rect 1825 1989 1838 2545
rect 1884 1989 1913 2545
rect 1825 1932 1913 1989
rect 1825 1886 1838 1932
rect 1884 1886 1913 1932
rect 1825 1829 1913 1886
rect 1825 1783 1838 1829
rect 1884 1783 1913 1829
rect 1825 1726 1913 1783
rect 1825 1680 1838 1726
rect 1884 1680 1913 1726
rect 1825 1623 1913 1680
rect 1825 1577 1838 1623
rect 1884 1577 1913 1623
rect 1825 1520 1913 1577
rect 1825 1474 1838 1520
rect 1884 1474 1913 1520
rect 1825 1417 1913 1474
rect 1825 1371 1838 1417
rect 1884 1371 1913 1417
rect 1825 1358 1913 1371
rect 2053 2545 2157 2558
rect 2053 1989 2082 2545
rect 2128 1989 2157 2545
rect 2053 1932 2157 1989
rect 2053 1886 2082 1932
rect 2128 1886 2157 1932
rect 2053 1829 2157 1886
rect 2053 1783 2082 1829
rect 2128 1783 2157 1829
rect 2053 1726 2157 1783
rect 2053 1680 2082 1726
rect 2128 1680 2157 1726
rect 2053 1623 2157 1680
rect 2053 1577 2082 1623
rect 2128 1577 2157 1623
rect 2053 1520 2157 1577
rect 2053 1474 2082 1520
rect 2128 1474 2157 1520
rect 2053 1417 2157 1474
rect 2053 1371 2082 1417
rect 2128 1371 2157 1417
rect 2053 1358 2157 1371
rect 2297 2545 2385 2558
rect 2297 1989 2326 2545
rect 2372 1989 2385 2545
rect 2297 1932 2385 1989
rect 2297 1886 2326 1932
rect 2372 1886 2385 1932
rect 2297 1829 2385 1886
rect 2297 1783 2326 1829
rect 2372 1783 2385 1829
rect 2297 1726 2385 1783
rect 2297 1680 2326 1726
rect 2372 1680 2385 1726
rect 2297 1623 2385 1680
rect 2297 1577 2326 1623
rect 2372 1577 2385 1623
rect 2297 1520 2385 1577
rect 2297 1474 2326 1520
rect 2372 1474 2385 1520
rect 2297 1417 2385 1474
rect 2297 1371 2326 1417
rect 2372 1371 2385 1417
rect 2297 1358 2385 1371
<< mvndiffc >>
rect 211 811 257 857
rect 211 706 257 752
rect 211 601 257 647
rect 211 495 257 541
rect 211 389 257 435
rect 211 283 257 329
rect 455 811 501 857
rect 455 706 501 752
rect 455 601 501 647
rect 455 495 501 541
rect 455 389 501 435
rect 455 283 501 329
rect 699 811 745 857
rect 699 706 745 752
rect 699 601 745 647
rect 699 495 745 541
rect 699 389 745 435
rect 699 283 745 329
rect 1838 811 1884 857
rect 1838 706 1884 752
rect 1838 601 1884 647
rect 1838 495 1884 541
rect 1838 389 1884 435
rect 1838 283 1884 329
rect 2082 811 2128 857
rect 2082 706 2128 752
rect 2082 601 2128 647
rect 2082 495 2128 541
rect 2082 389 2128 435
rect 2082 283 2128 329
rect 2326 811 2372 857
rect 2326 706 2372 752
rect 2326 601 2372 647
rect 2326 495 2372 541
rect 2326 389 2372 435
rect 2326 283 2372 329
<< mvpdiffc >>
rect 211 2499 257 2545
rect 211 2394 257 2440
rect 211 2289 257 2335
rect 211 2183 257 2229
rect 211 2077 257 2123
rect 211 1971 257 2017
rect 455 2499 501 2545
rect 455 2394 501 2440
rect 455 2289 501 2335
rect 455 2183 501 2229
rect 455 2077 501 2123
rect 455 1971 501 2017
rect 699 2499 745 2545
rect 699 2394 745 2440
rect 699 2289 745 2335
rect 699 2183 745 2229
rect 699 2077 745 2123
rect 699 1971 745 2017
rect 1838 1989 1884 2545
rect 1838 1886 1884 1932
rect 1838 1783 1884 1829
rect 1838 1680 1884 1726
rect 1838 1577 1884 1623
rect 1838 1474 1884 1520
rect 1838 1371 1884 1417
rect 2082 1989 2128 2545
rect 2082 1886 2128 1932
rect 2082 1783 2128 1829
rect 2082 1680 2128 1726
rect 2082 1577 2128 1623
rect 2082 1474 2128 1520
rect 2082 1371 2128 1417
rect 2326 1989 2372 2545
rect 2326 1886 2372 1932
rect 2326 1783 2372 1829
rect 2326 1680 2372 1726
rect 2326 1577 2372 1623
rect 2326 1474 2372 1520
rect 2326 1371 2372 1417
<< psubdiff >>
rect 0 1008 90 1030
rect 0 22 22 1008
rect 68 90 90 1008
rect 872 914 962 936
rect 872 90 894 914
rect 68 68 894 90
rect 68 22 176 68
rect 786 22 894 68
rect 940 22 962 914
rect 0 0 962 22
rect 1468 914 1558 936
rect 1468 22 1490 914
rect 1536 90 1558 914
rect 2528 1008 2618 1030
rect 2528 90 2550 1008
rect 1536 68 2550 90
rect 1536 22 1644 68
rect 2442 22 2550 68
rect 2596 22 2618 1008
rect 1468 0 2618 22
<< nsubdiff >>
rect 0 2806 962 2828
rect 0 1350 22 2806
rect 68 2760 176 2806
rect 786 2760 894 2806
rect 68 2738 894 2760
rect 68 1350 90 2738
rect 0 1328 90 1350
rect 872 1350 894 2738
rect 940 1350 962 2806
rect 872 1328 962 1350
rect 1468 2806 2618 2828
rect 1468 1350 1490 2806
rect 1536 2760 1644 2806
rect 2442 2760 2550 2806
rect 1536 2738 2550 2760
rect 1536 1350 1558 2738
rect 1468 1328 1558 1350
rect 2528 1350 2550 2738
rect 2596 1350 2618 2806
rect 2528 1328 2618 1350
<< psubdiffcont >>
rect 22 22 68 1008
rect 176 22 786 68
rect 894 22 940 914
rect 1490 22 1536 914
rect 1644 22 2442 68
rect 2550 22 2596 1008
<< nsubdiffcont >>
rect 22 1350 68 2806
rect 176 2760 786 2806
rect 894 1350 940 2806
rect 1490 1350 1536 2806
rect 1644 2760 2442 2806
rect 2550 1350 2596 2806
<< polysilicon >>
rect 286 2558 426 2602
rect 530 2558 670 2602
rect 286 1537 426 1958
rect 286 1397 333 1537
rect 379 1397 426 1537
rect 286 870 426 1397
rect 530 1537 670 1958
rect 530 1397 577 1537
rect 623 1397 670 1537
rect 530 870 670 1397
rect 1913 2558 2053 2602
rect 2157 2558 2297 2602
rect 1913 1213 2053 1358
rect 1697 1178 2053 1213
rect 1697 1038 1716 1178
rect 1762 1038 2053 1178
rect 1697 1002 2053 1038
rect 286 226 426 270
rect 530 226 670 270
rect 1913 870 2053 1002
rect 2157 1178 2297 1358
rect 2157 1038 2196 1178
rect 2242 1038 2297 1178
rect 2157 870 2297 1038
rect 1913 226 2053 270
rect 2157 226 2297 270
<< polycontact >>
rect 333 1397 379 1537
rect 577 1397 623 1537
rect 1716 1038 1762 1178
rect 2196 1038 2242 1178
<< metal1 >>
rect 11 2806 951 2817
rect 11 1350 22 2806
rect 68 2760 176 2806
rect 786 2760 894 2806
rect 68 2749 894 2760
rect 68 1350 79 2749
rect 196 2545 272 2749
rect 196 2499 211 2545
rect 257 2499 272 2545
rect 196 2440 272 2499
rect 196 2394 211 2440
rect 257 2394 272 2440
rect 196 2335 272 2394
rect 196 2289 211 2335
rect 257 2289 272 2335
rect 196 2229 272 2289
rect 196 2183 211 2229
rect 257 2183 272 2229
rect 196 2123 272 2183
rect 196 2077 211 2123
rect 257 2077 272 2123
rect 196 2017 272 2077
rect 196 1971 211 2017
rect 257 1971 272 2017
rect 196 1958 272 1971
rect 440 2545 516 2558
rect 440 2499 455 2545
rect 501 2499 516 2545
rect 440 2440 516 2499
rect 440 2394 455 2440
rect 501 2394 516 2440
rect 440 2335 516 2394
rect 440 2289 455 2335
rect 501 2289 516 2335
rect 440 2229 516 2289
rect 440 2183 455 2229
rect 501 2183 516 2229
rect 440 2123 516 2183
rect 440 2077 455 2123
rect 501 2077 516 2123
rect 440 2017 516 2077
rect 440 1971 455 2017
rect 501 1971 516 2017
rect 440 1794 516 1971
rect 684 2545 760 2749
rect 684 2499 699 2545
rect 745 2499 760 2545
rect 684 2440 760 2499
rect 684 2394 699 2440
rect 745 2394 760 2440
rect 684 2335 760 2394
rect 684 2289 699 2335
rect 745 2289 760 2335
rect 684 2229 760 2289
rect 684 2183 699 2229
rect 745 2183 760 2229
rect 684 2123 760 2183
rect 684 2077 699 2123
rect 745 2077 760 2123
rect 684 2017 760 2077
rect 684 1971 699 2017
rect 745 1971 760 2017
rect 684 1958 760 1971
rect 440 1718 760 1794
rect 322 1537 390 1548
rect 322 1397 333 1537
rect 379 1397 390 1537
rect 322 1386 390 1397
rect 566 1537 634 1548
rect 566 1397 577 1537
rect 623 1397 634 1537
rect 566 1386 634 1397
rect 11 1339 79 1350
rect 684 1197 760 1718
rect 883 1350 894 2749
rect 940 1350 951 2806
rect 883 1339 951 1350
rect 1479 2806 2607 2817
rect 1479 1350 1490 2806
rect 1536 2760 1644 2806
rect 2442 2760 2550 2806
rect 1536 2749 2550 2760
rect 1536 1350 1547 2749
rect 1479 1339 1547 1350
rect 1823 2545 1899 2558
rect 1823 1989 1838 2545
rect 1884 1989 1899 2545
rect 1823 1932 1899 1989
rect 1823 1886 1838 1932
rect 1884 1886 1899 1932
rect 1823 1829 1899 1886
rect 1823 1783 1838 1829
rect 1884 1783 1899 1829
rect 1823 1726 1899 1783
rect 1823 1680 1838 1726
rect 1884 1680 1899 1726
rect 1823 1623 1899 1680
rect 1823 1577 1838 1623
rect 1884 1577 1899 1623
rect 1823 1520 1899 1577
rect 1823 1474 1838 1520
rect 1884 1474 1899 1520
rect 1823 1417 1899 1474
rect 1823 1371 1838 1417
rect 1884 1371 1899 1417
rect 1823 1197 1899 1371
rect 2067 2545 2143 2749
rect 2067 1989 2082 2545
rect 2128 1989 2143 2545
rect 2067 1932 2143 1989
rect 2067 1886 2082 1932
rect 2128 1886 2143 1932
rect 2067 1829 2143 1886
rect 2067 1783 2082 1829
rect 2128 1783 2143 1829
rect 2067 1726 2143 1783
rect 2067 1680 2082 1726
rect 2128 1680 2143 1726
rect 2067 1623 2143 1680
rect 2067 1577 2082 1623
rect 2128 1577 2143 1623
rect 2067 1520 2143 1577
rect 2067 1474 2082 1520
rect 2128 1474 2143 1520
rect 2067 1417 2143 1474
rect 2067 1371 2082 1417
rect 2128 1371 2143 1417
rect 2067 1358 2143 1371
rect 2311 2545 2387 2558
rect 2311 1989 2326 2545
rect 2372 1989 2387 2545
rect 2311 1932 2387 1989
rect 2311 1886 2326 1932
rect 2372 1886 2387 1932
rect 2311 1829 2387 1886
rect 2311 1783 2326 1829
rect 2372 1783 2387 1829
rect 2311 1726 2387 1783
rect 2311 1680 2326 1726
rect 2372 1680 2387 1726
rect 2311 1623 2387 1680
rect 2311 1577 2326 1623
rect 2372 1577 2387 1623
rect 2311 1520 2387 1577
rect 2311 1474 2326 1520
rect 2372 1474 2387 1520
rect 2311 1417 2387 1474
rect 2311 1371 2326 1417
rect 2372 1371 2387 1417
rect 684 1178 1773 1197
rect 684 1038 1716 1178
rect 1762 1038 1773 1178
rect 684 1019 1773 1038
rect 1823 1178 2261 1197
rect 1823 1038 2196 1178
rect 2242 1038 2261 1178
rect 1823 1019 2261 1038
rect 11 1008 79 1019
rect 11 22 22 1008
rect 68 79 79 1008
rect 196 857 272 870
rect 196 811 211 857
rect 257 811 272 857
rect 196 752 272 811
rect 196 706 211 752
rect 257 706 272 752
rect 196 647 272 706
rect 196 601 211 647
rect 257 601 272 647
rect 196 541 272 601
rect 196 495 211 541
rect 257 495 272 541
rect 196 435 272 495
rect 196 389 211 435
rect 257 389 272 435
rect 196 329 272 389
rect 196 283 211 329
rect 257 283 272 329
rect 196 79 272 283
rect 455 857 501 870
rect 455 752 501 811
rect 455 647 501 706
rect 455 541 501 601
rect 455 435 501 495
rect 455 329 501 389
rect 455 270 501 283
rect 684 857 760 1019
rect 684 811 699 857
rect 745 811 760 857
rect 684 752 760 811
rect 684 706 699 752
rect 745 706 760 752
rect 684 647 760 706
rect 684 601 699 647
rect 745 601 760 647
rect 684 541 760 601
rect 684 495 699 541
rect 745 495 760 541
rect 684 435 760 495
rect 684 389 699 435
rect 745 389 760 435
rect 684 329 760 389
rect 684 283 699 329
rect 745 283 760 329
rect 684 270 760 283
rect 883 914 951 925
rect 883 79 894 914
rect 68 68 894 79
rect 68 22 176 68
rect 786 22 894 68
rect 940 22 951 914
rect 11 11 951 22
rect 1479 914 1547 925
rect 1479 22 1490 914
rect 1536 79 1547 914
rect 1823 857 1899 1019
rect 1823 811 1838 857
rect 1884 811 1899 857
rect 1823 752 1899 811
rect 1823 706 1838 752
rect 1884 706 1899 752
rect 1823 647 1899 706
rect 1823 601 1838 647
rect 1884 601 1899 647
rect 1823 541 1899 601
rect 1823 495 1838 541
rect 1884 495 1899 541
rect 1823 435 1899 495
rect 1823 389 1838 435
rect 1884 389 1899 435
rect 1823 329 1899 389
rect 1823 283 1838 329
rect 1884 283 1899 329
rect 1823 270 1899 283
rect 2067 857 2143 870
rect 2067 811 2082 857
rect 2128 811 2143 857
rect 2067 752 2143 811
rect 2067 706 2082 752
rect 2128 706 2143 752
rect 2067 647 2143 706
rect 2067 601 2082 647
rect 2128 601 2143 647
rect 2067 541 2143 601
rect 2067 495 2082 541
rect 2128 495 2143 541
rect 2067 435 2143 495
rect 2067 389 2082 435
rect 2128 389 2143 435
rect 2067 329 2143 389
rect 2067 283 2082 329
rect 2128 283 2143 329
rect 2067 79 2143 283
rect 2311 857 2387 1371
rect 2539 1350 2550 2749
rect 2596 1350 2607 2806
rect 2539 1339 2607 1350
rect 2311 811 2326 857
rect 2372 811 2387 857
rect 2311 752 2387 811
rect 2311 706 2326 752
rect 2372 706 2387 752
rect 2311 647 2387 706
rect 2311 601 2326 647
rect 2372 601 2387 647
rect 2311 541 2387 601
rect 2311 495 2326 541
rect 2372 495 2387 541
rect 2311 435 2387 495
rect 2311 389 2326 435
rect 2372 389 2387 435
rect 2311 329 2387 389
rect 2311 283 2326 329
rect 2372 283 2387 329
rect 2311 270 2387 283
rect 2539 1008 2607 1019
rect 2539 79 2550 1008
rect 1536 68 2550 79
rect 1536 22 1644 68
rect 2442 22 2550 68
rect 2596 22 2607 1008
rect 1479 11 2607 22
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_0
timestamp 1755005639
transform 1 0 917 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_1
timestamp 1755005639
transform 1 0 45 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_2
timestamp 1755005639
transform 1 0 1513 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145223  M1_NWELL_CDNS_40661953145223_3
timestamp 1755005639
transform 1 0 2573 0 1 2078
box 0 0 1 1
use M1_NWELL_CDNS_40661953145225  M1_NWELL_CDNS_40661953145225_0
timestamp 1755005639
transform 1 0 2043 0 1 2783
box 0 0 1 1
use M1_NWELL_CDNS_40661953145272  M1_NWELL_CDNS_40661953145272_0
timestamp 1755005639
transform 1 0 481 0 1 2783
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_0
timestamp 1755005639
transform -1 0 356 0 1 1467
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_1
timestamp 1755005639
transform -1 0 600 0 1 1467
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_2
timestamp 1755005639
transform 1 0 1739 0 1 1108
box 0 0 1 1
use M1_POLY2_CDNS_40661953145222  M1_POLY2_CDNS_40661953145222_3
timestamp 1755005639
transform 1 0 2219 0 1 1108
box 0 0 1 1
use M1_PSUB_CDNS_40661953145221  M1_PSUB_CDNS_40661953145221_0
timestamp 1755005639
transform 1 0 2043 0 -1 45
box 0 0 1 1
use M1_PSUB_CDNS_40661953145226  M1_PSUB_CDNS_40661953145226_0
timestamp 1755005639
transform 1 0 45 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661953145226  M1_PSUB_CDNS_40661953145226_1
timestamp 1755005639
transform 1 0 2573 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661953145228  M1_PSUB_CDNS_40661953145228_0
timestamp 1755005639
transform 1 0 917 0 -1 468
box 0 0 1 1
use M1_PSUB_CDNS_40661953145228  M1_PSUB_CDNS_40661953145228_1
timestamp 1755005639
transform 1 0 1513 0 -1 468
box 0 0 1 1
use M1_PSUB_CDNS_40661953145271  M1_PSUB_CDNS_40661953145271_0
timestamp 1755005639
transform 1 0 481 0 -1 45
box 0 0 1 1
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_0
timestamp 1755005639
transform 1 0 2157 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_1
timestamp 1755005639
transform 1 0 530 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_2
timestamp 1755005639
transform 1 0 286 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195314511  nmos_6p0_CDNS_4066195314511_3
timestamp 1755005639
transform 1 0 1913 0 1 270
box 0 0 1 1
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_0
timestamp 1755005639
transform -1 0 670 0 1 1958
box 0 0 1 1
use pmos_6p0_CDNS_4066195314512  pmos_6p0_CDNS_4066195314512_1
timestamp 1755005639
transform 1 0 286 0 1 1958
box 0 0 1 1
use pmos_6p0_CDNS_4066195314513  pmos_6p0_CDNS_4066195314513_0
timestamp 1755005639
transform 1 0 2157 0 1 1358
box 0 0 1 1
use pmos_6p0_CDNS_4066195314513  pmos_6p0_CDNS_4066195314513_1
timestamp 1755005639
transform 1 0 1913 0 1 1358
box 0 0 1 1
<< labels >>
rlabel metal1 s 263 45 263 45 4 VSS
port 1 nsew
rlabel metal1 s 2349 1100 2349 1100 4 AB
port 2 nsew
rlabel metal1 s 604 1468 604 1468 4 A
port 3 nsew
rlabel metal1 s 2245 45 2245 45 4 DVSS
port 4 nsew
rlabel metal1 s 2254 2788 2254 2788 4 DVDD
port 5 nsew
rlabel metal1 s 349 1468 349 1468 4 OE
port 6 nsew
rlabel metal1 s 92 2788 92 2788 4 VDD
port 7 nsew
<< properties >>
string GDS_END 1488392
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1484568
string path 5.850 1.050 5.850 21.750 
<< end >>
