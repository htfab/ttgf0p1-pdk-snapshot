* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__dfxtp_2.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__dfxtp_2 VDD VNW VPW VSS CLK D Q
X0 a_1709_68# a_28_68# a_1315_24# VNW pfet_03v3 ad=0.8418p pd=2.6u as=0.83145p ps=2.585u w=1.38u l=0.28u
X1 a_853_68# D a_629_68# VPW nfet_03v3 ad=0.875p pd=2.75u as=0.42p ps=1.84u w=1u l=0.28u
X2 VSS a_1315_24# a_1259_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.14p ps=1.28u w=1u l=0.28u
X3 a_1709_68# a_332_68# a_1315_24# VPW nfet_03v3 ad=0.625p pd=2.25u as=0.305p ps=1.61u w=1u l=0.28u
X4 a_2015_68# a_28_68# a_1709_68# VPW nfet_03v3 ad=0.43p pd=1.86u as=0.625p ps=2.25u w=1u l=0.28u
X5 a_332_68# a_28_68# VDD VNW pfet_03v3 ad=0.6693p pd=3.73u as=0.3588p ps=1.9u w=1.38u l=0.28u
X6 VSS CLK a_28_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X7 a_1259_68# a_332_68# a_853_68# VPW nfet_03v3 ad=0.14p pd=1.28u as=0.875p ps=2.75u w=1u l=0.28u
X8 VDD a_2187_24# a_2128_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.20355p ps=1.675u w=1.38u l=0.28u
X9 a_2187_24# a_1709_68# VSS VPW nfet_03v3 ad=0.55p pd=3.1u as=0.26p ps=1.52u w=1u l=0.28u
X10 VDD a_1315_24# a_1064_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.86595p ps=2.635u w=1.38u l=0.28u
X11 a_735_440# a_332_68# VDD VNW pfet_03v3 ad=0.2139p pd=1.69u as=1.3317p ps=4.69u w=1.38u l=0.285u
X12 a_853_68# D a_735_440# VNW pfet_03v3 ad=0.5313p pd=2.15u as=0.2139p ps=1.69u w=1.38u l=0.28u
X13 a_629_68# a_28_68# VSS VPW nfet_03v3 ad=0.42p pd=1.84u as=0.44p ps=2.88u w=1u l=0.28u
X14 VSS a_2187_24# Q VPW nfet_03v3 ad=0.615p pd=3.23u as=0.26p ps=1.52u w=1u l=0.28u
X15 VSS a_2187_24# a_2015_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.43p ps=1.86u w=1u l=0.28u
X16 a_1315_24# a_853_68# VDD VNW pfet_03v3 ad=0.83145p pd=2.585u as=0.3588p ps=1.9u w=1.38u l=0.28u
X17 Q a_2187_24# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X18 a_2187_24# a_1709_68# VDD VNW pfet_03v3 ad=0.759p pd=3.86u as=0.3588p ps=1.9u w=1.38u l=0.28u
X19 Q a_2187_24# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X20 a_1064_440# a_28_68# a_853_68# VNW pfet_03v3 ad=0.86595p pd=2.635u as=0.5313p ps=2.15u w=1.38u l=0.285u
X21 a_2128_440# a_332_68# a_1709_68# VNW pfet_03v3 ad=0.20355p pd=1.675u as=0.8418p ps=2.6u w=1.38u l=0.28u
X22 a_1315_24# a_853_68# VSS VPW nfet_03v3 ad=0.305p pd=1.61u as=0.26p ps=1.52u w=1u l=0.28u
X23 VDD a_2187_24# Q VNW pfet_03v3 ad=0.8487p pd=3.99u as=0.3588p ps=1.9u w=1.38u l=0.28u
X24 VDD CLK a_28_68# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X25 a_332_68# a_28_68# VSS VPW nfet_03v3 ad=0.485p pd=2.97u as=0.26p ps=1.52u w=1u l=0.28u
.ends

