magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 770 1486
<< nmos >>
rect 120 209 176 584
rect 280 209 336 584
rect 440 209 496 584
<< pmos >>
rect 120 776 176 1191
rect 280 776 336 1191
rect 440 776 496 1191
<< ndiff >>
rect 32 268 120 584
rect 32 222 45 268
rect 91 222 120 268
rect 32 209 120 222
rect 176 571 280 584
rect 176 325 205 571
rect 251 325 280 571
rect 176 209 280 325
rect 336 268 440 584
rect 336 222 365 268
rect 411 222 440 268
rect 336 209 440 222
rect 496 571 584 584
rect 496 325 525 571
rect 571 325 584 571
rect 496 209 584 325
<< pdiff >>
rect 32 1178 120 1191
rect 32 1132 45 1178
rect 91 1132 120 1178
rect 32 776 120 1132
rect 176 776 280 1191
rect 336 776 440 1191
rect 496 1055 584 1191
rect 496 809 525 1055
rect 571 809 584 1055
rect 496 776 584 809
<< ndiffc >>
rect 45 222 91 268
rect 205 325 251 571
rect 365 222 411 268
rect 525 325 571 571
<< pdiffc >>
rect 45 1132 91 1178
rect 525 809 571 1055
<< psubdiff >>
rect 28 87 656 100
rect 28 41 69 87
rect 615 41 656 87
rect 28 28 656 41
<< nsubdiff >>
rect 28 1359 656 1372
rect 28 1313 69 1359
rect 615 1313 656 1359
rect 28 1300 656 1313
<< psubdiffcont >>
rect 69 41 615 87
<< nsubdiffcont >>
rect 69 1313 615 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 120 716 176 776
rect 280 716 336 776
rect 440 716 496 776
rect 32 703 176 716
rect 32 657 45 703
rect 91 657 176 703
rect 32 644 176 657
rect 224 703 336 716
rect 224 657 237 703
rect 283 657 336 703
rect 224 644 336 657
rect 384 703 496 716
rect 384 657 397 703
rect 443 657 496 703
rect 384 644 496 657
rect 120 584 176 644
rect 280 584 336 644
rect 440 584 496 644
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
<< polycontact >>
rect 45 657 91 703
rect 237 657 283 703
rect 397 657 443 703
<< metal1 >>
rect 0 1359 684 1400
rect 0 1313 69 1359
rect 615 1313 684 1359
rect 0 1178 684 1313
rect 0 1132 45 1178
rect 91 1132 684 1178
rect 42 703 94 1086
rect 42 657 45 703
rect 91 657 94 703
rect 42 314 94 657
rect 234 703 286 1086
rect 234 657 237 703
rect 283 657 286 703
rect 234 628 286 657
rect 394 703 446 1086
rect 394 657 397 703
rect 443 657 446 703
rect 394 628 446 657
rect 522 1055 574 1086
rect 522 809 525 1055
rect 571 809 574 1055
rect 522 582 574 809
rect 205 571 574 582
rect 251 325 525 571
rect 571 325 574 571
rect 205 314 574 325
rect 0 222 45 268
rect 91 222 365 268
rect 411 222 684 268
rect 0 87 684 222
rect 0 41 69 87
rect 615 41 684 87
rect 0 0 684 41
<< labels >>
rlabel metal1 s 0 0 684 268 4 vss
port 3 nsew
rlabel metal1 s 0 1132 684 1400 4 vdd
port 5 nsew
rlabel metal1 s 522 314 574 1086 4 nq
port 7 nsew
rlabel metal1 s 42 314 94 1086 4 i0
port 9 nsew
rlabel metal1 s 234 628 286 1086 4 i1
port 11 nsew
rlabel metal1 s 394 628 446 1086 4 i2
port 13 nsew
<< end >>
