* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__buff_2.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__buff_2 VDD VNW VPW VSS A Y
X0 Y a_28_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X1 VSS A a_28_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X2 VDD a_28_68# Y VNW pfet_03v3 ad=1.0488p pd=4.28u as=0.3588p ps=1.9u w=1.38u l=0.28u
X3 VSS a_28_68# Y VPW nfet_03v3 ad=0.76p pd=3.52u as=0.26p ps=1.52u w=1u l=0.28u
X4 VDD A a_28_68# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X5 Y a_28_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

