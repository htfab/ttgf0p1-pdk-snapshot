* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__or2_4.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__or2_4 VDD VNW VPW VSS B A Y
X0 VSS a_28_440# Y VPW nfet_03v3 ad=0.6p pd=3.2u as=0.26p ps=1.52u w=1u l=0.28u
X1 VDD B a_172_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X2 Y a_28_440# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X3 a_28_440# A VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X4 Y a_28_440# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X5 Y a_28_440# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X6 VDD a_28_440# Y VNW pfet_03v3 ad=0.828p pd=3.96u as=0.3588p ps=1.9u w=1.38u l=0.28u
X7 VSS a_28_440# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X8 VDD a_28_440# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X9 Y a_28_440# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X10 a_172_440# A a_28_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X11 VSS B a_28_440# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

