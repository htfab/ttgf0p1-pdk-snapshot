magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 1226 1486
<< nmos >>
rect 120 209 176 452
rect 280 209 336 452
rect 440 209 496 452
rect 600 209 656 452
rect 760 209 816 452
<< pmos >>
rect 120 908 176 1191
rect 280 908 336 1191
rect 440 908 496 1191
rect 600 908 656 1191
rect 760 908 816 1191
<< ndiff >>
rect 32 405 120 452
rect 32 359 45 405
rect 91 359 120 405
rect 32 209 120 359
rect 176 268 280 452
rect 176 222 205 268
rect 251 222 280 268
rect 176 209 280 222
rect 336 405 440 452
rect 336 359 365 405
rect 411 359 440 405
rect 336 209 440 359
rect 496 268 600 452
rect 496 222 525 268
rect 571 222 600 268
rect 496 209 600 222
rect 656 405 760 452
rect 656 359 685 405
rect 731 359 760 405
rect 656 209 760 359
rect 816 268 904 452
rect 816 222 845 268
rect 891 222 904 268
rect 816 209 904 222
<< pdiff >>
rect 32 1071 120 1191
rect 32 925 45 1071
rect 91 925 120 1071
rect 32 908 120 925
rect 176 1178 280 1191
rect 176 1132 205 1178
rect 251 1132 280 1178
rect 176 908 280 1132
rect 336 1071 440 1191
rect 336 925 365 1071
rect 411 925 440 1071
rect 336 908 440 925
rect 496 1178 600 1191
rect 496 1132 525 1178
rect 571 1132 600 1178
rect 496 908 600 1132
rect 656 1071 760 1191
rect 656 925 685 1071
rect 731 925 760 1071
rect 656 908 760 925
rect 816 1178 904 1191
rect 816 1132 845 1178
rect 891 1132 904 1178
rect 816 908 904 1132
<< ndiffc >>
rect 45 359 91 405
rect 205 222 251 268
rect 365 359 411 405
rect 525 222 571 268
rect 685 359 731 405
rect 845 222 891 268
<< pdiffc >>
rect 45 925 91 1071
rect 205 1132 251 1178
rect 365 925 411 1071
rect 525 1132 571 1178
rect 685 925 731 1071
rect 845 1132 891 1178
<< psubdiff >>
rect 28 87 1112 100
rect 28 41 47 87
rect 1093 41 1112 87
rect 28 28 1112 41
<< nsubdiff >>
rect 28 1359 1112 1372
rect 28 1313 47 1359
rect 1093 1313 1112 1359
rect 28 1300 1112 1313
<< psubdiffcont >>
rect 47 41 1093 87
<< nsubdiffcont >>
rect 47 1313 1093 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 600 1191 656 1235
rect 760 1191 816 1235
rect 120 848 176 908
rect 120 835 202 848
rect 120 789 143 835
rect 189 789 202 835
rect 120 776 202 789
rect 280 716 336 908
rect 440 716 496 908
rect 600 716 656 908
rect 760 716 816 908
rect 32 703 816 716
rect 32 657 45 703
rect 91 657 816 703
rect 32 644 816 657
rect 120 571 202 584
rect 120 525 143 571
rect 189 525 202 571
rect 120 512 202 525
rect 120 452 176 512
rect 280 452 336 644
rect 440 452 496 644
rect 600 452 656 644
rect 760 452 816 644
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
rect 600 165 656 209
rect 760 165 816 209
<< polycontact >>
rect 143 789 189 835
rect 45 657 91 703
rect 143 525 189 571
<< metal1 >>
rect 0 1359 1140 1400
rect 0 1313 47 1359
rect 1093 1313 1140 1359
rect 0 1178 1140 1313
rect 0 1132 205 1178
rect 251 1132 525 1178
rect 571 1132 845 1178
rect 891 1132 1140 1178
rect 45 1071 91 1086
rect 42 925 45 982
rect 91 925 94 982
rect 42 703 94 925
rect 42 657 45 703
rect 91 657 94 703
rect 42 405 94 657
rect 42 359 45 405
rect 91 359 94 405
rect 42 348 94 359
rect 140 835 192 1086
rect 140 789 143 835
rect 189 789 192 835
rect 140 571 192 789
rect 140 525 143 571
rect 189 525 192 571
rect 45 314 91 348
rect 140 314 192 525
rect 362 1071 414 1086
rect 362 925 365 1071
rect 411 925 414 1071
rect 685 1071 731 1086
rect 362 714 414 925
rect 682 925 685 982
rect 731 925 734 982
rect 682 714 734 925
rect 362 646 734 714
rect 362 405 414 646
rect 362 359 365 405
rect 411 359 414 405
rect 362 314 414 359
rect 682 405 734 646
rect 682 359 685 405
rect 731 359 734 405
rect 682 348 734 359
rect 685 314 731 348
rect 0 222 205 268
rect 251 222 525 268
rect 571 222 845 268
rect 891 222 1140 268
rect 0 87 1140 222
rect 0 41 47 87
rect 1093 41 1140 87
rect 0 0 1140 41
<< labels >>
rlabel metal1 s 0 1132 1140 1400 4 vdd
port 3 nsew
rlabel metal1 s 0 0 1140 268 4 vss
port 5 nsew
rlabel metal1 s 140 314 192 1086 4 i
port 7 nsew
rlabel metal1 s 362 314 414 1086 4 q
port 9 nsew
<< end >>
