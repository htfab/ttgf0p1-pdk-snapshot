* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__fill_4.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__fill_4 VDD VNW VPW VSS
.ends

