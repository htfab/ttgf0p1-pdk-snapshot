magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect 5889 11760 13827 16428
rect 8785 9699 9384 9700
rect 13054 9699 13654 9700
rect 6493 7883 7347 7884
rect 4800 7122 5430 7790
rect 6493 7707 7861 7883
rect 6540 7412 7861 7707
rect 6493 7410 7861 7412
rect 6493 7185 7860 7410
rect 542 6727 5430 7122
rect 6234 6972 7860 7185
rect 542 6338 5654 6727
rect 4800 5991 5654 6338
rect 6234 6235 7861 6972
rect 6234 5995 7860 6235
rect 8785 5491 13654 9699
rect 9270 5490 13654 5491
rect 9271 5152 13654 5490
rect 10470 4675 13654 5152
rect 10470 4518 13057 4675
rect -73 2245 8748 3429
rect 7919 852 8748 2245
rect 7137 -1400 8748 852
<< mvnmos >>
rect 6700 9039 6820 11035
rect 6924 9039 7044 11035
rect 7148 9039 7268 11035
rect 7372 9039 7492 11035
rect 7596 9039 7716 11035
rect 8937 9839 9057 11313
rect 9161 9839 9281 11313
rect 9385 9839 9505 11313
rect 9609 9839 9729 11313
rect 9833 9839 9953 11313
rect 10057 9839 10177 11313
rect 10281 9839 10401 11313
rect 10505 9839 10625 11313
rect 10729 9839 10849 11313
rect 10953 9839 11073 11313
rect 11177 9839 11297 11313
rect 11401 9839 11521 11313
rect 11625 9839 11745 11313
rect 11849 9839 11969 11313
rect 12073 9839 12193 11313
rect 12297 9839 12417 11313
rect 12521 9839 12641 11313
rect 12745 9839 12865 11313
rect 12969 9839 13089 11313
rect 13193 9839 13313 11313
rect 5055 7941 5175 8133
rect 6972 8021 7092 8213
rect 7486 8021 7606 8213
rect 5055 5402 5175 5674
rect 5279 5402 5399 5674
rect 6748 5402 6868 5856
rect 6972 5402 7092 5856
rect 7486 5402 7606 5856
rect 5157 3772 5397 3892
rect 6235 3772 6475 3892
rect 6954 3777 7154 3897
rect 7600 3790 7720 3940
rect 8114 3789 8234 4393
rect 9526 262 9646 4798
rect 9750 262 9870 4798
rect 9974 262 10094 4798
rect 10725 484 10845 4113
rect 10949 484 11069 4113
rect 11173 484 11293 4113
rect 11397 484 11517 4113
rect 12010 3205 12130 4113
rect 12233 3205 12353 4113
rect 12458 3205 12578 4113
rect 12681 3205 12801 4113
<< mvpmos >>
rect 6408 13461 6528 15957
rect 6632 13461 6752 15957
rect 6856 13461 6976 15957
rect 7080 13461 7200 15957
rect 7304 13461 7424 15957
rect 7528 13461 7648 15957
rect 7752 13461 7872 15957
rect 7976 13461 8096 15957
rect 8200 13461 8320 15957
rect 8424 13461 8544 15957
rect 8937 12283 9057 15957
rect 9161 12283 9281 15957
rect 9385 12283 9505 15957
rect 9609 12283 9729 15957
rect 9833 12283 9953 15957
rect 10057 12283 10177 15957
rect 10281 12283 10401 15957
rect 10505 12283 10625 15957
rect 10729 12283 10849 15957
rect 10953 12283 11073 15957
rect 11177 12283 11297 15957
rect 11401 12283 11521 15957
rect 11625 12283 11745 15957
rect 11849 12283 11969 15957
rect 12073 12283 12193 15957
rect 12297 12283 12417 15957
rect 12521 12283 12641 15957
rect 12745 12283 12865 15957
rect 12969 12283 13089 15957
rect 13193 12283 13313 15957
rect 5055 7195 5175 7649
rect 6748 7514 6868 7742
rect 6972 7514 7092 7742
rect 7486 7550 7606 7742
rect 5055 6131 5174 6587
rect 5279 6131 5398 6587
rect 6748 6137 6868 7271
rect 6972 6137 7092 7271
rect 7486 6377 7606 6831
rect 9526 5293 9646 9193
rect 9750 5293 9870 9193
rect 9974 5293 10094 9193
rect 5157 3080 5397 3260
rect 6235 3080 6475 3260
rect 6954 3080 7154 3260
rect 7600 2882 7720 3260
rect 8114 2506 8234 3260
rect 8338 2506 8458 3260
rect 10725 4659 10845 9195
rect 10949 4659 11069 9195
rect 11173 4659 11293 9195
rect 11397 4659 11517 9195
rect 12010 4659 12130 9195
rect 12234 4659 12354 9195
rect 12458 4659 12578 9195
rect 12682 4659 12802 9195
<< mvndiff >>
rect 6612 11022 6700 11035
rect 6612 9052 6625 11022
rect 6671 9052 6700 11022
rect 6612 9039 6700 9052
rect 6820 11022 6924 11035
rect 6820 9052 6849 11022
rect 6895 9052 6924 11022
rect 6820 9039 6924 9052
rect 7044 11022 7148 11035
rect 7044 9052 7073 11022
rect 7119 9052 7148 11022
rect 7044 9039 7148 9052
rect 7268 11022 7372 11035
rect 7268 9052 7297 11022
rect 7343 9052 7372 11022
rect 7268 9039 7372 9052
rect 7492 11022 7596 11035
rect 7492 9052 7521 11022
rect 7567 9052 7596 11022
rect 7492 9039 7596 9052
rect 7716 11022 7804 11035
rect 7716 9052 7745 11022
rect 7791 9052 7804 11022
rect 7716 9039 7804 9052
rect 8849 11300 8937 11313
rect 8849 9852 8862 11300
rect 8908 9852 8937 11300
rect 8849 9839 8937 9852
rect 9057 11300 9161 11313
rect 9057 9852 9086 11300
rect 9132 9852 9161 11300
rect 9057 9839 9161 9852
rect 9281 11300 9385 11313
rect 9281 9852 9310 11300
rect 9356 9852 9385 11300
rect 9281 9839 9385 9852
rect 9505 11300 9609 11313
rect 9505 9852 9534 11300
rect 9580 9852 9609 11300
rect 9505 9839 9609 9852
rect 9729 11300 9833 11313
rect 9729 9852 9758 11300
rect 9804 9852 9833 11300
rect 9729 9839 9833 9852
rect 9953 11300 10057 11313
rect 9953 9852 9982 11300
rect 10028 9852 10057 11300
rect 9953 9839 10057 9852
rect 10177 11300 10281 11313
rect 10177 9852 10206 11300
rect 10252 9852 10281 11300
rect 10177 9839 10281 9852
rect 10401 11300 10505 11313
rect 10401 9852 10430 11300
rect 10476 9852 10505 11300
rect 10401 9839 10505 9852
rect 10625 11300 10729 11313
rect 10625 9852 10654 11300
rect 10700 9852 10729 11300
rect 10625 9839 10729 9852
rect 10849 11300 10953 11313
rect 10849 9852 10878 11300
rect 10924 9852 10953 11300
rect 10849 9839 10953 9852
rect 11073 11300 11177 11313
rect 11073 9852 11102 11300
rect 11148 9852 11177 11300
rect 11073 9839 11177 9852
rect 11297 11300 11401 11313
rect 11297 9852 11326 11300
rect 11372 9852 11401 11300
rect 11297 9839 11401 9852
rect 11521 11300 11625 11313
rect 11521 9852 11550 11300
rect 11596 9852 11625 11300
rect 11521 9839 11625 9852
rect 11745 11300 11849 11313
rect 11745 9852 11774 11300
rect 11820 9852 11849 11300
rect 11745 9839 11849 9852
rect 11969 11300 12073 11313
rect 11969 9852 11998 11300
rect 12044 9852 12073 11300
rect 11969 9839 12073 9852
rect 12193 11300 12297 11313
rect 12193 9852 12222 11300
rect 12268 9852 12297 11300
rect 12193 9839 12297 9852
rect 12417 11300 12521 11313
rect 12417 9852 12446 11300
rect 12492 9852 12521 11300
rect 12417 9839 12521 9852
rect 12641 11300 12745 11313
rect 12641 9852 12670 11300
rect 12716 9852 12745 11300
rect 12641 9839 12745 9852
rect 12865 11300 12969 11313
rect 12865 9852 12894 11300
rect 12940 9852 12969 11300
rect 12865 9839 12969 9852
rect 13089 11300 13193 11313
rect 13089 9852 13118 11300
rect 13164 9852 13193 11300
rect 13089 9839 13193 9852
rect 13313 11300 13401 11313
rect 13313 9852 13342 11300
rect 13388 9852 13401 11300
rect 13313 9839 13401 9852
rect 6884 8200 6972 8213
rect 6884 8154 6897 8200
rect 6943 8154 6972 8200
rect 4967 8120 5055 8133
rect 4967 8074 4980 8120
rect 5026 8074 5055 8120
rect 4967 8000 5055 8074
rect 4967 7954 4980 8000
rect 5026 7954 5055 8000
rect 4967 7941 5055 7954
rect 5175 8120 5263 8133
rect 5175 8074 5204 8120
rect 5250 8074 5263 8120
rect 5175 8000 5263 8074
rect 6884 8080 6972 8154
rect 6884 8034 6897 8080
rect 6943 8034 6972 8080
rect 6884 8021 6972 8034
rect 7092 8200 7180 8213
rect 7092 8154 7121 8200
rect 7167 8154 7180 8200
rect 7092 8080 7180 8154
rect 7092 8034 7121 8080
rect 7167 8034 7180 8080
rect 7092 8021 7180 8034
rect 7398 8200 7486 8213
rect 7398 8154 7411 8200
rect 7457 8154 7486 8200
rect 7398 8080 7486 8154
rect 7398 8034 7411 8080
rect 7457 8034 7486 8080
rect 7398 8021 7486 8034
rect 7606 8200 7694 8213
rect 7606 8154 7635 8200
rect 7681 8154 7694 8200
rect 7606 8080 7694 8154
rect 7606 8034 7635 8080
rect 7681 8034 7694 8080
rect 7606 8021 7694 8034
rect 5175 7954 5204 8000
rect 5250 7954 5263 8000
rect 5175 7941 5263 7954
rect 6660 5843 6748 5856
rect 6660 5797 6673 5843
rect 6719 5797 6748 5843
rect 4967 5661 5055 5674
rect 4967 5415 4980 5661
rect 5026 5415 5055 5661
rect 4967 5402 5055 5415
rect 5175 5661 5279 5674
rect 5175 5415 5204 5661
rect 5250 5415 5279 5661
rect 5175 5402 5279 5415
rect 5399 5661 5487 5674
rect 5399 5415 5428 5661
rect 5474 5415 5487 5661
rect 5399 5402 5487 5415
rect 6660 5716 6748 5797
rect 6660 5670 6673 5716
rect 6719 5670 6748 5716
rect 6660 5589 6748 5670
rect 6660 5543 6673 5589
rect 6719 5543 6748 5589
rect 6660 5461 6748 5543
rect 6660 5415 6673 5461
rect 6719 5415 6748 5461
rect 6660 5402 6748 5415
rect 6868 5843 6972 5856
rect 6868 5797 6897 5843
rect 6943 5797 6972 5843
rect 6868 5716 6972 5797
rect 6868 5670 6897 5716
rect 6943 5670 6972 5716
rect 6868 5589 6972 5670
rect 6868 5543 6897 5589
rect 6943 5543 6972 5589
rect 6868 5461 6972 5543
rect 6868 5415 6897 5461
rect 6943 5415 6972 5461
rect 6868 5402 6972 5415
rect 7092 5843 7180 5856
rect 7092 5797 7121 5843
rect 7167 5797 7180 5843
rect 7092 5716 7180 5797
rect 7092 5670 7121 5716
rect 7167 5670 7180 5716
rect 7092 5589 7180 5670
rect 7092 5543 7121 5589
rect 7167 5543 7180 5589
rect 7092 5461 7180 5543
rect 7092 5415 7121 5461
rect 7167 5415 7180 5461
rect 7092 5402 7180 5415
rect 7398 5843 7486 5856
rect 7398 5797 7411 5843
rect 7457 5797 7486 5843
rect 7398 5716 7486 5797
rect 7398 5670 7411 5716
rect 7457 5670 7486 5716
rect 7398 5589 7486 5670
rect 7398 5543 7411 5589
rect 7457 5543 7486 5589
rect 7398 5461 7486 5543
rect 7398 5415 7411 5461
rect 7457 5415 7486 5461
rect 7398 5402 7486 5415
rect 7606 5843 7694 5856
rect 7606 5797 7635 5843
rect 7681 5797 7694 5843
rect 7606 5716 7694 5797
rect 7606 5670 7635 5716
rect 7681 5670 7694 5716
rect 7606 5589 7694 5670
rect 7606 5543 7635 5589
rect 7681 5543 7694 5589
rect 7606 5461 7694 5543
rect 7606 5415 7635 5461
rect 7681 5415 7694 5461
rect 7606 5402 7694 5415
rect 8026 4380 8114 4393
rect 8026 4334 8039 4380
rect 8085 4334 8114 4380
rect 8026 4273 8114 4334
rect 8026 4227 8039 4273
rect 8085 4227 8114 4273
rect 8026 4166 8114 4227
rect 8026 4120 8039 4166
rect 8085 4120 8114 4166
rect 8026 4060 8114 4120
rect 8026 4014 8039 4060
rect 8085 4014 8114 4060
rect 8026 3954 8114 4014
rect 5069 3855 5157 3892
rect 5069 3809 5082 3855
rect 5128 3809 5157 3855
rect 5069 3772 5157 3809
rect 5397 3855 5485 3892
rect 5397 3809 5426 3855
rect 5472 3809 5485 3855
rect 5397 3772 5485 3809
rect 6147 3855 6235 3892
rect 6147 3809 6160 3855
rect 6206 3809 6235 3855
rect 6147 3772 6235 3809
rect 6475 3855 6563 3892
rect 6475 3809 6504 3855
rect 6550 3809 6563 3855
rect 6475 3772 6563 3809
rect 6866 3860 6954 3897
rect 6866 3814 6879 3860
rect 6925 3814 6954 3860
rect 6866 3777 6954 3814
rect 7154 3860 7242 3897
rect 7154 3814 7183 3860
rect 7229 3814 7242 3860
rect 7154 3777 7242 3814
rect 7512 3888 7600 3940
rect 7512 3842 7525 3888
rect 7571 3842 7600 3888
rect 7512 3790 7600 3842
rect 7720 3888 7808 3940
rect 7720 3842 7749 3888
rect 7795 3842 7808 3888
rect 7720 3790 7808 3842
rect 8026 3908 8039 3954
rect 8085 3908 8114 3954
rect 8026 3848 8114 3908
rect 8026 3802 8039 3848
rect 8085 3802 8114 3848
rect 8026 3789 8114 3802
rect 8234 4380 8322 4393
rect 8234 4334 8263 4380
rect 8309 4334 8322 4380
rect 8234 4273 8322 4334
rect 8234 4227 8263 4273
rect 8309 4227 8322 4273
rect 8234 4166 8322 4227
rect 8234 4120 8263 4166
rect 8309 4120 8322 4166
rect 8234 4060 8322 4120
rect 8234 4014 8263 4060
rect 8309 4014 8322 4060
rect 8234 3954 8322 4014
rect 8234 3908 8263 3954
rect 8309 3908 8322 3954
rect 8234 3848 8322 3908
rect 8234 3802 8263 3848
rect 8309 3802 8322 3848
rect 8234 3789 8322 3802
rect 9407 4752 9526 4798
rect 9407 4706 9451 4752
rect 9497 4706 9526 4752
rect 9407 4584 9526 4706
rect 9407 4538 9451 4584
rect 9497 4538 9526 4584
rect 9407 4417 9526 4538
rect 9407 4371 9451 4417
rect 9497 4371 9526 4417
rect 9407 4249 9526 4371
rect 9407 4203 9451 4249
rect 9497 4203 9526 4249
rect 9407 4081 9526 4203
rect 9407 4035 9451 4081
rect 9497 4035 9526 4081
rect 9407 3913 9526 4035
rect 9407 3867 9451 3913
rect 9497 3867 9526 3913
rect 9407 3746 9526 3867
rect 9407 3700 9451 3746
rect 9497 3700 9526 3746
rect 9407 3578 9526 3700
rect 9407 3532 9451 3578
rect 9497 3532 9526 3578
rect 9407 3410 9526 3532
rect 9407 3364 9451 3410
rect 9497 3364 9526 3410
rect 9407 3242 9526 3364
rect 9407 3196 9451 3242
rect 9497 3196 9526 3242
rect 9407 3075 9526 3196
rect 9407 3029 9451 3075
rect 9497 3029 9526 3075
rect 9407 2905 9526 3029
rect 9407 2859 9451 2905
rect 9497 2859 9526 2905
rect 9407 2735 9526 2859
rect 9407 2689 9451 2735
rect 9497 2689 9526 2735
rect 9407 2565 9526 2689
rect 9407 2519 9451 2565
rect 9497 2519 9526 2565
rect 9407 2395 9526 2519
rect 9407 2349 9451 2395
rect 9497 2349 9526 2395
rect 9407 2225 9526 2349
rect 9407 2179 9451 2225
rect 9497 2179 9526 2225
rect 9407 2055 9526 2179
rect 9407 2009 9451 2055
rect 9497 2009 9526 2055
rect 9407 1884 9526 2009
rect 9407 1838 9451 1884
rect 9497 1838 9526 1884
rect 9407 1714 9526 1838
rect 9407 1668 9451 1714
rect 9497 1668 9526 1714
rect 9407 1544 9526 1668
rect 9407 1498 9451 1544
rect 9497 1498 9526 1544
rect 9407 1374 9526 1498
rect 9407 1328 9451 1374
rect 9497 1328 9526 1374
rect 9407 1204 9526 1328
rect 9407 1158 9451 1204
rect 9497 1158 9526 1204
rect 9407 1034 9526 1158
rect 9407 988 9451 1034
rect 9497 988 9526 1034
rect 9407 864 9526 988
rect 9407 818 9451 864
rect 9497 818 9526 864
rect 9407 694 9526 818
rect 9407 648 9451 694
rect 9497 648 9526 694
rect 9407 524 9526 648
rect 9407 478 9451 524
rect 9497 478 9526 524
rect 9407 354 9526 478
rect 9407 308 9451 354
rect 9497 308 9526 354
rect 9407 262 9526 308
rect 9646 262 9750 4798
rect 9870 262 9974 4798
rect 10094 4584 10212 4798
rect 10094 4538 10123 4584
rect 10169 4538 10212 4584
rect 10094 4417 10212 4538
rect 10094 4371 10123 4417
rect 10169 4371 10212 4417
rect 10094 4249 10212 4371
rect 10094 4203 10123 4249
rect 10169 4203 10212 4249
rect 10094 4081 10212 4203
rect 10094 4035 10123 4081
rect 10169 4035 10212 4081
rect 10094 3913 10212 4035
rect 10094 3867 10123 3913
rect 10169 3867 10212 3913
rect 10094 3746 10212 3867
rect 10094 3700 10123 3746
rect 10169 3700 10212 3746
rect 10094 3578 10212 3700
rect 10094 3532 10123 3578
rect 10169 3532 10212 3578
rect 10094 3410 10212 3532
rect 10094 3364 10123 3410
rect 10169 3364 10212 3410
rect 10094 3242 10212 3364
rect 10094 3196 10123 3242
rect 10169 3196 10212 3242
rect 10094 3075 10212 3196
rect 10094 3029 10123 3075
rect 10169 3029 10212 3075
rect 10094 2905 10212 3029
rect 10094 2859 10123 2905
rect 10169 2859 10212 2905
rect 10094 2735 10212 2859
rect 10094 2689 10123 2735
rect 10169 2689 10212 2735
rect 10094 2565 10212 2689
rect 10094 2519 10123 2565
rect 10169 2519 10212 2565
rect 10094 2395 10212 2519
rect 10094 2349 10123 2395
rect 10169 2349 10212 2395
rect 10094 2225 10212 2349
rect 10094 2179 10123 2225
rect 10169 2179 10212 2225
rect 10094 2055 10212 2179
rect 10094 2009 10123 2055
rect 10169 2009 10212 2055
rect 10094 1884 10212 2009
rect 10094 1838 10123 1884
rect 10169 1838 10212 1884
rect 10094 1714 10212 1838
rect 10094 1668 10123 1714
rect 10169 1668 10212 1714
rect 10094 1544 10212 1668
rect 10094 1498 10123 1544
rect 10169 1498 10212 1544
rect 10094 1374 10212 1498
rect 10094 1328 10123 1374
rect 10169 1328 10212 1374
rect 10094 1204 10212 1328
rect 10094 1158 10123 1204
rect 10169 1158 10212 1204
rect 10094 1034 10212 1158
rect 10094 988 10123 1034
rect 10169 988 10212 1034
rect 10094 864 10212 988
rect 10094 818 10123 864
rect 10169 818 10212 864
rect 10094 694 10212 818
rect 10094 648 10123 694
rect 10169 648 10212 694
rect 10094 524 10212 648
rect 10094 478 10123 524
rect 10169 478 10212 524
rect 10606 4068 10725 4113
rect 10606 4022 10650 4068
rect 10696 4022 10725 4068
rect 10606 3900 10725 4022
rect 10606 3854 10650 3900
rect 10696 3854 10725 3900
rect 10606 3732 10725 3854
rect 10606 3686 10650 3732
rect 10696 3686 10725 3732
rect 10606 3564 10725 3686
rect 10606 3518 10650 3564
rect 10696 3518 10725 3564
rect 10606 3397 10725 3518
rect 10606 3351 10650 3397
rect 10696 3351 10725 3397
rect 10606 3229 10725 3351
rect 10606 3183 10650 3229
rect 10696 3183 10725 3229
rect 10606 3061 10725 3183
rect 10606 3015 10650 3061
rect 10696 3015 10725 3061
rect 10606 2893 10725 3015
rect 10606 2847 10650 2893
rect 10696 2847 10725 2893
rect 10606 2726 10725 2847
rect 10606 2680 10650 2726
rect 10696 2680 10725 2726
rect 10606 2558 10725 2680
rect 10606 2512 10650 2558
rect 10696 2512 10725 2558
rect 10606 2390 10725 2512
rect 10606 2344 10650 2390
rect 10696 2344 10725 2390
rect 10606 2220 10725 2344
rect 10606 2174 10650 2220
rect 10696 2174 10725 2220
rect 10606 2050 10725 2174
rect 10606 2004 10650 2050
rect 10696 2004 10725 2050
rect 10606 1880 10725 2004
rect 10606 1834 10650 1880
rect 10696 1834 10725 1880
rect 10606 1710 10725 1834
rect 10606 1664 10650 1710
rect 10696 1664 10725 1710
rect 10606 1540 10725 1664
rect 10606 1494 10650 1540
rect 10696 1494 10725 1540
rect 10606 1370 10725 1494
rect 10606 1324 10650 1370
rect 10696 1324 10725 1370
rect 10606 1200 10725 1324
rect 10606 1154 10650 1200
rect 10696 1154 10725 1200
rect 10606 1030 10725 1154
rect 10606 984 10650 1030
rect 10696 984 10725 1030
rect 10606 860 10725 984
rect 10606 814 10650 860
rect 10696 814 10725 860
rect 10606 690 10725 814
rect 10606 644 10650 690
rect 10696 644 10725 690
rect 10606 484 10725 644
rect 10845 484 10949 4113
rect 11069 4068 11173 4113
rect 11069 4022 11098 4068
rect 11144 4022 11173 4068
rect 11069 3900 11173 4022
rect 11069 3854 11098 3900
rect 11144 3854 11173 3900
rect 11069 3732 11173 3854
rect 11069 3686 11098 3732
rect 11144 3686 11173 3732
rect 11069 3564 11173 3686
rect 11069 3518 11098 3564
rect 11144 3518 11173 3564
rect 11069 3397 11173 3518
rect 11069 3351 11098 3397
rect 11144 3351 11173 3397
rect 11069 3229 11173 3351
rect 11069 3183 11098 3229
rect 11144 3183 11173 3229
rect 11069 3061 11173 3183
rect 11069 3015 11098 3061
rect 11144 3015 11173 3061
rect 11069 2893 11173 3015
rect 11069 2847 11098 2893
rect 11144 2847 11173 2893
rect 11069 2726 11173 2847
rect 11069 2680 11098 2726
rect 11144 2680 11173 2726
rect 11069 2558 11173 2680
rect 11069 2512 11098 2558
rect 11144 2512 11173 2558
rect 11069 2390 11173 2512
rect 11069 2344 11098 2390
rect 11144 2344 11173 2390
rect 11069 2220 11173 2344
rect 11069 2174 11098 2220
rect 11144 2174 11173 2220
rect 11069 2050 11173 2174
rect 11069 2004 11098 2050
rect 11144 2004 11173 2050
rect 11069 1880 11173 2004
rect 11069 1834 11098 1880
rect 11144 1834 11173 1880
rect 11069 1710 11173 1834
rect 11069 1664 11098 1710
rect 11144 1664 11173 1710
rect 11069 1540 11173 1664
rect 11069 1494 11098 1540
rect 11144 1494 11173 1540
rect 11069 1370 11173 1494
rect 11069 1324 11098 1370
rect 11144 1324 11173 1370
rect 11069 1200 11173 1324
rect 11069 1154 11098 1200
rect 11144 1154 11173 1200
rect 11069 1030 11173 1154
rect 11069 984 11098 1030
rect 11144 984 11173 1030
rect 11069 860 11173 984
rect 11069 814 11098 860
rect 11144 814 11173 860
rect 11069 690 11173 814
rect 11069 644 11098 690
rect 11144 644 11173 690
rect 11069 484 11173 644
rect 11293 484 11397 4113
rect 11517 4068 11635 4113
rect 11517 4022 11546 4068
rect 11592 4022 11635 4068
rect 11517 3900 11635 4022
rect 11517 3854 11546 3900
rect 11592 3854 11635 3900
rect 11517 3732 11635 3854
rect 11517 3686 11546 3732
rect 11592 3686 11635 3732
rect 11517 3564 11635 3686
rect 11517 3518 11546 3564
rect 11592 3518 11635 3564
rect 11517 3397 11635 3518
rect 11517 3351 11546 3397
rect 11592 3351 11635 3397
rect 11517 3229 11635 3351
rect 11517 3183 11546 3229
rect 11592 3183 11635 3229
rect 11891 4068 12010 4113
rect 11891 4022 11934 4068
rect 11980 4022 12010 4068
rect 11891 3900 12010 4022
rect 11891 3854 11934 3900
rect 11980 3854 12010 3900
rect 11891 3732 12010 3854
rect 11891 3686 11934 3732
rect 11980 3686 12010 3732
rect 11891 3564 12010 3686
rect 11891 3518 11934 3564
rect 11980 3518 12010 3564
rect 11891 3397 12010 3518
rect 11891 3351 11934 3397
rect 11980 3351 12010 3397
rect 11891 3205 12010 3351
rect 12130 3205 12233 4113
rect 12353 4068 12458 4113
rect 12353 4022 12382 4068
rect 12428 4022 12458 4068
rect 12353 3900 12458 4022
rect 12353 3854 12382 3900
rect 12428 3854 12458 3900
rect 12353 3732 12458 3854
rect 12353 3686 12382 3732
rect 12428 3686 12458 3732
rect 12353 3564 12458 3686
rect 12353 3518 12382 3564
rect 12428 3518 12458 3564
rect 12353 3397 12458 3518
rect 12353 3351 12382 3397
rect 12428 3351 12458 3397
rect 12353 3205 12458 3351
rect 12578 3205 12681 4113
rect 12801 4068 12920 4113
rect 12801 4022 12830 4068
rect 12876 4022 12920 4068
rect 12801 3732 12920 4022
rect 12801 3686 12830 3732
rect 12876 3686 12920 3732
rect 12801 3564 12920 3686
rect 12801 3518 12830 3564
rect 12876 3518 12920 3564
rect 12801 3397 12920 3518
rect 12801 3351 12830 3397
rect 12876 3351 12920 3397
rect 12801 3205 12920 3351
rect 11517 3061 11635 3183
rect 11517 3015 11546 3061
rect 11592 3015 11635 3061
rect 11517 2893 11635 3015
rect 11517 2847 11546 2893
rect 11592 2847 11635 2893
rect 11517 2726 11635 2847
rect 11517 2680 11546 2726
rect 11592 2680 11635 2726
rect 11517 2558 11635 2680
rect 11517 2512 11546 2558
rect 11592 2512 11635 2558
rect 11517 2390 11635 2512
rect 11517 2344 11546 2390
rect 11592 2344 11635 2390
rect 11517 2220 11635 2344
rect 11517 2174 11546 2220
rect 11592 2174 11635 2220
rect 11517 2050 11635 2174
rect 11517 2004 11546 2050
rect 11592 2004 11635 2050
rect 11517 1880 11635 2004
rect 11517 1834 11546 1880
rect 11592 1834 11635 1880
rect 11517 1710 11635 1834
rect 11517 1664 11546 1710
rect 11592 1664 11635 1710
rect 11517 1540 11635 1664
rect 11517 1494 11546 1540
rect 11592 1494 11635 1540
rect 11517 1370 11635 1494
rect 11517 1324 11546 1370
rect 11592 1324 11635 1370
rect 11517 1200 11635 1324
rect 11517 1154 11546 1200
rect 11592 1154 11635 1200
rect 11517 1030 11635 1154
rect 11517 984 11546 1030
rect 11592 984 11635 1030
rect 11517 860 11635 984
rect 11517 814 11546 860
rect 11592 814 11635 860
rect 11517 690 11635 814
rect 11517 644 11546 690
rect 11592 644 11635 690
rect 11517 484 11635 644
rect 10094 354 10212 478
rect 10094 308 10123 354
rect 10169 308 10212 354
rect 10094 262 10212 308
<< mvpdiff >>
rect 6320 15944 6408 15957
rect 6320 13474 6333 15944
rect 6379 13474 6408 15944
rect 6320 13461 6408 13474
rect 6528 15944 6632 15957
rect 6528 13474 6557 15944
rect 6603 13474 6632 15944
rect 6528 13461 6632 13474
rect 6752 15944 6856 15957
rect 6752 13474 6781 15944
rect 6827 13474 6856 15944
rect 6752 13461 6856 13474
rect 6976 15944 7080 15957
rect 6976 13474 7005 15944
rect 7051 13474 7080 15944
rect 6976 13461 7080 13474
rect 7200 15944 7304 15957
rect 7200 13474 7229 15944
rect 7275 13474 7304 15944
rect 7200 13461 7304 13474
rect 7424 15944 7528 15957
rect 7424 13474 7453 15944
rect 7499 13474 7528 15944
rect 7424 13461 7528 13474
rect 7648 15944 7752 15957
rect 7648 13474 7677 15944
rect 7723 13474 7752 15944
rect 7648 13461 7752 13474
rect 7872 15944 7976 15957
rect 7872 13474 7901 15944
rect 7947 13474 7976 15944
rect 7872 13461 7976 13474
rect 8096 15944 8200 15957
rect 8096 13474 8125 15944
rect 8171 13474 8200 15944
rect 8096 13461 8200 13474
rect 8320 15944 8424 15957
rect 8320 13474 8349 15944
rect 8395 13474 8424 15944
rect 8320 13461 8424 13474
rect 8544 15944 8632 15957
rect 8544 13474 8573 15944
rect 8619 13474 8632 15944
rect 8544 13461 8632 13474
rect 8849 15944 8937 15957
rect 8849 12296 8862 15944
rect 8908 12296 8937 15944
rect 8849 12283 8937 12296
rect 9057 15944 9161 15957
rect 9057 12296 9086 15944
rect 9132 12296 9161 15944
rect 9057 12283 9161 12296
rect 9281 15944 9385 15957
rect 9281 12296 9310 15944
rect 9356 12296 9385 15944
rect 9281 12283 9385 12296
rect 9505 15944 9609 15957
rect 9505 12296 9534 15944
rect 9580 12296 9609 15944
rect 9505 12283 9609 12296
rect 9729 15944 9833 15957
rect 9729 12296 9758 15944
rect 9804 12296 9833 15944
rect 9729 12283 9833 12296
rect 9953 15944 10057 15957
rect 9953 12296 9982 15944
rect 10028 12296 10057 15944
rect 9953 12283 10057 12296
rect 10177 15944 10281 15957
rect 10177 12296 10206 15944
rect 10252 12296 10281 15944
rect 10177 12283 10281 12296
rect 10401 15944 10505 15957
rect 10401 12296 10430 15944
rect 10476 12296 10505 15944
rect 10401 12283 10505 12296
rect 10625 15944 10729 15957
rect 10625 12296 10654 15944
rect 10700 12296 10729 15944
rect 10625 12283 10729 12296
rect 10849 15944 10953 15957
rect 10849 12296 10878 15944
rect 10924 12296 10953 15944
rect 10849 12283 10953 12296
rect 11073 15944 11177 15957
rect 11073 12296 11102 15944
rect 11148 12296 11177 15944
rect 11073 12283 11177 12296
rect 11297 15944 11401 15957
rect 11297 12296 11326 15944
rect 11372 12296 11401 15944
rect 11297 12283 11401 12296
rect 11521 15944 11625 15957
rect 11521 12296 11550 15944
rect 11596 12296 11625 15944
rect 11521 12283 11625 12296
rect 11745 15944 11849 15957
rect 11745 12296 11774 15944
rect 11820 12296 11849 15944
rect 11745 12283 11849 12296
rect 11969 15944 12073 15957
rect 11969 12296 11998 15944
rect 12044 12296 12073 15944
rect 11969 12283 12073 12296
rect 12193 15944 12297 15957
rect 12193 12296 12222 15944
rect 12268 12296 12297 15944
rect 12193 12283 12297 12296
rect 12417 15944 12521 15957
rect 12417 12296 12446 15944
rect 12492 12296 12521 15944
rect 12417 12283 12521 12296
rect 12641 15944 12745 15957
rect 12641 12296 12670 15944
rect 12716 12296 12745 15944
rect 12641 12283 12745 12296
rect 12865 15944 12969 15957
rect 12865 12296 12894 15944
rect 12940 12296 12969 15944
rect 12865 12283 12969 12296
rect 13089 15944 13193 15957
rect 13089 12296 13118 15944
rect 13164 12296 13193 15944
rect 13089 12283 13193 12296
rect 13313 15944 13401 15957
rect 13313 12296 13342 15944
rect 13388 12296 13401 15944
rect 13313 12283 13401 12296
rect 6660 7729 6748 7742
rect 6660 7683 6673 7729
rect 6719 7683 6748 7729
rect 4967 7636 5055 7649
rect 4967 7590 4980 7636
rect 5026 7590 5055 7636
rect 4967 7509 5055 7590
rect 4967 7463 4980 7509
rect 5026 7463 5055 7509
rect 4967 7382 5055 7463
rect 4967 7336 4980 7382
rect 5026 7336 5055 7382
rect 4967 7254 5055 7336
rect 4967 7208 4980 7254
rect 5026 7208 5055 7254
rect 4967 7195 5055 7208
rect 5175 7636 5263 7649
rect 5175 7590 5204 7636
rect 5250 7590 5263 7636
rect 5175 7509 5263 7590
rect 6660 7573 6748 7683
rect 6660 7527 6673 7573
rect 6719 7527 6748 7573
rect 6660 7514 6748 7527
rect 6868 7729 6972 7742
rect 6868 7683 6897 7729
rect 6943 7683 6972 7729
rect 6868 7573 6972 7683
rect 6868 7527 6897 7573
rect 6943 7527 6972 7573
rect 6868 7514 6972 7527
rect 7092 7729 7180 7742
rect 7092 7683 7121 7729
rect 7167 7683 7180 7729
rect 7092 7573 7180 7683
rect 7092 7527 7121 7573
rect 7167 7527 7180 7573
rect 7398 7729 7486 7742
rect 7398 7683 7411 7729
rect 7457 7683 7486 7729
rect 7398 7609 7486 7683
rect 7398 7563 7411 7609
rect 7457 7563 7486 7609
rect 7398 7550 7486 7563
rect 7606 7729 7694 7742
rect 7606 7683 7635 7729
rect 7681 7683 7694 7729
rect 7606 7609 7694 7683
rect 7606 7563 7635 7609
rect 7681 7563 7694 7609
rect 7606 7550 7694 7563
rect 7092 7514 7180 7527
rect 5175 7463 5204 7509
rect 5250 7463 5263 7509
rect 5175 7382 5263 7463
rect 5175 7336 5204 7382
rect 5250 7336 5263 7382
rect 5175 7254 5263 7336
rect 5175 7208 5204 7254
rect 5250 7208 5263 7254
rect 5175 7195 5263 7208
rect 6660 7258 6748 7271
rect 6660 7212 6673 7258
rect 6719 7212 6748 7258
rect 6660 7152 6748 7212
rect 6660 7106 6673 7152
rect 6719 7106 6748 7152
rect 6660 7046 6748 7106
rect 4936 6405 5055 6587
rect 4936 6359 4980 6405
rect 5026 6359 5055 6405
rect 4936 6224 5055 6359
rect 4936 6178 4980 6224
rect 5026 6178 5055 6224
rect 4936 6131 5055 6178
rect 5174 6131 5279 6587
rect 5398 6405 5517 6587
rect 5398 6359 5428 6405
rect 5474 6359 5517 6405
rect 5398 6224 5517 6359
rect 5398 6178 5428 6224
rect 5474 6178 5517 6224
rect 6660 7000 6673 7046
rect 6719 7000 6748 7046
rect 6660 6940 6748 7000
rect 6660 6894 6673 6940
rect 6719 6894 6748 6940
rect 6660 6834 6748 6894
rect 6660 6788 6673 6834
rect 6719 6788 6748 6834
rect 6660 6728 6748 6788
rect 6660 6682 6673 6728
rect 6719 6682 6748 6728
rect 6660 6622 6748 6682
rect 6660 6576 6673 6622
rect 6719 6576 6748 6622
rect 6660 6516 6748 6576
rect 6660 6470 6673 6516
rect 6719 6470 6748 6516
rect 6660 6410 6748 6470
rect 6660 6364 6673 6410
rect 6719 6364 6748 6410
rect 6660 6303 6748 6364
rect 6660 6257 6673 6303
rect 6719 6257 6748 6303
rect 5398 6131 5517 6178
rect 6660 6196 6748 6257
rect 6660 6150 6673 6196
rect 6719 6150 6748 6196
rect 6660 6137 6748 6150
rect 6868 7258 6972 7271
rect 6868 7212 6897 7258
rect 6943 7212 6972 7258
rect 6868 7152 6972 7212
rect 6868 7106 6897 7152
rect 6943 7106 6972 7152
rect 6868 7046 6972 7106
rect 6868 7000 6897 7046
rect 6943 7000 6972 7046
rect 6868 6940 6972 7000
rect 6868 6894 6897 6940
rect 6943 6894 6972 6940
rect 6868 6834 6972 6894
rect 6868 6788 6897 6834
rect 6943 6788 6972 6834
rect 6868 6728 6972 6788
rect 6868 6682 6897 6728
rect 6943 6682 6972 6728
rect 6868 6622 6972 6682
rect 6868 6576 6897 6622
rect 6943 6576 6972 6622
rect 6868 6516 6972 6576
rect 6868 6470 6897 6516
rect 6943 6470 6972 6516
rect 6868 6410 6972 6470
rect 6868 6364 6897 6410
rect 6943 6364 6972 6410
rect 6868 6303 6972 6364
rect 6868 6257 6897 6303
rect 6943 6257 6972 6303
rect 6868 6196 6972 6257
rect 6868 6150 6897 6196
rect 6943 6150 6972 6196
rect 6868 6137 6972 6150
rect 7092 7258 7180 7271
rect 7092 7212 7121 7258
rect 7167 7212 7180 7258
rect 7092 7152 7180 7212
rect 7092 7106 7121 7152
rect 7167 7106 7180 7152
rect 7092 7046 7180 7106
rect 7092 7000 7121 7046
rect 7167 7000 7180 7046
rect 7092 6940 7180 7000
rect 7092 6894 7121 6940
rect 7167 6894 7180 6940
rect 7092 6834 7180 6894
rect 7092 6788 7121 6834
rect 7167 6788 7180 6834
rect 7092 6728 7180 6788
rect 7092 6682 7121 6728
rect 7167 6682 7180 6728
rect 7092 6622 7180 6682
rect 7092 6576 7121 6622
rect 7167 6576 7180 6622
rect 7092 6516 7180 6576
rect 7092 6470 7121 6516
rect 7167 6470 7180 6516
rect 7092 6410 7180 6470
rect 7092 6364 7121 6410
rect 7167 6364 7180 6410
rect 7398 6818 7486 6831
rect 7398 6772 7411 6818
rect 7457 6772 7486 6818
rect 7398 6691 7486 6772
rect 7398 6645 7411 6691
rect 7457 6645 7486 6691
rect 7398 6564 7486 6645
rect 7398 6518 7411 6564
rect 7457 6518 7486 6564
rect 7398 6436 7486 6518
rect 7398 6390 7411 6436
rect 7457 6390 7486 6436
rect 7398 6377 7486 6390
rect 7606 6818 7694 6831
rect 7606 6772 7635 6818
rect 7681 6772 7694 6818
rect 7606 6691 7694 6772
rect 7606 6645 7635 6691
rect 7681 6645 7694 6691
rect 7606 6564 7694 6645
rect 7606 6518 7635 6564
rect 7681 6518 7694 6564
rect 7606 6436 7694 6518
rect 7606 6390 7635 6436
rect 7681 6390 7694 6436
rect 7606 6377 7694 6390
rect 7092 6303 7180 6364
rect 7092 6257 7121 6303
rect 7167 6257 7180 6303
rect 7092 6196 7180 6257
rect 7092 6150 7121 6196
rect 7167 6150 7180 6196
rect 7092 6137 7180 6150
rect 9438 9180 9526 9193
rect 9438 5306 9451 9180
rect 9497 5306 9526 9180
rect 9438 5293 9526 5306
rect 9646 9180 9750 9193
rect 9646 5306 9675 9180
rect 9721 5306 9750 9180
rect 9646 5293 9750 5306
rect 9870 9180 9974 9193
rect 9870 5306 9899 9180
rect 9945 5306 9974 9180
rect 9870 5293 9974 5306
rect 10094 9180 10182 9193
rect 10094 5306 10123 9180
rect 10169 5306 10182 9180
rect 10094 5293 10182 5306
rect 10637 9182 10725 9195
rect 5069 3247 5157 3260
rect 5069 3201 5082 3247
rect 5128 3201 5157 3247
rect 5069 3139 5157 3201
rect 5069 3093 5082 3139
rect 5128 3093 5157 3139
rect 5069 3080 5157 3093
rect 5397 3247 5485 3260
rect 5397 3201 5426 3247
rect 5472 3201 5485 3247
rect 5397 3139 5485 3201
rect 5397 3093 5426 3139
rect 5472 3093 5485 3139
rect 5397 3080 5485 3093
rect 6147 3247 6235 3260
rect 6147 3201 6160 3247
rect 6206 3201 6235 3247
rect 6147 3139 6235 3201
rect 6147 3093 6160 3139
rect 6206 3093 6235 3139
rect 6147 3080 6235 3093
rect 6475 3247 6563 3260
rect 6475 3201 6504 3247
rect 6550 3201 6563 3247
rect 6475 3139 6563 3201
rect 6475 3093 6504 3139
rect 6550 3093 6563 3139
rect 6475 3080 6563 3093
rect 6866 3247 6954 3260
rect 6866 3201 6879 3247
rect 6925 3201 6954 3247
rect 6866 3139 6954 3201
rect 6866 3093 6879 3139
rect 6925 3093 6954 3139
rect 6866 3080 6954 3093
rect 7154 3247 7242 3260
rect 7154 3201 7183 3247
rect 7229 3201 7242 3247
rect 7154 3139 7242 3201
rect 7154 3093 7183 3139
rect 7229 3093 7242 3139
rect 7154 3080 7242 3093
rect 7512 3247 7600 3260
rect 7512 2895 7525 3247
rect 7571 2895 7600 3247
rect 7512 2882 7600 2895
rect 7720 3247 7808 3260
rect 7720 2895 7749 3247
rect 7795 2895 7808 3247
rect 7720 2882 7808 2895
rect 8026 3247 8114 3260
rect 8026 3201 8039 3247
rect 8085 3201 8114 3247
rect 8026 3133 8114 3201
rect 8026 3087 8039 3133
rect 8085 3087 8114 3133
rect 8026 3019 8114 3087
rect 8026 2973 8039 3019
rect 8085 2973 8114 3019
rect 8026 2905 8114 2973
rect 8026 2859 8039 2905
rect 8085 2859 8114 2905
rect 8026 2791 8114 2859
rect 8026 2745 8039 2791
rect 8085 2745 8114 2791
rect 8026 2678 8114 2745
rect 8026 2632 8039 2678
rect 8085 2632 8114 2678
rect 8026 2565 8114 2632
rect 8026 2519 8039 2565
rect 8085 2519 8114 2565
rect 8026 2506 8114 2519
rect 8234 3247 8338 3260
rect 8234 3201 8263 3247
rect 8309 3201 8338 3247
rect 8234 3133 8338 3201
rect 8234 3087 8263 3133
rect 8309 3087 8338 3133
rect 8234 3019 8338 3087
rect 8234 2973 8263 3019
rect 8309 2973 8338 3019
rect 8234 2905 8338 2973
rect 8234 2859 8263 2905
rect 8309 2859 8338 2905
rect 8234 2791 8338 2859
rect 8234 2745 8263 2791
rect 8309 2745 8338 2791
rect 8234 2678 8338 2745
rect 8234 2632 8263 2678
rect 8309 2632 8338 2678
rect 8234 2565 8338 2632
rect 8234 2519 8263 2565
rect 8309 2519 8338 2565
rect 8234 2506 8338 2519
rect 8458 3247 8546 3260
rect 8458 3201 8487 3247
rect 8533 3201 8546 3247
rect 8458 3133 8546 3201
rect 8458 3087 8487 3133
rect 8533 3087 8546 3133
rect 8458 3019 8546 3087
rect 8458 2973 8487 3019
rect 8533 2973 8546 3019
rect 8458 2905 8546 2973
rect 8458 2859 8487 2905
rect 8533 2859 8546 2905
rect 8458 2791 8546 2859
rect 8458 2745 8487 2791
rect 8533 2745 8546 2791
rect 8458 2678 8546 2745
rect 8458 2632 8487 2678
rect 8533 2632 8546 2678
rect 8458 2565 8546 2632
rect 8458 2519 8487 2565
rect 8533 2519 8546 2565
rect 8458 2506 8546 2519
rect 10637 4672 10650 9182
rect 10696 4672 10725 9182
rect 10637 4659 10725 4672
rect 10845 9182 10949 9195
rect 10845 4672 10874 9182
rect 10920 4672 10949 9182
rect 10845 4659 10949 4672
rect 11069 9182 11173 9195
rect 11069 4672 11098 9182
rect 11144 4672 11173 9182
rect 11069 4659 11173 4672
rect 11293 9182 11397 9195
rect 11293 4672 11322 9182
rect 11368 4672 11397 9182
rect 11293 4659 11397 4672
rect 11517 9182 11605 9195
rect 11517 4672 11546 9182
rect 11592 4672 11605 9182
rect 11517 4659 11605 4672
rect 11922 9182 12010 9195
rect 11922 4672 11935 9182
rect 11981 4672 12010 9182
rect 11922 4659 12010 4672
rect 12130 9182 12234 9195
rect 12130 4672 12159 9182
rect 12205 4672 12234 9182
rect 12130 4659 12234 4672
rect 12354 9182 12458 9195
rect 12354 4672 12383 9182
rect 12429 4672 12458 9182
rect 12354 4659 12458 4672
rect 12578 9182 12682 9195
rect 12578 4672 12607 9182
rect 12653 4672 12682 9182
rect 12578 4659 12682 4672
rect 12802 9182 12890 9195
rect 12802 4672 12831 9182
rect 12877 4672 12890 9182
rect 12802 4659 12890 4672
<< mvndiffc >>
rect 6625 9052 6671 11022
rect 6849 9052 6895 11022
rect 7073 9052 7119 11022
rect 7297 9052 7343 11022
rect 7521 9052 7567 11022
rect 7745 9052 7791 11022
rect 8862 9852 8908 11300
rect 9086 9852 9132 11300
rect 9310 9852 9356 11300
rect 9534 9852 9580 11300
rect 9758 9852 9804 11300
rect 9982 9852 10028 11300
rect 10206 9852 10252 11300
rect 10430 9852 10476 11300
rect 10654 9852 10700 11300
rect 10878 9852 10924 11300
rect 11102 9852 11148 11300
rect 11326 9852 11372 11300
rect 11550 9852 11596 11300
rect 11774 9852 11820 11300
rect 11998 9852 12044 11300
rect 12222 9852 12268 11300
rect 12446 9852 12492 11300
rect 12670 9852 12716 11300
rect 12894 9852 12940 11300
rect 13118 9852 13164 11300
rect 13342 9852 13388 11300
rect 6897 8154 6943 8200
rect 4980 8074 5026 8120
rect 4980 7954 5026 8000
rect 5204 8074 5250 8120
rect 6897 8034 6943 8080
rect 7121 8154 7167 8200
rect 7121 8034 7167 8080
rect 7411 8154 7457 8200
rect 7411 8034 7457 8080
rect 7635 8154 7681 8200
rect 7635 8034 7681 8080
rect 5204 7954 5250 8000
rect 6673 5797 6719 5843
rect 4980 5415 5026 5661
rect 5204 5415 5250 5661
rect 5428 5415 5474 5661
rect 6673 5670 6719 5716
rect 6673 5543 6719 5589
rect 6673 5415 6719 5461
rect 6897 5797 6943 5843
rect 6897 5670 6943 5716
rect 6897 5543 6943 5589
rect 6897 5415 6943 5461
rect 7121 5797 7167 5843
rect 7121 5670 7167 5716
rect 7121 5543 7167 5589
rect 7121 5415 7167 5461
rect 7411 5797 7457 5843
rect 7411 5670 7457 5716
rect 7411 5543 7457 5589
rect 7411 5415 7457 5461
rect 7635 5797 7681 5843
rect 7635 5670 7681 5716
rect 7635 5543 7681 5589
rect 7635 5415 7681 5461
rect 8039 4334 8085 4380
rect 8039 4227 8085 4273
rect 8039 4120 8085 4166
rect 8039 4014 8085 4060
rect 5082 3809 5128 3855
rect 5426 3809 5472 3855
rect 6160 3809 6206 3855
rect 6504 3809 6550 3855
rect 6879 3814 6925 3860
rect 7183 3814 7229 3860
rect 7525 3842 7571 3888
rect 7749 3842 7795 3888
rect 8039 3908 8085 3954
rect 8039 3802 8085 3848
rect 8263 4334 8309 4380
rect 8263 4227 8309 4273
rect 8263 4120 8309 4166
rect 8263 4014 8309 4060
rect 8263 3908 8309 3954
rect 8263 3802 8309 3848
rect 9451 4706 9497 4752
rect 9451 4538 9497 4584
rect 9451 4371 9497 4417
rect 9451 4203 9497 4249
rect 9451 4035 9497 4081
rect 9451 3867 9497 3913
rect 9451 3700 9497 3746
rect 9451 3532 9497 3578
rect 9451 3364 9497 3410
rect 9451 3196 9497 3242
rect 9451 3029 9497 3075
rect 9451 2859 9497 2905
rect 9451 2689 9497 2735
rect 9451 2519 9497 2565
rect 9451 2349 9497 2395
rect 9451 2179 9497 2225
rect 9451 2009 9497 2055
rect 9451 1838 9497 1884
rect 9451 1668 9497 1714
rect 9451 1498 9497 1544
rect 9451 1328 9497 1374
rect 9451 1158 9497 1204
rect 9451 988 9497 1034
rect 9451 818 9497 864
rect 9451 648 9497 694
rect 9451 478 9497 524
rect 9451 308 9497 354
rect 10123 4538 10169 4584
rect 10123 4371 10169 4417
rect 10123 4203 10169 4249
rect 10123 4035 10169 4081
rect 10123 3867 10169 3913
rect 10123 3700 10169 3746
rect 10123 3532 10169 3578
rect 10123 3364 10169 3410
rect 10123 3196 10169 3242
rect 10123 3029 10169 3075
rect 10123 2859 10169 2905
rect 10123 2689 10169 2735
rect 10123 2519 10169 2565
rect 10123 2349 10169 2395
rect 10123 2179 10169 2225
rect 10123 2009 10169 2055
rect 10123 1838 10169 1884
rect 10123 1668 10169 1714
rect 10123 1498 10169 1544
rect 10123 1328 10169 1374
rect 10123 1158 10169 1204
rect 10123 988 10169 1034
rect 10123 818 10169 864
rect 10123 648 10169 694
rect 10123 478 10169 524
rect 10650 4022 10696 4068
rect 10650 3854 10696 3900
rect 10650 3686 10696 3732
rect 10650 3518 10696 3564
rect 10650 3351 10696 3397
rect 10650 3183 10696 3229
rect 10650 3015 10696 3061
rect 10650 2847 10696 2893
rect 10650 2680 10696 2726
rect 10650 2512 10696 2558
rect 10650 2344 10696 2390
rect 10650 2174 10696 2220
rect 10650 2004 10696 2050
rect 10650 1834 10696 1880
rect 10650 1664 10696 1710
rect 10650 1494 10696 1540
rect 10650 1324 10696 1370
rect 10650 1154 10696 1200
rect 10650 984 10696 1030
rect 10650 814 10696 860
rect 10650 644 10696 690
rect 11098 4022 11144 4068
rect 11098 3854 11144 3900
rect 11098 3686 11144 3732
rect 11098 3518 11144 3564
rect 11098 3351 11144 3397
rect 11098 3183 11144 3229
rect 11098 3015 11144 3061
rect 11098 2847 11144 2893
rect 11098 2680 11144 2726
rect 11098 2512 11144 2558
rect 11098 2344 11144 2390
rect 11098 2174 11144 2220
rect 11098 2004 11144 2050
rect 11098 1834 11144 1880
rect 11098 1664 11144 1710
rect 11098 1494 11144 1540
rect 11098 1324 11144 1370
rect 11098 1154 11144 1200
rect 11098 984 11144 1030
rect 11098 814 11144 860
rect 11098 644 11144 690
rect 11546 4022 11592 4068
rect 11546 3854 11592 3900
rect 11546 3686 11592 3732
rect 11546 3518 11592 3564
rect 11546 3351 11592 3397
rect 11546 3183 11592 3229
rect 11934 4022 11980 4068
rect 11934 3854 11980 3900
rect 11934 3686 11980 3732
rect 11934 3518 11980 3564
rect 11934 3351 11980 3397
rect 12382 4022 12428 4068
rect 12382 3854 12428 3900
rect 12382 3686 12428 3732
rect 12382 3518 12428 3564
rect 12382 3351 12428 3397
rect 12830 4022 12876 4068
rect 12830 3686 12876 3732
rect 12830 3518 12876 3564
rect 12830 3351 12876 3397
rect 11546 3015 11592 3061
rect 11546 2847 11592 2893
rect 11546 2680 11592 2726
rect 11546 2512 11592 2558
rect 11546 2344 11592 2390
rect 11546 2174 11592 2220
rect 11546 2004 11592 2050
rect 11546 1834 11592 1880
rect 11546 1664 11592 1710
rect 11546 1494 11592 1540
rect 11546 1324 11592 1370
rect 11546 1154 11592 1200
rect 11546 984 11592 1030
rect 11546 814 11592 860
rect 11546 644 11592 690
rect 10123 308 10169 354
<< mvpdiffc >>
rect 6333 13474 6379 15944
rect 6557 13474 6603 15944
rect 6781 13474 6827 15944
rect 7005 13474 7051 15944
rect 7229 13474 7275 15944
rect 7453 13474 7499 15944
rect 7677 13474 7723 15944
rect 7901 13474 7947 15944
rect 8125 13474 8171 15944
rect 8349 13474 8395 15944
rect 8573 13474 8619 15944
rect 8862 12296 8908 15944
rect 9086 12296 9132 15944
rect 9310 12296 9356 15944
rect 9534 12296 9580 15944
rect 9758 12296 9804 15944
rect 9982 12296 10028 15944
rect 10206 12296 10252 15944
rect 10430 12296 10476 15944
rect 10654 12296 10700 15944
rect 10878 12296 10924 15944
rect 11102 12296 11148 15944
rect 11326 12296 11372 15944
rect 11550 12296 11596 15944
rect 11774 12296 11820 15944
rect 11998 12296 12044 15944
rect 12222 12296 12268 15944
rect 12446 12296 12492 15944
rect 12670 12296 12716 15944
rect 12894 12296 12940 15944
rect 13118 12296 13164 15944
rect 13342 12296 13388 15944
rect 6673 7683 6719 7729
rect 4980 7590 5026 7636
rect 4980 7463 5026 7509
rect 4980 7336 5026 7382
rect 4980 7208 5026 7254
rect 5204 7590 5250 7636
rect 6673 7527 6719 7573
rect 6897 7683 6943 7729
rect 6897 7527 6943 7573
rect 7121 7683 7167 7729
rect 7121 7527 7167 7573
rect 7411 7683 7457 7729
rect 7411 7563 7457 7609
rect 7635 7683 7681 7729
rect 7635 7563 7681 7609
rect 5204 7463 5250 7509
rect 5204 7336 5250 7382
rect 5204 7208 5250 7254
rect 6673 7212 6719 7258
rect 6673 7106 6719 7152
rect 4980 6359 5026 6405
rect 4980 6178 5026 6224
rect 5428 6359 5474 6405
rect 5428 6178 5474 6224
rect 6673 7000 6719 7046
rect 6673 6894 6719 6940
rect 6673 6788 6719 6834
rect 6673 6682 6719 6728
rect 6673 6576 6719 6622
rect 6673 6470 6719 6516
rect 6673 6364 6719 6410
rect 6673 6257 6719 6303
rect 6673 6150 6719 6196
rect 6897 7212 6943 7258
rect 6897 7106 6943 7152
rect 6897 7000 6943 7046
rect 6897 6894 6943 6940
rect 6897 6788 6943 6834
rect 6897 6682 6943 6728
rect 6897 6576 6943 6622
rect 6897 6470 6943 6516
rect 6897 6364 6943 6410
rect 6897 6257 6943 6303
rect 6897 6150 6943 6196
rect 7121 7212 7167 7258
rect 7121 7106 7167 7152
rect 7121 7000 7167 7046
rect 7121 6894 7167 6940
rect 7121 6788 7167 6834
rect 7121 6682 7167 6728
rect 7121 6576 7167 6622
rect 7121 6470 7167 6516
rect 7121 6364 7167 6410
rect 7411 6772 7457 6818
rect 7411 6645 7457 6691
rect 7411 6518 7457 6564
rect 7411 6390 7457 6436
rect 7635 6772 7681 6818
rect 7635 6645 7681 6691
rect 7635 6518 7681 6564
rect 7635 6390 7681 6436
rect 7121 6257 7167 6303
rect 7121 6150 7167 6196
rect 9451 5306 9497 9180
rect 9675 5306 9721 9180
rect 9899 5306 9945 9180
rect 10123 5306 10169 9180
rect 5082 3201 5128 3247
rect 5082 3093 5128 3139
rect 5426 3201 5472 3247
rect 5426 3093 5472 3139
rect 6160 3201 6206 3247
rect 6160 3093 6206 3139
rect 6504 3201 6550 3247
rect 6504 3093 6550 3139
rect 6879 3201 6925 3247
rect 6879 3093 6925 3139
rect 7183 3201 7229 3247
rect 7183 3093 7229 3139
rect 7525 2895 7571 3247
rect 7749 2895 7795 3247
rect 8039 3201 8085 3247
rect 8039 3087 8085 3133
rect 8039 2973 8085 3019
rect 8039 2859 8085 2905
rect 8039 2745 8085 2791
rect 8039 2632 8085 2678
rect 8039 2519 8085 2565
rect 8263 3201 8309 3247
rect 8263 3087 8309 3133
rect 8263 2973 8309 3019
rect 8263 2859 8309 2905
rect 8263 2745 8309 2791
rect 8263 2632 8309 2678
rect 8263 2519 8309 2565
rect 8487 3201 8533 3247
rect 8487 3087 8533 3133
rect 8487 2973 8533 3019
rect 8487 2859 8533 2905
rect 8487 2745 8533 2791
rect 8487 2632 8533 2678
rect 8487 2519 8533 2565
rect 10650 4672 10696 9182
rect 10874 4672 10920 9182
rect 11098 4672 11144 9182
rect 11322 4672 11368 9182
rect 11546 4672 11592 9182
rect 11935 4672 11981 9182
rect 12159 4672 12205 9182
rect 12383 4672 12429 9182
rect 12607 4672 12653 9182
rect 12831 4672 12877 9182
<< mvpsubdiff >>
rect 7991 11596 13744 11653
rect 7991 11550 13643 11596
rect 13689 11550 13744 11596
rect 7991 11543 13744 11550
rect 7991 11536 8304 11543
rect 7990 11535 8304 11536
rect 6269 11478 8304 11535
rect 6269 11432 6323 11478
rect 6369 11432 6481 11478
rect 6527 11432 6639 11478
rect 6685 11432 6798 11478
rect 6844 11432 6956 11478
rect 7002 11432 7114 11478
rect 7160 11432 7272 11478
rect 7318 11432 7430 11478
rect 7476 11432 7588 11478
rect 7634 11432 7747 11478
rect 7793 11432 7905 11478
rect 7951 11432 8063 11478
rect 8109 11432 8304 11478
rect 6269 11375 8304 11432
rect 6269 11315 6424 11375
rect 6269 11269 6323 11315
rect 6369 11269 6424 11315
rect 6269 11152 6424 11269
rect 7991 11243 8304 11375
rect 13588 11433 13744 11543
rect 13588 11387 13643 11433
rect 13689 11387 13744 11433
rect 7991 11197 8045 11243
rect 8091 11197 8203 11243
rect 8249 11197 8304 11243
rect 6269 11106 6323 11152
rect 6369 11106 6424 11152
rect 6269 10988 6424 11106
rect 7991 11080 8304 11197
rect 6269 10942 6323 10988
rect 6369 10942 6424 10988
rect 6269 10825 6424 10942
rect 6269 10779 6323 10825
rect 6369 10779 6424 10825
rect 6269 10662 6424 10779
rect 6269 10616 6323 10662
rect 6369 10616 6424 10662
rect 6269 10499 6424 10616
rect 6269 10453 6323 10499
rect 6369 10453 6424 10499
rect 6269 10335 6424 10453
rect 6269 10289 6323 10335
rect 6369 10289 6424 10335
rect 6269 10172 6424 10289
rect 6269 10126 6323 10172
rect 6369 10126 6424 10172
rect 6269 10009 6424 10126
rect 6269 9963 6323 10009
rect 6369 9963 6424 10009
rect 6269 9845 6424 9963
rect 6269 9799 6323 9845
rect 6369 9799 6424 9845
rect 6269 9682 6424 9799
rect 6269 9636 6323 9682
rect 6369 9636 6424 9682
rect 6269 9519 6424 9636
rect 6269 9473 6323 9519
rect 6369 9473 6424 9519
rect 6269 9356 6424 9473
rect 6269 9310 6323 9356
rect 6369 9310 6424 9356
rect 6269 9192 6424 9310
rect 6269 9146 6323 9192
rect 6369 9146 6424 9192
rect 6269 9029 6424 9146
rect 7991 11034 8045 11080
rect 8091 11034 8203 11080
rect 8249 11034 8304 11080
rect 7991 10917 8304 11034
rect 7991 10871 8045 10917
rect 8091 10871 8203 10917
rect 8249 10871 8304 10917
rect 7991 10753 8304 10871
rect 7991 10707 8045 10753
rect 8091 10707 8203 10753
rect 8249 10707 8304 10753
rect 7991 10590 8304 10707
rect 7991 10544 8045 10590
rect 8091 10544 8203 10590
rect 8249 10544 8304 10590
rect 7991 10427 8304 10544
rect 7991 10381 8045 10427
rect 8091 10381 8203 10427
rect 8249 10381 8304 10427
rect 7991 10264 8304 10381
rect 7991 10218 8045 10264
rect 8091 10218 8203 10264
rect 8249 10218 8304 10264
rect 7991 10100 8304 10218
rect 7991 10054 8045 10100
rect 8091 10054 8203 10100
rect 8249 10054 8304 10100
rect 7991 9937 8304 10054
rect 7991 9891 8045 9937
rect 8091 9891 8203 9937
rect 8249 9891 8304 9937
rect 7991 9774 8304 9891
rect 13588 11270 13744 11387
rect 13588 11224 13643 11270
rect 13689 11224 13744 11270
rect 13588 11107 13744 11224
rect 13588 11061 13643 11107
rect 13689 11061 13744 11107
rect 13588 10943 13744 11061
rect 13588 10897 13643 10943
rect 13689 10897 13744 10943
rect 13588 10780 13744 10897
rect 13588 10734 13643 10780
rect 13689 10734 13744 10780
rect 13588 10617 13744 10734
rect 13588 10571 13643 10617
rect 13689 10571 13744 10617
rect 13588 10453 13744 10571
rect 13588 10407 13643 10453
rect 13689 10407 13744 10453
rect 13588 10290 13744 10407
rect 13588 10244 13643 10290
rect 13689 10244 13744 10290
rect 13588 10127 13744 10244
rect 13588 10081 13643 10127
rect 13689 10081 13744 10127
rect 13588 9964 13744 10081
rect 13588 9918 13643 9964
rect 13689 9918 13744 9964
rect 13588 9861 13744 9918
rect 7991 9728 8045 9774
rect 8091 9728 8203 9774
rect 8249 9728 8304 9774
rect 7991 9610 8304 9728
rect 7991 9564 8045 9610
rect 8091 9564 8203 9610
rect 8249 9564 8304 9610
rect 7991 9447 8304 9564
rect 7991 9401 8045 9447
rect 8091 9401 8203 9447
rect 8249 9401 8304 9447
rect 7991 9284 8304 9401
rect 7991 9238 8045 9284
rect 8091 9238 8203 9284
rect 8249 9238 8304 9284
rect 7991 9121 8304 9238
rect 7991 9075 8045 9121
rect 8091 9075 8203 9121
rect 8249 9075 8304 9121
rect 6269 8983 6323 9029
rect 6369 8983 6424 9029
rect 6269 8866 6424 8983
rect 6269 8820 6323 8866
rect 6369 8820 6424 8866
rect 6269 8688 6424 8820
rect 7991 8957 8304 9075
rect 7991 8911 8045 8957
rect 8091 8911 8203 8957
rect 8249 8911 8304 8957
rect 7991 8794 8304 8911
rect 7991 8748 8045 8794
rect 8091 8748 8203 8794
rect 8249 8748 8304 8794
rect 7991 8688 8304 8748
rect 346 8631 8304 8688
rect 346 8585 400 8631
rect 446 8585 558 8631
rect 604 8585 716 8631
rect 762 8585 875 8631
rect 921 8585 1033 8631
rect 1079 8585 1191 8631
rect 1237 8585 1349 8631
rect 1395 8585 1507 8631
rect 1553 8585 1665 8631
rect 1711 8585 1823 8631
rect 1869 8585 1981 8631
rect 2027 8585 2139 8631
rect 2185 8585 2298 8631
rect 2344 8585 2456 8631
rect 2502 8585 2614 8631
rect 2660 8585 2772 8631
rect 2818 8585 2930 8631
rect 2976 8585 3088 8631
rect 3134 8585 3246 8631
rect 3292 8585 3404 8631
rect 3450 8585 3562 8631
rect 3608 8585 3721 8631
rect 3767 8585 3879 8631
rect 3925 8585 4037 8631
rect 4083 8585 4195 8631
rect 4241 8585 4353 8631
rect 4399 8585 4511 8631
rect 4557 8585 4670 8631
rect 4716 8585 4828 8631
rect 4874 8585 4986 8631
rect 5032 8585 5144 8631
rect 5190 8585 5302 8631
rect 5348 8585 5460 8631
rect 5506 8585 5618 8631
rect 5664 8585 5776 8631
rect 5822 8585 5934 8631
rect 5980 8585 6093 8631
rect 6139 8585 6251 8631
rect 6297 8585 6409 8631
rect 6455 8585 6567 8631
rect 6613 8585 6725 8631
rect 6771 8585 6883 8631
rect 6929 8585 7041 8631
rect 7087 8585 7199 8631
rect 7245 8585 7357 8631
rect 7403 8585 7516 8631
rect 7562 8585 7674 8631
rect 7720 8585 7832 8631
rect 7878 8585 8045 8631
rect 8091 8585 8203 8631
rect 8249 8585 8304 8631
rect 346 8528 8304 8585
rect 346 8306 4301 8528
rect 6269 8523 6424 8528
rect 346 8260 403 8306
rect 449 8260 561 8306
rect 607 8260 719 8306
rect 765 8260 877 8306
rect 923 8260 1035 8306
rect 1081 8260 1193 8306
rect 1239 8260 1351 8306
rect 1397 8260 1509 8306
rect 1555 8260 1667 8306
rect 1713 8260 1826 8306
rect 1872 8260 1984 8306
rect 2030 8260 2142 8306
rect 2188 8260 2300 8306
rect 2346 8260 2458 8306
rect 2504 8260 2616 8306
rect 2662 8260 2774 8306
rect 2820 8260 2933 8306
rect 2979 8260 3091 8306
rect 3137 8260 3249 8306
rect 3295 8260 3407 8306
rect 3453 8260 3565 8306
rect 3611 8260 3723 8306
rect 3769 8260 3881 8306
rect 3927 8260 4039 8306
rect 4085 8260 4197 8306
rect 4243 8260 4301 8306
rect 346 8143 4301 8260
rect 346 8097 403 8143
rect 449 8097 561 8143
rect 607 8097 719 8143
rect 765 8097 877 8143
rect 923 8097 1035 8143
rect 1081 8097 1193 8143
rect 1239 8097 1351 8143
rect 1397 8097 1509 8143
rect 1555 8097 1667 8143
rect 1713 8097 1826 8143
rect 1872 8097 1984 8143
rect 2030 8097 2142 8143
rect 2188 8097 2300 8143
rect 2346 8097 2458 8143
rect 2504 8097 2616 8143
rect 2662 8097 2774 8143
rect 2820 8097 2933 8143
rect 2979 8097 3091 8143
rect 3137 8097 3249 8143
rect 3295 8097 3407 8143
rect 3453 8097 3565 8143
rect 3611 8097 3723 8143
rect 3769 8097 3881 8143
rect 3927 8097 4039 8143
rect 4085 8097 4197 8143
rect 4243 8097 4301 8143
rect 346 7980 4301 8097
rect 346 7934 403 7980
rect 449 7934 561 7980
rect 607 7934 719 7980
rect 765 7934 877 7980
rect 923 7934 1035 7980
rect 1081 7934 1193 7980
rect 1239 7934 1351 7980
rect 1397 7934 1509 7980
rect 1555 7934 1667 7980
rect 1713 7934 1826 7980
rect 1872 7934 1984 7980
rect 2030 7934 2142 7980
rect 2188 7934 2300 7980
rect 2346 7934 2458 7980
rect 2504 7934 2616 7980
rect 2662 7934 2774 7980
rect 2820 7934 2933 7980
rect 2979 7934 3091 7980
rect 3137 7934 3249 7980
rect 3295 7934 3407 7980
rect 3453 7934 3565 7980
rect 3611 7934 3723 7980
rect 3769 7934 3881 7980
rect 3927 7934 4039 7980
rect 4085 7934 4197 7980
rect 4243 7934 4301 7980
rect 346 7875 4301 7934
rect 685 5931 4476 5988
rect 685 5885 739 5931
rect 785 5885 897 5931
rect 943 5885 1055 5931
rect 1101 5885 1213 5931
rect 1259 5885 1371 5931
rect 1417 5885 1529 5931
rect 1575 5885 1687 5931
rect 1733 5885 1845 5931
rect 1891 5885 2003 5931
rect 2049 5885 2162 5931
rect 2208 5885 2320 5931
rect 2366 5885 2478 5931
rect 2524 5885 2636 5931
rect 2682 5885 2794 5931
rect 2840 5885 2952 5931
rect 2998 5885 3111 5931
rect 3157 5885 3269 5931
rect 3315 5885 3427 5931
rect 3473 5885 3585 5931
rect 3631 5885 3743 5931
rect 3789 5885 3901 5931
rect 3947 5885 4059 5931
rect 4105 5885 4217 5931
rect 4263 5885 4375 5931
rect 4421 5885 4476 5931
rect 685 5768 4476 5885
rect 685 5722 739 5768
rect 785 5722 897 5768
rect 943 5722 1055 5768
rect 1101 5722 1213 5768
rect 1259 5722 1371 5768
rect 1417 5722 1529 5768
rect 1575 5722 1687 5768
rect 1733 5722 1845 5768
rect 1891 5722 2003 5768
rect 2049 5722 2162 5768
rect 2208 5722 2320 5768
rect 2366 5722 2478 5768
rect 2524 5722 2636 5768
rect 2682 5722 2794 5768
rect 2840 5722 2952 5768
rect 2998 5722 3111 5768
rect 3157 5722 3269 5768
rect 3315 5722 3427 5768
rect 3473 5722 3585 5768
rect 3631 5722 3743 5768
rect 3789 5722 3901 5768
rect 3947 5722 4059 5768
rect 4105 5722 4217 5768
rect 4263 5722 4375 5768
rect 4421 5722 4476 5768
rect 685 5605 4476 5722
rect 6339 5707 6473 5766
rect 685 5559 739 5605
rect 785 5559 897 5605
rect 943 5559 1055 5605
rect 1101 5559 1213 5605
rect 1259 5559 1371 5605
rect 1417 5559 1529 5605
rect 1575 5559 1687 5605
rect 1733 5559 1845 5605
rect 1891 5559 2003 5605
rect 2049 5559 2162 5605
rect 2208 5559 2320 5605
rect 2366 5559 2478 5605
rect 2524 5559 2636 5605
rect 2682 5559 2794 5605
rect 2840 5559 2952 5605
rect 2998 5559 3111 5605
rect 3157 5559 3269 5605
rect 3315 5559 3427 5605
rect 3473 5559 3585 5605
rect 3631 5559 3743 5605
rect 3789 5559 3901 5605
rect 3947 5559 4059 5605
rect 4105 5559 4217 5605
rect 4263 5559 4375 5605
rect 4421 5559 4476 5605
rect 685 5501 4476 5559
rect 6339 5661 6383 5707
rect 6429 5661 6473 5707
rect 6339 5543 6473 5661
rect 6339 5497 6383 5543
rect 6429 5497 6473 5543
rect 6339 5016 6473 5497
rect 295 4997 7779 5016
rect 295 4351 314 4997
rect 7760 4351 7779 4997
rect 8869 4720 9187 4779
rect 8869 4674 8926 4720
rect 8972 4674 9084 4720
rect 9130 4674 9187 4720
rect 8869 4557 9187 4674
rect 8869 4511 8926 4557
rect 8972 4511 9084 4557
rect 9130 4511 9187 4557
rect 8869 4394 9187 4511
rect 295 4332 7779 4351
rect 8869 4348 8926 4394
rect 8972 4348 9084 4394
rect 9130 4348 9187 4394
rect 8869 4230 9187 4348
rect 8869 4184 8926 4230
rect 8972 4184 9084 4230
rect 9130 4184 9187 4230
rect 8869 4067 9187 4184
rect 8869 4021 8926 4067
rect 8972 4021 9084 4067
rect 9130 4021 9187 4067
rect 8869 3904 9187 4021
rect 8869 3858 8926 3904
rect 8972 3858 9084 3904
rect 9130 3858 9187 3904
rect 8869 3741 9187 3858
rect 8869 3695 8926 3741
rect 8972 3695 9084 3741
rect 9130 3695 9187 3741
rect 8869 3577 9187 3695
rect 8869 3531 8926 3577
rect 8972 3531 9084 3577
rect 9130 3531 9187 3577
rect 8869 3414 9187 3531
rect 8869 3368 8926 3414
rect 8972 3368 9084 3414
rect 9130 3368 9187 3414
rect 8869 3251 9187 3368
rect 8869 3205 8926 3251
rect 8972 3205 9084 3251
rect 9130 3205 9187 3251
rect 8869 3088 9187 3205
rect 8869 3042 8926 3088
rect 8972 3042 9084 3088
rect 9130 3042 9187 3088
rect 8869 2925 9187 3042
rect 8869 2879 8926 2925
rect 8972 2879 9084 2925
rect 9130 2879 9187 2925
rect 8869 2761 9187 2879
rect 8869 2715 8926 2761
rect 8972 2715 9084 2761
rect 9130 2715 9187 2761
rect 8869 2598 9187 2715
rect 8869 2552 8926 2598
rect 8972 2552 9084 2598
rect 9130 2552 9187 2598
rect 8869 2435 9187 2552
rect 8869 2389 8926 2435
rect 8972 2389 9084 2435
rect 9130 2389 9187 2435
rect 8869 2271 9187 2389
rect 8869 2225 8926 2271
rect 8972 2225 9084 2271
rect 9130 2225 9187 2271
rect 8869 2108 9187 2225
rect 8869 2062 8926 2108
rect 8972 2062 9084 2108
rect 9130 2062 9187 2108
rect 8869 1945 9187 2062
rect 8869 1899 8926 1945
rect 8972 1899 9084 1945
rect 9130 1899 9187 1945
rect 8869 1781 9187 1899
rect 8869 1735 8926 1781
rect 8972 1735 9084 1781
rect 9130 1735 9187 1781
rect 8869 1618 9187 1735
rect 8869 1572 8926 1618
rect 8972 1572 9084 1618
rect 9130 1572 9187 1618
rect 8869 1455 9187 1572
rect 8869 1409 8926 1455
rect 8972 1409 9084 1455
rect 9130 1409 9187 1455
rect 8869 1292 9187 1409
rect 8869 1246 8926 1292
rect 8972 1246 9084 1292
rect 9130 1246 9187 1292
rect 8869 1129 9187 1246
rect 8869 1083 8926 1129
rect 8972 1083 9084 1129
rect 9130 1083 9187 1129
rect 8869 965 9187 1083
rect 8869 919 8926 965
rect 8972 919 9084 965
rect 9130 919 9187 965
rect 8869 802 9187 919
rect 8869 756 8926 802
rect 8972 756 9084 802
rect 9130 756 9187 802
rect 8869 639 9187 756
rect 8869 593 8926 639
rect 8972 593 9084 639
rect 9130 593 9187 639
rect 8869 476 9187 593
rect 8869 430 8926 476
rect 8972 430 9084 476
rect 9130 430 9187 476
rect 8869 312 9187 430
rect 8869 266 8926 312
rect 8972 266 9084 312
rect 9130 266 9187 312
rect 8869 149 9187 266
rect 13296 4237 13614 4290
rect 13296 4191 13353 4237
rect 13399 4191 13511 4237
rect 13557 4191 13614 4237
rect 13296 4074 13614 4191
rect 13296 4028 13353 4074
rect 13399 4028 13511 4074
rect 13557 4028 13614 4074
rect 13296 3905 13614 4028
rect 13296 3859 13353 3905
rect 13399 3859 13511 3905
rect 13557 3859 13614 3905
rect 13296 3742 13614 3859
rect 13296 3696 13353 3742
rect 13399 3696 13511 3742
rect 13557 3696 13614 3742
rect 13296 3578 13614 3696
rect 13296 3532 13353 3578
rect 13399 3532 13511 3578
rect 13557 3532 13614 3578
rect 13296 3415 13614 3532
rect 13296 3369 13353 3415
rect 13399 3369 13511 3415
rect 13557 3369 13614 3415
rect 13296 3252 13614 3369
rect 13296 3206 13353 3252
rect 13399 3206 13511 3252
rect 13557 3206 13614 3252
rect 13296 3089 13614 3206
rect 13296 3043 13353 3089
rect 13399 3043 13511 3089
rect 13557 3043 13614 3089
rect 13296 2925 13614 3043
rect 13296 2879 13353 2925
rect 13399 2879 13511 2925
rect 13557 2879 13614 2925
rect 13296 2762 13614 2879
rect 13296 2716 13353 2762
rect 13399 2716 13511 2762
rect 13557 2716 13614 2762
rect 13296 2599 13614 2716
rect 13296 2553 13353 2599
rect 13399 2553 13511 2599
rect 13557 2553 13614 2599
rect 13296 2436 13614 2553
rect 13296 2390 13353 2436
rect 13399 2390 13511 2436
rect 13557 2390 13614 2436
rect 13296 2272 13614 2390
rect 13296 2226 13353 2272
rect 13399 2226 13511 2272
rect 13557 2226 13614 2272
rect 13296 2109 13614 2226
rect 13296 2063 13353 2109
rect 13399 2063 13511 2109
rect 13557 2063 13614 2109
rect 13296 1946 13614 2063
rect 13296 1900 13353 1946
rect 13399 1900 13511 1946
rect 13557 1900 13614 1946
rect 13296 1782 13614 1900
rect 13296 1736 13353 1782
rect 13399 1736 13511 1782
rect 13557 1736 13614 1782
rect 13296 1619 13614 1736
rect 13296 1573 13353 1619
rect 13399 1573 13511 1619
rect 13557 1573 13614 1619
rect 13296 1456 13614 1573
rect 13296 1410 13353 1456
rect 13399 1410 13511 1456
rect 13557 1410 13614 1456
rect 13296 1293 13614 1410
rect 13296 1247 13353 1293
rect 13399 1247 13511 1293
rect 13557 1247 13614 1293
rect 13296 1129 13614 1247
rect 13296 1083 13353 1129
rect 13399 1083 13511 1129
rect 13557 1083 13614 1129
rect 13296 966 13614 1083
rect 13296 920 13353 966
rect 13399 920 13511 966
rect 13557 920 13614 966
rect 13296 803 13614 920
rect 13296 757 13353 803
rect 13399 757 13511 803
rect 13557 757 13614 803
rect 13296 640 13614 757
rect 13296 594 13353 640
rect 13399 594 13511 640
rect 13557 594 13614 640
rect 13296 476 13614 594
rect 13296 430 13353 476
rect 13399 430 13511 476
rect 13557 430 13614 476
rect 13296 313 13614 430
rect 13296 267 13353 313
rect 13399 267 13511 313
rect 13557 267 13614 313
rect 8869 103 8926 149
rect 8972 103 9084 149
rect 9130 103 9187 149
rect 8869 46 9187 103
rect 13296 150 13614 267
rect 13296 104 13353 150
rect 13399 104 13511 150
rect 13557 104 13614 150
rect 13296 46 13614 104
rect 8869 45 9188 46
rect 13296 45 13615 46
rect 8869 -13 13615 45
rect 8869 -14 13353 -13
rect 8869 -60 8926 -14
rect 8972 -60 9084 -14
rect 9130 -60 9401 -14
rect 9447 -60 9559 -14
rect 9605 -60 9717 -14
rect 9763 -60 9875 -14
rect 9921 -60 10033 -14
rect 10079 -60 10191 -14
rect 10237 -60 10349 -14
rect 10395 -60 10507 -14
rect 10553 -60 10665 -14
rect 10711 -60 10824 -14
rect 10870 -60 10982 -14
rect 11028 -60 11140 -14
rect 11186 -60 11298 -14
rect 11344 -60 11456 -14
rect 11502 -60 11614 -14
rect 11660 -60 11772 -14
rect 11818 -60 11931 -14
rect 11977 -60 12089 -14
rect 12135 -60 12247 -14
rect 12293 -60 12405 -14
rect 12451 -60 12563 -14
rect 12609 -60 12721 -14
rect 12767 -60 12879 -14
rect 12925 -60 13037 -14
rect 13083 -60 13195 -14
rect 13241 -59 13353 -14
rect 13399 -59 13511 -13
rect 13557 -59 13615 -13
rect 13241 -60 13615 -59
rect 8869 -119 13615 -60
rect 9027 -120 13615 -119
<< mvnsubdiff >>
rect 5994 16273 13722 16319
rect 5994 16227 6192 16273
rect 6238 16227 6350 16273
rect 6396 16227 6508 16273
rect 6554 16227 6666 16273
rect 6712 16227 6824 16273
rect 6870 16227 6982 16273
rect 7028 16227 7140 16273
rect 7186 16227 7298 16273
rect 7344 16227 7457 16273
rect 7503 16227 7615 16273
rect 7661 16227 7773 16273
rect 7819 16227 7931 16273
rect 7977 16227 8089 16273
rect 8135 16227 8247 16273
rect 8293 16227 8405 16273
rect 8451 16227 8563 16273
rect 8609 16227 8721 16273
rect 8767 16227 8880 16273
rect 8926 16227 9038 16273
rect 9084 16227 9196 16273
rect 9242 16227 9354 16273
rect 9400 16227 9512 16273
rect 9558 16227 9670 16273
rect 9716 16227 9828 16273
rect 9874 16227 9986 16273
rect 10032 16227 10144 16273
rect 10190 16227 10303 16273
rect 10349 16227 10461 16273
rect 10507 16227 10619 16273
rect 10665 16227 10777 16273
rect 10823 16227 10935 16273
rect 10981 16227 11093 16273
rect 11139 16227 11251 16273
rect 11297 16227 11409 16273
rect 11455 16227 11567 16273
rect 11613 16227 11726 16273
rect 11772 16227 11884 16273
rect 11930 16227 12042 16273
rect 12088 16227 12200 16273
rect 12246 16227 12358 16273
rect 12404 16227 12516 16273
rect 12562 16227 12674 16273
rect 12720 16227 12832 16273
rect 12878 16227 12990 16273
rect 13036 16227 13149 16273
rect 13195 16227 13307 16273
rect 13353 16227 13465 16273
rect 13511 16227 13722 16273
rect 5994 16181 13722 16227
rect 5994 16092 6128 16181
rect 5994 16046 6038 16092
rect 6084 16046 6128 16092
rect 5994 15928 6128 16046
rect 13588 16092 13722 16181
rect 13588 16046 13632 16092
rect 13678 16046 13722 16092
rect 5994 15882 6038 15928
rect 6084 15882 6128 15928
rect 5994 15765 6128 15882
rect 5994 15719 6038 15765
rect 6084 15719 6128 15765
rect 5994 15602 6128 15719
rect 5994 15556 6038 15602
rect 6084 15556 6128 15602
rect 5994 15439 6128 15556
rect 5994 15393 6038 15439
rect 6084 15393 6128 15439
rect 5994 15275 6128 15393
rect 5994 15229 6038 15275
rect 6084 15229 6128 15275
rect 5994 15112 6128 15229
rect 5994 15066 6038 15112
rect 6084 15066 6128 15112
rect 5994 14949 6128 15066
rect 5994 14903 6038 14949
rect 6084 14903 6128 14949
rect 5994 14786 6128 14903
rect 5994 14740 6038 14786
rect 6084 14740 6128 14786
rect 5994 14622 6128 14740
rect 5994 14576 6038 14622
rect 6084 14576 6128 14622
rect 5994 14459 6128 14576
rect 5994 14413 6038 14459
rect 6084 14413 6128 14459
rect 5994 14296 6128 14413
rect 5994 14250 6038 14296
rect 6084 14250 6128 14296
rect 5994 14133 6128 14250
rect 5994 14087 6038 14133
rect 6084 14087 6128 14133
rect 5994 13970 6128 14087
rect 5994 13924 6038 13970
rect 6084 13924 6128 13970
rect 5994 13806 6128 13924
rect 5994 13760 6038 13806
rect 6084 13760 6128 13806
rect 5994 13643 6128 13760
rect 5994 13597 6038 13643
rect 6084 13597 6128 13643
rect 5994 13480 6128 13597
rect 5994 13434 6038 13480
rect 6084 13434 6128 13480
rect 5994 13317 6128 13434
rect 5994 13271 6038 13317
rect 6084 13271 6128 13317
rect 5994 13161 6128 13271
rect 5994 13153 8664 13161
rect 5994 13107 6038 13153
rect 6084 13107 8664 13153
rect 5994 13104 8664 13107
rect 5994 13058 6349 13104
rect 6395 13058 6507 13104
rect 6553 13058 6665 13104
rect 6711 13058 6823 13104
rect 6869 13058 6982 13104
rect 7028 13058 7140 13104
rect 7186 13058 7298 13104
rect 7344 13058 7456 13104
rect 7502 13058 7614 13104
rect 7660 13058 7772 13104
rect 7818 13058 7930 13104
rect 7976 13058 8089 13104
rect 8135 13058 8247 13104
rect 8293 13058 8405 13104
rect 8451 13058 8563 13104
rect 8609 13058 8664 13104
rect 5994 12990 8664 13058
rect 5994 12944 6038 12990
rect 6084 12944 8664 12990
rect 5994 12941 8664 12944
rect 5994 12895 6349 12941
rect 6395 12895 6507 12941
rect 6553 12895 6665 12941
rect 6711 12895 6823 12941
rect 6869 12895 6982 12941
rect 7028 12895 7140 12941
rect 7186 12895 7298 12941
rect 7344 12895 7456 12941
rect 7502 12895 7614 12941
rect 7660 12895 7772 12941
rect 7818 12895 7930 12941
rect 7976 12895 8089 12941
rect 8135 12895 8247 12941
rect 8293 12895 8405 12941
rect 8451 12895 8563 12941
rect 8609 12895 8664 12941
rect 5994 12827 8664 12895
rect 5994 12781 6038 12827
rect 6084 12781 8664 12827
rect 5994 12777 8664 12781
rect 5994 12731 6349 12777
rect 6395 12731 6507 12777
rect 6553 12731 6665 12777
rect 6711 12731 6823 12777
rect 6869 12731 6982 12777
rect 7028 12731 7140 12777
rect 7186 12731 7298 12777
rect 7344 12731 7456 12777
rect 7502 12731 7614 12777
rect 7660 12731 7772 12777
rect 7818 12731 7930 12777
rect 7976 12731 8089 12777
rect 8135 12731 8247 12777
rect 8293 12731 8405 12777
rect 8451 12731 8563 12777
rect 8609 12731 8664 12777
rect 5994 12664 8664 12731
rect 5994 12618 6038 12664
rect 6084 12618 8664 12664
rect 5994 12614 8664 12618
rect 5994 12568 6349 12614
rect 6395 12568 6507 12614
rect 6553 12568 6665 12614
rect 6711 12568 6823 12614
rect 6869 12568 6982 12614
rect 7028 12568 7140 12614
rect 7186 12568 7298 12614
rect 7344 12568 7456 12614
rect 7502 12568 7614 12614
rect 7660 12568 7772 12614
rect 7818 12568 7930 12614
rect 7976 12568 8089 12614
rect 8135 12568 8247 12614
rect 8293 12568 8405 12614
rect 8451 12568 8563 12614
rect 8609 12568 8664 12614
rect 5994 12501 8664 12568
rect 5994 12455 6038 12501
rect 6084 12455 8664 12501
rect 5994 12451 8664 12455
rect 5994 12405 6349 12451
rect 6395 12405 6507 12451
rect 6553 12405 6665 12451
rect 6711 12405 6823 12451
rect 6869 12405 6982 12451
rect 7028 12405 7140 12451
rect 7186 12405 7298 12451
rect 7344 12405 7456 12451
rect 7502 12405 7614 12451
rect 7660 12405 7772 12451
rect 7818 12405 7930 12451
rect 7976 12405 8089 12451
rect 8135 12405 8247 12451
rect 8293 12405 8405 12451
rect 8451 12405 8563 12451
rect 8609 12405 8664 12451
rect 5994 12337 8664 12405
rect 5994 12291 6038 12337
rect 6084 12291 8664 12337
rect 5994 12287 8664 12291
rect 5994 12241 6349 12287
rect 6395 12241 6507 12287
rect 6553 12241 6665 12287
rect 6711 12241 6823 12287
rect 6869 12241 6982 12287
rect 7028 12241 7140 12287
rect 7186 12241 7298 12287
rect 7344 12241 7456 12287
rect 7502 12241 7614 12287
rect 7660 12241 7772 12287
rect 7818 12241 7930 12287
rect 7976 12241 8089 12287
rect 8135 12241 8247 12287
rect 8293 12241 8405 12287
rect 8451 12241 8563 12287
rect 8609 12241 8664 12287
rect 13588 15928 13722 16046
rect 13588 15882 13632 15928
rect 13678 15882 13722 15928
rect 13588 15765 13722 15882
rect 13588 15719 13632 15765
rect 13678 15719 13722 15765
rect 13588 15602 13722 15719
rect 13588 15556 13632 15602
rect 13678 15556 13722 15602
rect 13588 15439 13722 15556
rect 13588 15393 13632 15439
rect 13678 15393 13722 15439
rect 13588 15275 13722 15393
rect 13588 15229 13632 15275
rect 13678 15229 13722 15275
rect 13588 15112 13722 15229
rect 13588 15066 13632 15112
rect 13678 15066 13722 15112
rect 13588 14949 13722 15066
rect 13588 14903 13632 14949
rect 13678 14903 13722 14949
rect 13588 14786 13722 14903
rect 13588 14740 13632 14786
rect 13678 14740 13722 14786
rect 13588 14622 13722 14740
rect 13588 14576 13632 14622
rect 13678 14576 13722 14622
rect 13588 14459 13722 14576
rect 13588 14413 13632 14459
rect 13678 14413 13722 14459
rect 13588 14296 13722 14413
rect 13588 14250 13632 14296
rect 13678 14250 13722 14296
rect 13588 14133 13722 14250
rect 13588 14087 13632 14133
rect 13678 14087 13722 14133
rect 13588 13970 13722 14087
rect 13588 13924 13632 13970
rect 13678 13924 13722 13970
rect 13588 13806 13722 13924
rect 13588 13760 13632 13806
rect 13678 13760 13722 13806
rect 13588 13643 13722 13760
rect 13588 13597 13632 13643
rect 13678 13597 13722 13643
rect 13588 13480 13722 13597
rect 13588 13434 13632 13480
rect 13678 13434 13722 13480
rect 13588 13317 13722 13434
rect 13588 13271 13632 13317
rect 13678 13271 13722 13317
rect 13588 13153 13722 13271
rect 13588 13107 13632 13153
rect 13678 13107 13722 13153
rect 13588 12990 13722 13107
rect 13588 12944 13632 12990
rect 13678 12944 13722 12990
rect 13588 12827 13722 12944
rect 13588 12781 13632 12827
rect 13678 12781 13722 12827
rect 13588 12664 13722 12781
rect 13588 12618 13632 12664
rect 13678 12618 13722 12664
rect 13588 12501 13722 12618
rect 13588 12455 13632 12501
rect 13678 12455 13722 12501
rect 13588 12337 13722 12455
rect 13588 12291 13632 12337
rect 13678 12291 13722 12337
rect 5994 12174 8664 12241
rect 5994 12128 6038 12174
rect 6084 12128 8664 12174
rect 13588 12174 13722 12291
rect 5994 12124 8664 12128
rect 5994 12078 6349 12124
rect 6395 12078 6507 12124
rect 6553 12078 6665 12124
rect 6711 12078 6823 12124
rect 6869 12078 6982 12124
rect 7028 12078 7140 12124
rect 7186 12078 7298 12124
rect 7344 12078 7456 12124
rect 7502 12078 7614 12124
rect 7660 12078 7772 12124
rect 7818 12078 7930 12124
rect 7976 12078 8089 12124
rect 8135 12078 8247 12124
rect 8293 12078 8405 12124
rect 8451 12078 8563 12124
rect 8609 12078 8664 12124
rect 5994 12011 8664 12078
rect 5994 11965 6038 12011
rect 6084 12007 8664 12011
rect 13588 12128 13632 12174
rect 13678 12128 13722 12174
rect 13588 12011 13722 12128
rect 13588 12007 13632 12011
rect 6084 11965 13632 12007
rect 13678 11965 13722 12011
rect 5994 11961 13722 11965
rect 5994 11915 6192 11961
rect 6238 11915 6350 11961
rect 6396 11915 6508 11961
rect 6554 11915 6666 11961
rect 6712 11915 6824 11961
rect 6870 11915 6982 11961
rect 7028 11915 7140 11961
rect 7186 11915 7298 11961
rect 7344 11915 7457 11961
rect 7503 11915 7615 11961
rect 7661 11915 7773 11961
rect 7819 11915 7931 11961
rect 7977 11915 8089 11961
rect 8135 11915 8247 11961
rect 8293 11915 8405 11961
rect 8451 11915 8563 11961
rect 8609 11915 8721 11961
rect 8767 11915 8880 11961
rect 8926 11915 9038 11961
rect 9084 11915 9196 11961
rect 9242 11915 9354 11961
rect 9400 11915 9512 11961
rect 9558 11915 9670 11961
rect 9716 11915 9828 11961
rect 9874 11915 9986 11961
rect 10032 11915 10144 11961
rect 10190 11915 10303 11961
rect 10349 11915 10461 11961
rect 10507 11915 10619 11961
rect 10665 11915 10777 11961
rect 10823 11915 10935 11961
rect 10981 11915 11093 11961
rect 11139 11915 11251 11961
rect 11297 11915 11409 11961
rect 11455 11915 11567 11961
rect 11613 11915 11726 11961
rect 11772 11915 11884 11961
rect 11930 11915 12042 11961
rect 12088 11915 12200 11961
rect 12246 11915 12358 11961
rect 12404 11915 12516 11961
rect 12562 11915 12674 11961
rect 12720 11915 12832 11961
rect 12878 11915 12990 11961
rect 13036 11915 13149 11961
rect 13195 11915 13307 11961
rect 13353 11915 13465 11961
rect 13511 11915 13722 11961
rect 5994 11869 13722 11915
rect 8927 9495 13511 9552
rect 8927 9449 8982 9495
rect 9028 9449 9140 9495
rect 9186 9449 9299 9495
rect 9345 9449 9457 9495
rect 9503 9449 9615 9495
rect 9661 9449 9773 9495
rect 9819 9449 9931 9495
rect 9977 9449 10089 9495
rect 10135 9449 10247 9495
rect 10293 9449 10405 9495
rect 10451 9449 10563 9495
rect 10609 9449 10722 9495
rect 10768 9449 10880 9495
rect 10926 9449 11038 9495
rect 11084 9449 11196 9495
rect 11242 9449 11354 9495
rect 11400 9449 11512 9495
rect 11558 9449 11671 9495
rect 11717 9449 11829 9495
rect 11875 9449 11987 9495
rect 12033 9449 12145 9495
rect 12191 9449 12303 9495
rect 12349 9449 12461 9495
rect 12507 9449 12619 9495
rect 12665 9449 12777 9495
rect 12823 9449 12935 9495
rect 12981 9449 13094 9495
rect 13140 9449 13252 9495
rect 13298 9449 13410 9495
rect 13456 9449 13511 9495
rect 8927 9392 13511 9449
rect 8927 9332 9241 9392
rect 8927 9286 8982 9332
rect 9028 9286 9140 9332
rect 9186 9286 9241 9332
rect 8927 9169 9241 9286
rect 13197 9332 13511 9392
rect 13197 9286 13252 9332
rect 13298 9286 13410 9332
rect 13456 9286 13511 9332
rect 8927 9123 8982 9169
rect 9028 9123 9140 9169
rect 9186 9123 9241 9169
rect 8927 9006 9241 9123
rect 8927 8960 8982 9006
rect 9028 8960 9140 9006
rect 9186 8960 9241 9006
rect 8927 8842 9241 8960
rect 8927 8796 8982 8842
rect 9028 8796 9140 8842
rect 9186 8796 9241 8842
rect 8927 8679 9241 8796
rect 8927 8633 8982 8679
rect 9028 8633 9140 8679
rect 9186 8633 9241 8679
rect 8927 8516 9241 8633
rect 8927 8470 8982 8516
rect 9028 8470 9140 8516
rect 9186 8470 9241 8516
rect 8927 8353 9241 8470
rect 8927 8307 8982 8353
rect 9028 8307 9140 8353
rect 9186 8307 9241 8353
rect 8927 8190 9241 8307
rect 8927 8144 8982 8190
rect 9028 8144 9140 8190
rect 9186 8144 9241 8190
rect 8927 8026 9241 8144
rect 8927 7980 8982 8026
rect 9028 7980 9140 8026
rect 9186 7980 9241 8026
rect 8927 7863 9241 7980
rect 8927 7817 8982 7863
rect 9028 7817 9140 7863
rect 9186 7817 9241 7863
rect 685 6914 4476 6972
rect 685 6868 739 6914
rect 785 6868 897 6914
rect 943 6868 1055 6914
rect 1101 6868 1213 6914
rect 1259 6868 1371 6914
rect 1417 6868 1529 6914
rect 1575 6868 1687 6914
rect 1733 6868 1845 6914
rect 1891 6868 2003 6914
rect 2049 6868 2162 6914
rect 2208 6868 2320 6914
rect 2366 6868 2478 6914
rect 2524 6868 2636 6914
rect 2682 6868 2794 6914
rect 2840 6868 2952 6914
rect 2998 6868 3111 6914
rect 3157 6868 3269 6914
rect 3315 6868 3427 6914
rect 3473 6868 3585 6914
rect 3631 6868 3743 6914
rect 3789 6868 3901 6914
rect 3947 6868 4059 6914
rect 4105 6868 4217 6914
rect 4263 6868 4375 6914
rect 4421 6868 4476 6914
rect 685 6751 4476 6868
rect 685 6705 739 6751
rect 785 6705 897 6751
rect 943 6705 1055 6751
rect 1101 6705 1213 6751
rect 1259 6705 1371 6751
rect 1417 6705 1529 6751
rect 1575 6705 1687 6751
rect 1733 6705 1845 6751
rect 1891 6705 2003 6751
rect 2049 6705 2162 6751
rect 2208 6705 2320 6751
rect 2366 6705 2478 6751
rect 2524 6705 2636 6751
rect 2682 6705 2794 6751
rect 2840 6705 2952 6751
rect 2998 6705 3111 6751
rect 3157 6705 3269 6751
rect 3315 6705 3427 6751
rect 3473 6705 3585 6751
rect 3631 6705 3743 6751
rect 3789 6705 3901 6751
rect 3947 6705 4059 6751
rect 4105 6705 4217 6751
rect 4263 6705 4375 6751
rect 4421 6705 4476 6751
rect 685 6588 4476 6705
rect 6339 6969 6473 7045
rect 6339 6923 6383 6969
rect 6429 6923 6473 6969
rect 6339 6777 6473 6923
rect 6339 6731 6383 6777
rect 6429 6731 6473 6777
rect 685 6542 739 6588
rect 785 6542 897 6588
rect 943 6542 1055 6588
rect 1101 6542 1213 6588
rect 1259 6542 1371 6588
rect 1417 6542 1529 6588
rect 1575 6542 1687 6588
rect 1733 6542 1845 6588
rect 1891 6542 2003 6588
rect 2049 6542 2162 6588
rect 2208 6542 2320 6588
rect 2366 6542 2478 6588
rect 2524 6542 2636 6588
rect 2682 6542 2794 6588
rect 2840 6542 2952 6588
rect 2998 6542 3111 6588
rect 3157 6542 3269 6588
rect 3315 6542 3427 6588
rect 3473 6542 3585 6588
rect 3631 6542 3743 6588
rect 3789 6542 3901 6588
rect 3947 6542 4059 6588
rect 4105 6542 4217 6588
rect 4263 6542 4375 6588
rect 4421 6542 4476 6588
rect 685 6485 4476 6542
rect 6339 6584 6473 6731
rect 6339 6538 6383 6584
rect 6429 6538 6473 6584
rect 6339 6421 6473 6538
rect 6339 6375 6383 6421
rect 6429 6375 6473 6421
rect 6339 6213 6473 6375
rect 8927 7700 9241 7817
rect 8927 7654 8982 7700
rect 9028 7654 9140 7700
rect 9186 7654 9241 7700
rect 8927 7536 9241 7654
rect 8927 7490 8982 7536
rect 9028 7490 9140 7536
rect 9186 7490 9241 7536
rect 8927 7373 9241 7490
rect 8927 7327 8982 7373
rect 9028 7327 9140 7373
rect 9186 7327 9241 7373
rect 8927 7210 9241 7327
rect 8927 7164 8982 7210
rect 9028 7164 9140 7210
rect 9186 7164 9241 7210
rect 8927 7046 9241 7164
rect 8927 7000 8982 7046
rect 9028 7000 9140 7046
rect 9186 7000 9241 7046
rect 8927 6883 9241 7000
rect 8927 6837 8982 6883
rect 9028 6837 9140 6883
rect 9186 6837 9241 6883
rect 8927 6720 9241 6837
rect 8927 6674 8982 6720
rect 9028 6674 9140 6720
rect 9186 6674 9241 6720
rect 8927 6557 9241 6674
rect 8927 6511 8982 6557
rect 9028 6511 9140 6557
rect 9186 6511 9241 6557
rect 8927 6394 9241 6511
rect 8927 6348 8982 6394
rect 9028 6348 9140 6394
rect 9186 6348 9241 6394
rect 8927 6230 9241 6348
rect 8927 6184 8982 6230
rect 9028 6184 9140 6230
rect 9186 6184 9241 6230
rect 8927 6067 9241 6184
rect 8927 6021 8982 6067
rect 9028 6021 9140 6067
rect 9186 6021 9241 6067
rect 8927 5904 9241 6021
rect 8927 5858 8982 5904
rect 9028 5858 9140 5904
rect 9186 5858 9241 5904
rect 8927 5741 9241 5858
rect 8927 5695 8982 5741
rect 9028 5695 9140 5741
rect 9186 5695 9241 5741
rect 8927 5638 9241 5695
rect 3753 2719 7433 2738
rect 3753 2673 3772 2719
rect 3818 2673 3896 2719
rect 3942 2673 4020 2719
rect 4066 2673 4144 2719
rect 4190 2673 4268 2719
rect 4314 2673 4392 2719
rect 4438 2673 4516 2719
rect 4562 2673 4640 2719
rect 4686 2673 4764 2719
rect 4810 2673 4888 2719
rect 4934 2673 5012 2719
rect 5058 2673 5136 2719
rect 5182 2673 5260 2719
rect 5306 2673 5384 2719
rect 5430 2673 5508 2719
rect 5554 2673 5632 2719
rect 5678 2673 5756 2719
rect 5802 2673 5880 2719
rect 5926 2673 6004 2719
rect 6050 2673 6128 2719
rect 6174 2673 6252 2719
rect 6298 2673 6376 2719
rect 6422 2673 6500 2719
rect 6546 2673 6624 2719
rect 6670 2673 6748 2719
rect 6794 2673 6872 2719
rect 6918 2673 6996 2719
rect 7042 2673 7120 2719
rect 7166 2673 7244 2719
rect 7290 2673 7368 2719
rect 7414 2673 7433 2719
rect 3753 2595 7433 2673
rect 3753 2549 3772 2595
rect 3818 2549 3896 2595
rect 3942 2549 4020 2595
rect 4066 2549 4144 2595
rect 4190 2549 4268 2595
rect 4314 2549 4392 2595
rect 4438 2549 4516 2595
rect 4562 2549 4640 2595
rect 4686 2549 4764 2595
rect 4810 2549 4888 2595
rect 4934 2549 5012 2595
rect 5058 2549 5136 2595
rect 5182 2549 5260 2595
rect 5306 2549 5384 2595
rect 5430 2549 5508 2595
rect 5554 2549 5632 2595
rect 5678 2549 5756 2595
rect 5802 2549 5880 2595
rect 5926 2549 6004 2595
rect 6050 2549 6128 2595
rect 6174 2549 6252 2595
rect 6298 2549 6376 2595
rect 6422 2549 6500 2595
rect 6546 2549 6624 2595
rect 6670 2549 6748 2595
rect 6794 2549 6872 2595
rect 6918 2549 6996 2595
rect 7042 2549 7120 2595
rect 7166 2549 7244 2595
rect 7290 2549 7368 2595
rect 7414 2549 7433 2595
rect 3753 2471 7433 2549
rect 3753 2425 3772 2471
rect 3818 2425 3896 2471
rect 3942 2425 4020 2471
rect 4066 2425 4144 2471
rect 4190 2425 4268 2471
rect 4314 2425 4392 2471
rect 4438 2425 4516 2471
rect 4562 2425 4640 2471
rect 4686 2425 4764 2471
rect 4810 2425 4888 2471
rect 4934 2425 5012 2471
rect 5058 2425 5136 2471
rect 5182 2425 5260 2471
rect 5306 2425 5384 2471
rect 5430 2425 5508 2471
rect 5554 2425 5632 2471
rect 5678 2425 5756 2471
rect 5802 2425 5880 2471
rect 5926 2425 6004 2471
rect 6050 2425 6128 2471
rect 6174 2425 6252 2471
rect 6298 2425 6376 2471
rect 6422 2425 6500 2471
rect 6546 2425 6624 2471
rect 6670 2425 6748 2471
rect 6794 2425 6872 2471
rect 6918 2425 6996 2471
rect 7042 2425 7120 2471
rect 7166 2425 7244 2471
rect 7290 2425 7368 2471
rect 7414 2425 7433 2471
rect 3753 2347 7433 2425
rect 3753 2301 3772 2347
rect 3818 2301 3896 2347
rect 3942 2301 4020 2347
rect 4066 2301 4144 2347
rect 4190 2301 4268 2347
rect 4314 2301 4392 2347
rect 4438 2301 4516 2347
rect 4562 2301 4640 2347
rect 4686 2301 4764 2347
rect 4810 2301 4888 2347
rect 4934 2301 5012 2347
rect 5058 2301 5136 2347
rect 5182 2301 5260 2347
rect 5306 2301 5384 2347
rect 5430 2301 5508 2347
rect 5554 2301 5632 2347
rect 5678 2301 5756 2347
rect 5802 2301 5880 2347
rect 5926 2301 6004 2347
rect 6050 2301 6128 2347
rect 6174 2301 6252 2347
rect 6298 2301 6376 2347
rect 6422 2301 6500 2347
rect 6546 2301 6624 2347
rect 6670 2301 6748 2347
rect 6794 2301 6872 2347
rect 6918 2301 6996 2347
rect 7042 2301 7120 2347
rect 7166 2301 7244 2347
rect 7290 2301 7368 2347
rect 7414 2301 7433 2347
rect 3753 2282 7433 2301
rect 13197 9169 13511 9286
rect 13197 9123 13252 9169
rect 13298 9123 13410 9169
rect 13456 9123 13511 9169
rect 13197 9006 13511 9123
rect 13197 8960 13252 9006
rect 13298 8960 13410 9006
rect 13456 8960 13511 9006
rect 13197 8843 13511 8960
rect 13197 8797 13252 8843
rect 13298 8797 13410 8843
rect 13456 8797 13511 8843
rect 13197 8679 13511 8797
rect 13197 8633 13252 8679
rect 13298 8633 13410 8679
rect 13456 8633 13511 8679
rect 13197 8516 13511 8633
rect 13197 8470 13252 8516
rect 13298 8470 13410 8516
rect 13456 8470 13511 8516
rect 13197 8353 13511 8470
rect 13197 8307 13252 8353
rect 13298 8307 13410 8353
rect 13456 8307 13511 8353
rect 13197 8190 13511 8307
rect 13197 8144 13252 8190
rect 13298 8144 13410 8190
rect 13456 8144 13511 8190
rect 13197 8026 13511 8144
rect 13197 7980 13252 8026
rect 13298 7980 13410 8026
rect 13456 7980 13511 8026
rect 13197 7863 13511 7980
rect 13197 7817 13252 7863
rect 13298 7817 13410 7863
rect 13456 7817 13511 7863
rect 13197 7700 13511 7817
rect 13197 7654 13252 7700
rect 13298 7654 13410 7700
rect 13456 7654 13511 7700
rect 13197 7537 13511 7654
rect 13197 7491 13252 7537
rect 13298 7491 13410 7537
rect 13456 7491 13511 7537
rect 13197 7373 13511 7491
rect 13197 7327 13252 7373
rect 13298 7327 13410 7373
rect 13456 7327 13511 7373
rect 13197 7210 13511 7327
rect 13197 7164 13252 7210
rect 13298 7164 13410 7210
rect 13456 7164 13511 7210
rect 13197 7047 13511 7164
rect 13197 7001 13252 7047
rect 13298 7001 13410 7047
rect 13456 7001 13511 7047
rect 13197 6883 13511 7001
rect 13197 6837 13252 6883
rect 13298 6837 13410 6883
rect 13456 6837 13511 6883
rect 13197 6720 13511 6837
rect 13197 6674 13252 6720
rect 13298 6674 13410 6720
rect 13456 6674 13511 6720
rect 13197 6557 13511 6674
rect 13197 6511 13252 6557
rect 13298 6511 13410 6557
rect 13456 6511 13511 6557
rect 13197 6394 13511 6511
rect 13197 6348 13252 6394
rect 13298 6348 13410 6394
rect 13456 6348 13511 6394
rect 13197 6230 13511 6348
rect 13197 6184 13252 6230
rect 13298 6184 13410 6230
rect 13456 6184 13511 6230
rect 13197 6067 13511 6184
rect 13197 6021 13252 6067
rect 13298 6021 13410 6067
rect 13456 6021 13511 6067
rect 13197 5904 13511 6021
rect 13197 5858 13252 5904
rect 13298 5858 13410 5904
rect 13456 5858 13511 5904
rect 13197 5741 13511 5858
rect 13197 5695 13252 5741
rect 13298 5695 13410 5741
rect 13456 5695 13511 5741
rect 13197 5577 13511 5695
rect 13197 5531 13252 5577
rect 13298 5531 13410 5577
rect 13456 5531 13511 5577
rect 13197 5414 13511 5531
rect 13197 5368 13252 5414
rect 13298 5368 13410 5414
rect 13456 5368 13511 5414
rect 13197 5251 13511 5368
rect 13197 5205 13252 5251
rect 13298 5205 13410 5251
rect 13456 5205 13511 5251
rect 13197 5088 13511 5205
rect 13197 5042 13252 5088
rect 13298 5042 13410 5088
rect 13456 5042 13511 5088
rect 13197 4925 13511 5042
rect 13197 4879 13252 4925
rect 13298 4879 13410 4925
rect 13456 4879 13511 4925
rect 13197 4822 13511 4879
<< mvpsubdiffcont >>
rect 13643 11550 13689 11596
rect 6323 11432 6369 11478
rect 6481 11432 6527 11478
rect 6639 11432 6685 11478
rect 6798 11432 6844 11478
rect 6956 11432 7002 11478
rect 7114 11432 7160 11478
rect 7272 11432 7318 11478
rect 7430 11432 7476 11478
rect 7588 11432 7634 11478
rect 7747 11432 7793 11478
rect 7905 11432 7951 11478
rect 8063 11432 8109 11478
rect 6323 11269 6369 11315
rect 13643 11387 13689 11433
rect 8045 11197 8091 11243
rect 8203 11197 8249 11243
rect 6323 11106 6369 11152
rect 6323 10942 6369 10988
rect 6323 10779 6369 10825
rect 6323 10616 6369 10662
rect 6323 10453 6369 10499
rect 6323 10289 6369 10335
rect 6323 10126 6369 10172
rect 6323 9963 6369 10009
rect 6323 9799 6369 9845
rect 6323 9636 6369 9682
rect 6323 9473 6369 9519
rect 6323 9310 6369 9356
rect 6323 9146 6369 9192
rect 8045 11034 8091 11080
rect 8203 11034 8249 11080
rect 8045 10871 8091 10917
rect 8203 10871 8249 10917
rect 8045 10707 8091 10753
rect 8203 10707 8249 10753
rect 8045 10544 8091 10590
rect 8203 10544 8249 10590
rect 8045 10381 8091 10427
rect 8203 10381 8249 10427
rect 8045 10218 8091 10264
rect 8203 10218 8249 10264
rect 8045 10054 8091 10100
rect 8203 10054 8249 10100
rect 8045 9891 8091 9937
rect 8203 9891 8249 9937
rect 13643 11224 13689 11270
rect 13643 11061 13689 11107
rect 13643 10897 13689 10943
rect 13643 10734 13689 10780
rect 13643 10571 13689 10617
rect 13643 10407 13689 10453
rect 13643 10244 13689 10290
rect 13643 10081 13689 10127
rect 13643 9918 13689 9964
rect 8045 9728 8091 9774
rect 8203 9728 8249 9774
rect 8045 9564 8091 9610
rect 8203 9564 8249 9610
rect 8045 9401 8091 9447
rect 8203 9401 8249 9447
rect 8045 9238 8091 9284
rect 8203 9238 8249 9284
rect 8045 9075 8091 9121
rect 8203 9075 8249 9121
rect 6323 8983 6369 9029
rect 6323 8820 6369 8866
rect 8045 8911 8091 8957
rect 8203 8911 8249 8957
rect 8045 8748 8091 8794
rect 8203 8748 8249 8794
rect 400 8585 446 8631
rect 558 8585 604 8631
rect 716 8585 762 8631
rect 875 8585 921 8631
rect 1033 8585 1079 8631
rect 1191 8585 1237 8631
rect 1349 8585 1395 8631
rect 1507 8585 1553 8631
rect 1665 8585 1711 8631
rect 1823 8585 1869 8631
rect 1981 8585 2027 8631
rect 2139 8585 2185 8631
rect 2298 8585 2344 8631
rect 2456 8585 2502 8631
rect 2614 8585 2660 8631
rect 2772 8585 2818 8631
rect 2930 8585 2976 8631
rect 3088 8585 3134 8631
rect 3246 8585 3292 8631
rect 3404 8585 3450 8631
rect 3562 8585 3608 8631
rect 3721 8585 3767 8631
rect 3879 8585 3925 8631
rect 4037 8585 4083 8631
rect 4195 8585 4241 8631
rect 4353 8585 4399 8631
rect 4511 8585 4557 8631
rect 4670 8585 4716 8631
rect 4828 8585 4874 8631
rect 4986 8585 5032 8631
rect 5144 8585 5190 8631
rect 5302 8585 5348 8631
rect 5460 8585 5506 8631
rect 5618 8585 5664 8631
rect 5776 8585 5822 8631
rect 5934 8585 5980 8631
rect 6093 8585 6139 8631
rect 6251 8585 6297 8631
rect 6409 8585 6455 8631
rect 6567 8585 6613 8631
rect 6725 8585 6771 8631
rect 6883 8585 6929 8631
rect 7041 8585 7087 8631
rect 7199 8585 7245 8631
rect 7357 8585 7403 8631
rect 7516 8585 7562 8631
rect 7674 8585 7720 8631
rect 7832 8585 7878 8631
rect 8045 8585 8091 8631
rect 8203 8585 8249 8631
rect 403 8260 449 8306
rect 561 8260 607 8306
rect 719 8260 765 8306
rect 877 8260 923 8306
rect 1035 8260 1081 8306
rect 1193 8260 1239 8306
rect 1351 8260 1397 8306
rect 1509 8260 1555 8306
rect 1667 8260 1713 8306
rect 1826 8260 1872 8306
rect 1984 8260 2030 8306
rect 2142 8260 2188 8306
rect 2300 8260 2346 8306
rect 2458 8260 2504 8306
rect 2616 8260 2662 8306
rect 2774 8260 2820 8306
rect 2933 8260 2979 8306
rect 3091 8260 3137 8306
rect 3249 8260 3295 8306
rect 3407 8260 3453 8306
rect 3565 8260 3611 8306
rect 3723 8260 3769 8306
rect 3881 8260 3927 8306
rect 4039 8260 4085 8306
rect 4197 8260 4243 8306
rect 403 8097 449 8143
rect 561 8097 607 8143
rect 719 8097 765 8143
rect 877 8097 923 8143
rect 1035 8097 1081 8143
rect 1193 8097 1239 8143
rect 1351 8097 1397 8143
rect 1509 8097 1555 8143
rect 1667 8097 1713 8143
rect 1826 8097 1872 8143
rect 1984 8097 2030 8143
rect 2142 8097 2188 8143
rect 2300 8097 2346 8143
rect 2458 8097 2504 8143
rect 2616 8097 2662 8143
rect 2774 8097 2820 8143
rect 2933 8097 2979 8143
rect 3091 8097 3137 8143
rect 3249 8097 3295 8143
rect 3407 8097 3453 8143
rect 3565 8097 3611 8143
rect 3723 8097 3769 8143
rect 3881 8097 3927 8143
rect 4039 8097 4085 8143
rect 4197 8097 4243 8143
rect 403 7934 449 7980
rect 561 7934 607 7980
rect 719 7934 765 7980
rect 877 7934 923 7980
rect 1035 7934 1081 7980
rect 1193 7934 1239 7980
rect 1351 7934 1397 7980
rect 1509 7934 1555 7980
rect 1667 7934 1713 7980
rect 1826 7934 1872 7980
rect 1984 7934 2030 7980
rect 2142 7934 2188 7980
rect 2300 7934 2346 7980
rect 2458 7934 2504 7980
rect 2616 7934 2662 7980
rect 2774 7934 2820 7980
rect 2933 7934 2979 7980
rect 3091 7934 3137 7980
rect 3249 7934 3295 7980
rect 3407 7934 3453 7980
rect 3565 7934 3611 7980
rect 3723 7934 3769 7980
rect 3881 7934 3927 7980
rect 4039 7934 4085 7980
rect 4197 7934 4243 7980
rect 739 5885 785 5931
rect 897 5885 943 5931
rect 1055 5885 1101 5931
rect 1213 5885 1259 5931
rect 1371 5885 1417 5931
rect 1529 5885 1575 5931
rect 1687 5885 1733 5931
rect 1845 5885 1891 5931
rect 2003 5885 2049 5931
rect 2162 5885 2208 5931
rect 2320 5885 2366 5931
rect 2478 5885 2524 5931
rect 2636 5885 2682 5931
rect 2794 5885 2840 5931
rect 2952 5885 2998 5931
rect 3111 5885 3157 5931
rect 3269 5885 3315 5931
rect 3427 5885 3473 5931
rect 3585 5885 3631 5931
rect 3743 5885 3789 5931
rect 3901 5885 3947 5931
rect 4059 5885 4105 5931
rect 4217 5885 4263 5931
rect 4375 5885 4421 5931
rect 739 5722 785 5768
rect 897 5722 943 5768
rect 1055 5722 1101 5768
rect 1213 5722 1259 5768
rect 1371 5722 1417 5768
rect 1529 5722 1575 5768
rect 1687 5722 1733 5768
rect 1845 5722 1891 5768
rect 2003 5722 2049 5768
rect 2162 5722 2208 5768
rect 2320 5722 2366 5768
rect 2478 5722 2524 5768
rect 2636 5722 2682 5768
rect 2794 5722 2840 5768
rect 2952 5722 2998 5768
rect 3111 5722 3157 5768
rect 3269 5722 3315 5768
rect 3427 5722 3473 5768
rect 3585 5722 3631 5768
rect 3743 5722 3789 5768
rect 3901 5722 3947 5768
rect 4059 5722 4105 5768
rect 4217 5722 4263 5768
rect 4375 5722 4421 5768
rect 739 5559 785 5605
rect 897 5559 943 5605
rect 1055 5559 1101 5605
rect 1213 5559 1259 5605
rect 1371 5559 1417 5605
rect 1529 5559 1575 5605
rect 1687 5559 1733 5605
rect 1845 5559 1891 5605
rect 2003 5559 2049 5605
rect 2162 5559 2208 5605
rect 2320 5559 2366 5605
rect 2478 5559 2524 5605
rect 2636 5559 2682 5605
rect 2794 5559 2840 5605
rect 2952 5559 2998 5605
rect 3111 5559 3157 5605
rect 3269 5559 3315 5605
rect 3427 5559 3473 5605
rect 3585 5559 3631 5605
rect 3743 5559 3789 5605
rect 3901 5559 3947 5605
rect 4059 5559 4105 5605
rect 4217 5559 4263 5605
rect 4375 5559 4421 5605
rect 6383 5661 6429 5707
rect 6383 5497 6429 5543
rect 314 4351 7760 4997
rect 8926 4674 8972 4720
rect 9084 4674 9130 4720
rect 8926 4511 8972 4557
rect 9084 4511 9130 4557
rect 8926 4348 8972 4394
rect 9084 4348 9130 4394
rect 8926 4184 8972 4230
rect 9084 4184 9130 4230
rect 8926 4021 8972 4067
rect 9084 4021 9130 4067
rect 8926 3858 8972 3904
rect 9084 3858 9130 3904
rect 8926 3695 8972 3741
rect 9084 3695 9130 3741
rect 8926 3531 8972 3577
rect 9084 3531 9130 3577
rect 8926 3368 8972 3414
rect 9084 3368 9130 3414
rect 8926 3205 8972 3251
rect 9084 3205 9130 3251
rect 8926 3042 8972 3088
rect 9084 3042 9130 3088
rect 8926 2879 8972 2925
rect 9084 2879 9130 2925
rect 8926 2715 8972 2761
rect 9084 2715 9130 2761
rect 8926 2552 8972 2598
rect 9084 2552 9130 2598
rect 8926 2389 8972 2435
rect 9084 2389 9130 2435
rect 8926 2225 8972 2271
rect 9084 2225 9130 2271
rect 8926 2062 8972 2108
rect 9084 2062 9130 2108
rect 8926 1899 8972 1945
rect 9084 1899 9130 1945
rect 8926 1735 8972 1781
rect 9084 1735 9130 1781
rect 8926 1572 8972 1618
rect 9084 1572 9130 1618
rect 8926 1409 8972 1455
rect 9084 1409 9130 1455
rect 8926 1246 8972 1292
rect 9084 1246 9130 1292
rect 8926 1083 8972 1129
rect 9084 1083 9130 1129
rect 8926 919 8972 965
rect 9084 919 9130 965
rect 8926 756 8972 802
rect 9084 756 9130 802
rect 8926 593 8972 639
rect 9084 593 9130 639
rect 8926 430 8972 476
rect 9084 430 9130 476
rect 8926 266 8972 312
rect 9084 266 9130 312
rect 13353 4191 13399 4237
rect 13511 4191 13557 4237
rect 13353 4028 13399 4074
rect 13511 4028 13557 4074
rect 13353 3859 13399 3905
rect 13511 3859 13557 3905
rect 13353 3696 13399 3742
rect 13511 3696 13557 3742
rect 13353 3532 13399 3578
rect 13511 3532 13557 3578
rect 13353 3369 13399 3415
rect 13511 3369 13557 3415
rect 13353 3206 13399 3252
rect 13511 3206 13557 3252
rect 13353 3043 13399 3089
rect 13511 3043 13557 3089
rect 13353 2879 13399 2925
rect 13511 2879 13557 2925
rect 13353 2716 13399 2762
rect 13511 2716 13557 2762
rect 13353 2553 13399 2599
rect 13511 2553 13557 2599
rect 13353 2390 13399 2436
rect 13511 2390 13557 2436
rect 13353 2226 13399 2272
rect 13511 2226 13557 2272
rect 13353 2063 13399 2109
rect 13511 2063 13557 2109
rect 13353 1900 13399 1946
rect 13511 1900 13557 1946
rect 13353 1736 13399 1782
rect 13511 1736 13557 1782
rect 13353 1573 13399 1619
rect 13511 1573 13557 1619
rect 13353 1410 13399 1456
rect 13511 1410 13557 1456
rect 13353 1247 13399 1293
rect 13511 1247 13557 1293
rect 13353 1083 13399 1129
rect 13511 1083 13557 1129
rect 13353 920 13399 966
rect 13511 920 13557 966
rect 13353 757 13399 803
rect 13511 757 13557 803
rect 13353 594 13399 640
rect 13511 594 13557 640
rect 13353 430 13399 476
rect 13511 430 13557 476
rect 13353 267 13399 313
rect 13511 267 13557 313
rect 8926 103 8972 149
rect 9084 103 9130 149
rect 13353 104 13399 150
rect 13511 104 13557 150
rect 8926 -60 8972 -14
rect 9084 -60 9130 -14
rect 9401 -60 9447 -14
rect 9559 -60 9605 -14
rect 9717 -60 9763 -14
rect 9875 -60 9921 -14
rect 10033 -60 10079 -14
rect 10191 -60 10237 -14
rect 10349 -60 10395 -14
rect 10507 -60 10553 -14
rect 10665 -60 10711 -14
rect 10824 -60 10870 -14
rect 10982 -60 11028 -14
rect 11140 -60 11186 -14
rect 11298 -60 11344 -14
rect 11456 -60 11502 -14
rect 11614 -60 11660 -14
rect 11772 -60 11818 -14
rect 11931 -60 11977 -14
rect 12089 -60 12135 -14
rect 12247 -60 12293 -14
rect 12405 -60 12451 -14
rect 12563 -60 12609 -14
rect 12721 -60 12767 -14
rect 12879 -60 12925 -14
rect 13037 -60 13083 -14
rect 13195 -60 13241 -14
rect 13353 -59 13399 -13
rect 13511 -59 13557 -13
<< mvnsubdiffcont >>
rect 6192 16227 6238 16273
rect 6350 16227 6396 16273
rect 6508 16227 6554 16273
rect 6666 16227 6712 16273
rect 6824 16227 6870 16273
rect 6982 16227 7028 16273
rect 7140 16227 7186 16273
rect 7298 16227 7344 16273
rect 7457 16227 7503 16273
rect 7615 16227 7661 16273
rect 7773 16227 7819 16273
rect 7931 16227 7977 16273
rect 8089 16227 8135 16273
rect 8247 16227 8293 16273
rect 8405 16227 8451 16273
rect 8563 16227 8609 16273
rect 8721 16227 8767 16273
rect 8880 16227 8926 16273
rect 9038 16227 9084 16273
rect 9196 16227 9242 16273
rect 9354 16227 9400 16273
rect 9512 16227 9558 16273
rect 9670 16227 9716 16273
rect 9828 16227 9874 16273
rect 9986 16227 10032 16273
rect 10144 16227 10190 16273
rect 10303 16227 10349 16273
rect 10461 16227 10507 16273
rect 10619 16227 10665 16273
rect 10777 16227 10823 16273
rect 10935 16227 10981 16273
rect 11093 16227 11139 16273
rect 11251 16227 11297 16273
rect 11409 16227 11455 16273
rect 11567 16227 11613 16273
rect 11726 16227 11772 16273
rect 11884 16227 11930 16273
rect 12042 16227 12088 16273
rect 12200 16227 12246 16273
rect 12358 16227 12404 16273
rect 12516 16227 12562 16273
rect 12674 16227 12720 16273
rect 12832 16227 12878 16273
rect 12990 16227 13036 16273
rect 13149 16227 13195 16273
rect 13307 16227 13353 16273
rect 13465 16227 13511 16273
rect 6038 16046 6084 16092
rect 13632 16046 13678 16092
rect 6038 15882 6084 15928
rect 6038 15719 6084 15765
rect 6038 15556 6084 15602
rect 6038 15393 6084 15439
rect 6038 15229 6084 15275
rect 6038 15066 6084 15112
rect 6038 14903 6084 14949
rect 6038 14740 6084 14786
rect 6038 14576 6084 14622
rect 6038 14413 6084 14459
rect 6038 14250 6084 14296
rect 6038 14087 6084 14133
rect 6038 13924 6084 13970
rect 6038 13760 6084 13806
rect 6038 13597 6084 13643
rect 6038 13434 6084 13480
rect 6038 13271 6084 13317
rect 6038 13107 6084 13153
rect 6349 13058 6395 13104
rect 6507 13058 6553 13104
rect 6665 13058 6711 13104
rect 6823 13058 6869 13104
rect 6982 13058 7028 13104
rect 7140 13058 7186 13104
rect 7298 13058 7344 13104
rect 7456 13058 7502 13104
rect 7614 13058 7660 13104
rect 7772 13058 7818 13104
rect 7930 13058 7976 13104
rect 8089 13058 8135 13104
rect 8247 13058 8293 13104
rect 8405 13058 8451 13104
rect 8563 13058 8609 13104
rect 6038 12944 6084 12990
rect 6349 12895 6395 12941
rect 6507 12895 6553 12941
rect 6665 12895 6711 12941
rect 6823 12895 6869 12941
rect 6982 12895 7028 12941
rect 7140 12895 7186 12941
rect 7298 12895 7344 12941
rect 7456 12895 7502 12941
rect 7614 12895 7660 12941
rect 7772 12895 7818 12941
rect 7930 12895 7976 12941
rect 8089 12895 8135 12941
rect 8247 12895 8293 12941
rect 8405 12895 8451 12941
rect 8563 12895 8609 12941
rect 6038 12781 6084 12827
rect 6349 12731 6395 12777
rect 6507 12731 6553 12777
rect 6665 12731 6711 12777
rect 6823 12731 6869 12777
rect 6982 12731 7028 12777
rect 7140 12731 7186 12777
rect 7298 12731 7344 12777
rect 7456 12731 7502 12777
rect 7614 12731 7660 12777
rect 7772 12731 7818 12777
rect 7930 12731 7976 12777
rect 8089 12731 8135 12777
rect 8247 12731 8293 12777
rect 8405 12731 8451 12777
rect 8563 12731 8609 12777
rect 6038 12618 6084 12664
rect 6349 12568 6395 12614
rect 6507 12568 6553 12614
rect 6665 12568 6711 12614
rect 6823 12568 6869 12614
rect 6982 12568 7028 12614
rect 7140 12568 7186 12614
rect 7298 12568 7344 12614
rect 7456 12568 7502 12614
rect 7614 12568 7660 12614
rect 7772 12568 7818 12614
rect 7930 12568 7976 12614
rect 8089 12568 8135 12614
rect 8247 12568 8293 12614
rect 8405 12568 8451 12614
rect 8563 12568 8609 12614
rect 6038 12455 6084 12501
rect 6349 12405 6395 12451
rect 6507 12405 6553 12451
rect 6665 12405 6711 12451
rect 6823 12405 6869 12451
rect 6982 12405 7028 12451
rect 7140 12405 7186 12451
rect 7298 12405 7344 12451
rect 7456 12405 7502 12451
rect 7614 12405 7660 12451
rect 7772 12405 7818 12451
rect 7930 12405 7976 12451
rect 8089 12405 8135 12451
rect 8247 12405 8293 12451
rect 8405 12405 8451 12451
rect 8563 12405 8609 12451
rect 6038 12291 6084 12337
rect 6349 12241 6395 12287
rect 6507 12241 6553 12287
rect 6665 12241 6711 12287
rect 6823 12241 6869 12287
rect 6982 12241 7028 12287
rect 7140 12241 7186 12287
rect 7298 12241 7344 12287
rect 7456 12241 7502 12287
rect 7614 12241 7660 12287
rect 7772 12241 7818 12287
rect 7930 12241 7976 12287
rect 8089 12241 8135 12287
rect 8247 12241 8293 12287
rect 8405 12241 8451 12287
rect 8563 12241 8609 12287
rect 13632 15882 13678 15928
rect 13632 15719 13678 15765
rect 13632 15556 13678 15602
rect 13632 15393 13678 15439
rect 13632 15229 13678 15275
rect 13632 15066 13678 15112
rect 13632 14903 13678 14949
rect 13632 14740 13678 14786
rect 13632 14576 13678 14622
rect 13632 14413 13678 14459
rect 13632 14250 13678 14296
rect 13632 14087 13678 14133
rect 13632 13924 13678 13970
rect 13632 13760 13678 13806
rect 13632 13597 13678 13643
rect 13632 13434 13678 13480
rect 13632 13271 13678 13317
rect 13632 13107 13678 13153
rect 13632 12944 13678 12990
rect 13632 12781 13678 12827
rect 13632 12618 13678 12664
rect 13632 12455 13678 12501
rect 13632 12291 13678 12337
rect 6038 12128 6084 12174
rect 6349 12078 6395 12124
rect 6507 12078 6553 12124
rect 6665 12078 6711 12124
rect 6823 12078 6869 12124
rect 6982 12078 7028 12124
rect 7140 12078 7186 12124
rect 7298 12078 7344 12124
rect 7456 12078 7502 12124
rect 7614 12078 7660 12124
rect 7772 12078 7818 12124
rect 7930 12078 7976 12124
rect 8089 12078 8135 12124
rect 8247 12078 8293 12124
rect 8405 12078 8451 12124
rect 8563 12078 8609 12124
rect 6038 11965 6084 12011
rect 13632 12128 13678 12174
rect 13632 11965 13678 12011
rect 6192 11915 6238 11961
rect 6350 11915 6396 11961
rect 6508 11915 6554 11961
rect 6666 11915 6712 11961
rect 6824 11915 6870 11961
rect 6982 11915 7028 11961
rect 7140 11915 7186 11961
rect 7298 11915 7344 11961
rect 7457 11915 7503 11961
rect 7615 11915 7661 11961
rect 7773 11915 7819 11961
rect 7931 11915 7977 11961
rect 8089 11915 8135 11961
rect 8247 11915 8293 11961
rect 8405 11915 8451 11961
rect 8563 11915 8609 11961
rect 8721 11915 8767 11961
rect 8880 11915 8926 11961
rect 9038 11915 9084 11961
rect 9196 11915 9242 11961
rect 9354 11915 9400 11961
rect 9512 11915 9558 11961
rect 9670 11915 9716 11961
rect 9828 11915 9874 11961
rect 9986 11915 10032 11961
rect 10144 11915 10190 11961
rect 10303 11915 10349 11961
rect 10461 11915 10507 11961
rect 10619 11915 10665 11961
rect 10777 11915 10823 11961
rect 10935 11915 10981 11961
rect 11093 11915 11139 11961
rect 11251 11915 11297 11961
rect 11409 11915 11455 11961
rect 11567 11915 11613 11961
rect 11726 11915 11772 11961
rect 11884 11915 11930 11961
rect 12042 11915 12088 11961
rect 12200 11915 12246 11961
rect 12358 11915 12404 11961
rect 12516 11915 12562 11961
rect 12674 11915 12720 11961
rect 12832 11915 12878 11961
rect 12990 11915 13036 11961
rect 13149 11915 13195 11961
rect 13307 11915 13353 11961
rect 13465 11915 13511 11961
rect 8982 9449 9028 9495
rect 9140 9449 9186 9495
rect 9299 9449 9345 9495
rect 9457 9449 9503 9495
rect 9615 9449 9661 9495
rect 9773 9449 9819 9495
rect 9931 9449 9977 9495
rect 10089 9449 10135 9495
rect 10247 9449 10293 9495
rect 10405 9449 10451 9495
rect 10563 9449 10609 9495
rect 10722 9449 10768 9495
rect 10880 9449 10926 9495
rect 11038 9449 11084 9495
rect 11196 9449 11242 9495
rect 11354 9449 11400 9495
rect 11512 9449 11558 9495
rect 11671 9449 11717 9495
rect 11829 9449 11875 9495
rect 11987 9449 12033 9495
rect 12145 9449 12191 9495
rect 12303 9449 12349 9495
rect 12461 9449 12507 9495
rect 12619 9449 12665 9495
rect 12777 9449 12823 9495
rect 12935 9449 12981 9495
rect 13094 9449 13140 9495
rect 13252 9449 13298 9495
rect 13410 9449 13456 9495
rect 8982 9286 9028 9332
rect 9140 9286 9186 9332
rect 13252 9286 13298 9332
rect 13410 9286 13456 9332
rect 8982 9123 9028 9169
rect 9140 9123 9186 9169
rect 8982 8960 9028 9006
rect 9140 8960 9186 9006
rect 8982 8796 9028 8842
rect 9140 8796 9186 8842
rect 8982 8633 9028 8679
rect 9140 8633 9186 8679
rect 8982 8470 9028 8516
rect 9140 8470 9186 8516
rect 8982 8307 9028 8353
rect 9140 8307 9186 8353
rect 8982 8144 9028 8190
rect 9140 8144 9186 8190
rect 8982 7980 9028 8026
rect 9140 7980 9186 8026
rect 8982 7817 9028 7863
rect 9140 7817 9186 7863
rect 739 6868 785 6914
rect 897 6868 943 6914
rect 1055 6868 1101 6914
rect 1213 6868 1259 6914
rect 1371 6868 1417 6914
rect 1529 6868 1575 6914
rect 1687 6868 1733 6914
rect 1845 6868 1891 6914
rect 2003 6868 2049 6914
rect 2162 6868 2208 6914
rect 2320 6868 2366 6914
rect 2478 6868 2524 6914
rect 2636 6868 2682 6914
rect 2794 6868 2840 6914
rect 2952 6868 2998 6914
rect 3111 6868 3157 6914
rect 3269 6868 3315 6914
rect 3427 6868 3473 6914
rect 3585 6868 3631 6914
rect 3743 6868 3789 6914
rect 3901 6868 3947 6914
rect 4059 6868 4105 6914
rect 4217 6868 4263 6914
rect 4375 6868 4421 6914
rect 739 6705 785 6751
rect 897 6705 943 6751
rect 1055 6705 1101 6751
rect 1213 6705 1259 6751
rect 1371 6705 1417 6751
rect 1529 6705 1575 6751
rect 1687 6705 1733 6751
rect 1845 6705 1891 6751
rect 2003 6705 2049 6751
rect 2162 6705 2208 6751
rect 2320 6705 2366 6751
rect 2478 6705 2524 6751
rect 2636 6705 2682 6751
rect 2794 6705 2840 6751
rect 2952 6705 2998 6751
rect 3111 6705 3157 6751
rect 3269 6705 3315 6751
rect 3427 6705 3473 6751
rect 3585 6705 3631 6751
rect 3743 6705 3789 6751
rect 3901 6705 3947 6751
rect 4059 6705 4105 6751
rect 4217 6705 4263 6751
rect 4375 6705 4421 6751
rect 6383 6923 6429 6969
rect 6383 6731 6429 6777
rect 739 6542 785 6588
rect 897 6542 943 6588
rect 1055 6542 1101 6588
rect 1213 6542 1259 6588
rect 1371 6542 1417 6588
rect 1529 6542 1575 6588
rect 1687 6542 1733 6588
rect 1845 6542 1891 6588
rect 2003 6542 2049 6588
rect 2162 6542 2208 6588
rect 2320 6542 2366 6588
rect 2478 6542 2524 6588
rect 2636 6542 2682 6588
rect 2794 6542 2840 6588
rect 2952 6542 2998 6588
rect 3111 6542 3157 6588
rect 3269 6542 3315 6588
rect 3427 6542 3473 6588
rect 3585 6542 3631 6588
rect 3743 6542 3789 6588
rect 3901 6542 3947 6588
rect 4059 6542 4105 6588
rect 4217 6542 4263 6588
rect 4375 6542 4421 6588
rect 6383 6538 6429 6584
rect 6383 6375 6429 6421
rect 8982 7654 9028 7700
rect 9140 7654 9186 7700
rect 8982 7490 9028 7536
rect 9140 7490 9186 7536
rect 8982 7327 9028 7373
rect 9140 7327 9186 7373
rect 8982 7164 9028 7210
rect 9140 7164 9186 7210
rect 8982 7000 9028 7046
rect 9140 7000 9186 7046
rect 8982 6837 9028 6883
rect 9140 6837 9186 6883
rect 8982 6674 9028 6720
rect 9140 6674 9186 6720
rect 8982 6511 9028 6557
rect 9140 6511 9186 6557
rect 8982 6348 9028 6394
rect 9140 6348 9186 6394
rect 8982 6184 9028 6230
rect 9140 6184 9186 6230
rect 8982 6021 9028 6067
rect 9140 6021 9186 6067
rect 8982 5858 9028 5904
rect 9140 5858 9186 5904
rect 8982 5695 9028 5741
rect 9140 5695 9186 5741
rect 3772 2673 3818 2719
rect 3896 2673 3942 2719
rect 4020 2673 4066 2719
rect 4144 2673 4190 2719
rect 4268 2673 4314 2719
rect 4392 2673 4438 2719
rect 4516 2673 4562 2719
rect 4640 2673 4686 2719
rect 4764 2673 4810 2719
rect 4888 2673 4934 2719
rect 5012 2673 5058 2719
rect 5136 2673 5182 2719
rect 5260 2673 5306 2719
rect 5384 2673 5430 2719
rect 5508 2673 5554 2719
rect 5632 2673 5678 2719
rect 5756 2673 5802 2719
rect 5880 2673 5926 2719
rect 6004 2673 6050 2719
rect 6128 2673 6174 2719
rect 6252 2673 6298 2719
rect 6376 2673 6422 2719
rect 6500 2673 6546 2719
rect 6624 2673 6670 2719
rect 6748 2673 6794 2719
rect 6872 2673 6918 2719
rect 6996 2673 7042 2719
rect 7120 2673 7166 2719
rect 7244 2673 7290 2719
rect 7368 2673 7414 2719
rect 3772 2549 3818 2595
rect 3896 2549 3942 2595
rect 4020 2549 4066 2595
rect 4144 2549 4190 2595
rect 4268 2549 4314 2595
rect 4392 2549 4438 2595
rect 4516 2549 4562 2595
rect 4640 2549 4686 2595
rect 4764 2549 4810 2595
rect 4888 2549 4934 2595
rect 5012 2549 5058 2595
rect 5136 2549 5182 2595
rect 5260 2549 5306 2595
rect 5384 2549 5430 2595
rect 5508 2549 5554 2595
rect 5632 2549 5678 2595
rect 5756 2549 5802 2595
rect 5880 2549 5926 2595
rect 6004 2549 6050 2595
rect 6128 2549 6174 2595
rect 6252 2549 6298 2595
rect 6376 2549 6422 2595
rect 6500 2549 6546 2595
rect 6624 2549 6670 2595
rect 6748 2549 6794 2595
rect 6872 2549 6918 2595
rect 6996 2549 7042 2595
rect 7120 2549 7166 2595
rect 7244 2549 7290 2595
rect 7368 2549 7414 2595
rect 3772 2425 3818 2471
rect 3896 2425 3942 2471
rect 4020 2425 4066 2471
rect 4144 2425 4190 2471
rect 4268 2425 4314 2471
rect 4392 2425 4438 2471
rect 4516 2425 4562 2471
rect 4640 2425 4686 2471
rect 4764 2425 4810 2471
rect 4888 2425 4934 2471
rect 5012 2425 5058 2471
rect 5136 2425 5182 2471
rect 5260 2425 5306 2471
rect 5384 2425 5430 2471
rect 5508 2425 5554 2471
rect 5632 2425 5678 2471
rect 5756 2425 5802 2471
rect 5880 2425 5926 2471
rect 6004 2425 6050 2471
rect 6128 2425 6174 2471
rect 6252 2425 6298 2471
rect 6376 2425 6422 2471
rect 6500 2425 6546 2471
rect 6624 2425 6670 2471
rect 6748 2425 6794 2471
rect 6872 2425 6918 2471
rect 6996 2425 7042 2471
rect 7120 2425 7166 2471
rect 7244 2425 7290 2471
rect 7368 2425 7414 2471
rect 3772 2301 3818 2347
rect 3896 2301 3942 2347
rect 4020 2301 4066 2347
rect 4144 2301 4190 2347
rect 4268 2301 4314 2347
rect 4392 2301 4438 2347
rect 4516 2301 4562 2347
rect 4640 2301 4686 2347
rect 4764 2301 4810 2347
rect 4888 2301 4934 2347
rect 5012 2301 5058 2347
rect 5136 2301 5182 2347
rect 5260 2301 5306 2347
rect 5384 2301 5430 2347
rect 5508 2301 5554 2347
rect 5632 2301 5678 2347
rect 5756 2301 5802 2347
rect 5880 2301 5926 2347
rect 6004 2301 6050 2347
rect 6128 2301 6174 2347
rect 6252 2301 6298 2347
rect 6376 2301 6422 2347
rect 6500 2301 6546 2347
rect 6624 2301 6670 2347
rect 6748 2301 6794 2347
rect 6872 2301 6918 2347
rect 6996 2301 7042 2347
rect 7120 2301 7166 2347
rect 7244 2301 7290 2347
rect 7368 2301 7414 2347
rect 13252 9123 13298 9169
rect 13410 9123 13456 9169
rect 13252 8960 13298 9006
rect 13410 8960 13456 9006
rect 13252 8797 13298 8843
rect 13410 8797 13456 8843
rect 13252 8633 13298 8679
rect 13410 8633 13456 8679
rect 13252 8470 13298 8516
rect 13410 8470 13456 8516
rect 13252 8307 13298 8353
rect 13410 8307 13456 8353
rect 13252 8144 13298 8190
rect 13410 8144 13456 8190
rect 13252 7980 13298 8026
rect 13410 7980 13456 8026
rect 13252 7817 13298 7863
rect 13410 7817 13456 7863
rect 13252 7654 13298 7700
rect 13410 7654 13456 7700
rect 13252 7491 13298 7537
rect 13410 7491 13456 7537
rect 13252 7327 13298 7373
rect 13410 7327 13456 7373
rect 13252 7164 13298 7210
rect 13410 7164 13456 7210
rect 13252 7001 13298 7047
rect 13410 7001 13456 7047
rect 13252 6837 13298 6883
rect 13410 6837 13456 6883
rect 13252 6674 13298 6720
rect 13410 6674 13456 6720
rect 13252 6511 13298 6557
rect 13410 6511 13456 6557
rect 13252 6348 13298 6394
rect 13410 6348 13456 6394
rect 13252 6184 13298 6230
rect 13410 6184 13456 6230
rect 13252 6021 13298 6067
rect 13410 6021 13456 6067
rect 13252 5858 13298 5904
rect 13410 5858 13456 5904
rect 13252 5695 13298 5741
rect 13410 5695 13456 5741
rect 13252 5531 13298 5577
rect 13410 5531 13456 5577
rect 13252 5368 13298 5414
rect 13410 5368 13456 5414
rect 13252 5205 13298 5251
rect 13410 5205 13456 5251
rect 13252 5042 13298 5088
rect 13410 5042 13456 5088
rect 13252 4879 13298 4925
rect 13410 4879 13456 4925
<< polysilicon >>
rect 6408 16001 6527 16028
rect 6632 16001 6751 16028
rect 6856 16001 6975 16028
rect 7080 16001 7199 16028
rect 7304 16001 7423 16028
rect 7528 16001 7647 16028
rect 7752 16001 7871 16028
rect 7976 16001 8095 16028
rect 8200 16001 8319 16028
rect 8424 16001 8543 16028
rect 6408 15957 6528 16001
rect 6632 15957 6752 16001
rect 6856 15957 6976 16001
rect 7080 15957 7200 16001
rect 7304 15957 7424 16001
rect 7528 15957 7648 16001
rect 7752 15957 7872 16001
rect 7976 15957 8096 16001
rect 8200 15957 8320 16001
rect 8424 15957 8544 16001
rect 8937 15957 9057 16001
rect 9161 15957 9281 16001
rect 9385 15957 9505 16001
rect 9609 15957 9729 16001
rect 9833 15957 9953 16001
rect 10057 15957 10177 16001
rect 10281 15957 10401 16001
rect 10505 15957 10625 16001
rect 10729 15957 10849 16001
rect 10953 15957 11073 16001
rect 11177 15957 11297 16001
rect 11401 15957 11521 16001
rect 11625 15957 11745 16001
rect 11849 15957 11969 16001
rect 12073 15957 12193 16001
rect 12297 15957 12417 16001
rect 12521 15957 12641 16001
rect 12745 15957 12865 16001
rect 12969 15957 13089 16001
rect 13193 15957 13313 16001
rect 6408 13401 6528 13461
rect 6632 13401 6752 13461
rect 6856 13401 6976 13461
rect 7080 13401 7200 13461
rect 7304 13401 7424 13461
rect 7528 13401 7648 13461
rect 7752 13401 7872 13461
rect 7976 13401 8096 13461
rect 8200 13401 8320 13461
rect 8424 13401 8544 13461
rect 6408 13382 8544 13401
rect 6408 13336 6474 13382
rect 8494 13336 8544 13382
rect 6408 13317 8544 13336
rect 8937 12223 9057 12283
rect 9161 12223 9281 12283
rect 9385 12223 9505 12283
rect 9609 12223 9729 12283
rect 9833 12223 9953 12283
rect 10057 12223 10177 12283
rect 10281 12223 10401 12283
rect 10505 12223 10625 12283
rect 10729 12223 10849 12283
rect 10953 12223 11073 12283
rect 11177 12223 11297 12283
rect 11401 12223 11521 12283
rect 11625 12223 11745 12283
rect 11849 12223 11969 12283
rect 12073 12223 12193 12283
rect 12297 12223 12417 12283
rect 12521 12223 12641 12283
rect 12745 12223 12865 12283
rect 12969 12223 13089 12283
rect 13193 12223 13313 12283
rect 8937 12204 13313 12223
rect 8937 12158 9003 12204
rect 13279 12158 13313 12204
rect 8937 12139 13313 12158
rect 8905 11438 13313 11457
rect 8905 11392 8924 11438
rect 13294 11392 13313 11438
rect 8905 11373 13313 11392
rect 8937 11313 9057 11373
rect 9161 11313 9281 11373
rect 9385 11313 9505 11373
rect 9609 11313 9729 11373
rect 9833 11313 9953 11373
rect 10057 11313 10177 11373
rect 10281 11313 10401 11373
rect 10505 11313 10625 11373
rect 10729 11313 10849 11373
rect 10953 11313 11073 11373
rect 11177 11313 11297 11373
rect 11401 11313 11521 11373
rect 11625 11313 11745 11373
rect 11849 11313 11969 11373
rect 12073 11313 12193 11373
rect 12297 11313 12417 11373
rect 12521 11313 12641 11373
rect 12745 11313 12865 11373
rect 12969 11313 13089 11373
rect 13193 11313 13313 11373
rect 6700 11160 7716 11179
rect 6700 11114 6766 11160
rect 7658 11114 7716 11160
rect 6700 11095 7716 11114
rect 6700 11035 6820 11095
rect 6924 11035 7044 11095
rect 7148 11035 7268 11095
rect 7372 11035 7492 11095
rect 7596 11035 7716 11095
rect 8937 9795 9057 9839
rect 9161 9795 9281 9839
rect 9385 9795 9505 9839
rect 9609 9795 9729 9839
rect 9833 9795 9953 9839
rect 10057 9795 10177 9839
rect 10281 9795 10401 9839
rect 10505 9795 10625 9839
rect 10729 9795 10849 9839
rect 10953 9795 11073 9839
rect 11177 9795 11297 9839
rect 11401 9795 11521 9839
rect 11625 9795 11745 9839
rect 11849 9795 11969 9839
rect 12073 9795 12193 9839
rect 12297 9795 12417 9839
rect 12521 9795 12641 9839
rect 12745 9795 12865 9839
rect 12969 9795 13089 9839
rect 13193 9795 13313 9839
rect 6700 8995 6820 9039
rect 6924 8995 7044 9039
rect 7148 8995 7268 9039
rect 7372 8995 7492 9039
rect 7596 8995 7716 9039
rect 6700 8965 6819 8995
rect 6924 8965 7043 8995
rect 7148 8965 7267 8995
rect 7372 8965 7491 8995
rect 7596 8965 7715 8995
rect 9526 9237 9645 9266
rect 9750 9237 9869 9266
rect 9974 9237 10093 9266
rect 9526 9193 9646 9237
rect 9750 9193 9870 9237
rect 9974 9193 10094 9237
rect 10725 9195 10845 9266
rect 10949 9195 11069 9266
rect 11173 9195 11293 9266
rect 11397 9195 11517 9266
rect 12010 9195 12130 9266
rect 12234 9195 12354 9266
rect 12458 9195 12578 9266
rect 12682 9195 12802 9266
rect 6972 8213 7092 8287
rect 7486 8213 7606 8287
rect 5055 8133 5175 8205
rect 5055 7867 5175 7941
rect 5055 7722 5174 7867
rect 6748 7742 6868 7816
rect 6972 7742 7092 8021
rect 7486 7961 7606 8021
rect 7755 7985 7947 8031
rect 7755 7961 7828 7985
rect 7486 7939 7828 7961
rect 7874 7939 7947 7985
rect 7486 7896 7947 7939
rect 7755 7821 7947 7896
rect 7486 7786 7605 7815
rect 7486 7742 7606 7786
rect 7755 7775 7828 7821
rect 7874 7775 7947 7821
rect 5055 7649 5175 7722
rect 7755 7729 7947 7775
rect 6748 7454 6868 7514
rect 6972 7454 7092 7514
rect 6166 7394 7092 7454
rect 7486 7477 7606 7550
rect 7486 7432 7723 7477
rect 6166 7393 6519 7394
rect 6166 7391 6518 7393
rect 6166 7345 6240 7391
rect 6286 7345 6398 7391
rect 6444 7345 6518 7391
rect 6166 7299 6518 7345
rect 7486 7386 7604 7432
rect 7650 7386 7723 7432
rect 7486 7340 7723 7386
rect 6748 7271 6868 7315
rect 6972 7271 7092 7315
rect 5055 7123 5175 7195
rect 5055 7078 5376 7123
rect 5055 7032 5256 7078
rect 5302 7032 5376 7078
rect 5055 6986 5376 7032
rect 5055 6587 5174 6659
rect 5279 6587 5398 6659
rect 7791 6978 7911 7729
rect 7486 6891 7911 6978
rect 7486 6831 7606 6891
rect 7486 6304 7606 6377
rect 5055 6069 5174 6131
rect 4981 6024 5174 6069
rect 4981 5978 5054 6024
rect 5100 5978 5174 6024
rect 4981 5932 5174 5978
rect 5055 5718 5174 5932
rect 5279 5857 5398 6131
rect 6748 6063 6868 6137
rect 6972 6063 7092 6137
rect 6748 6017 7254 6063
rect 6748 5971 7134 6017
rect 7180 5971 7254 6017
rect 7719 6033 7912 6078
rect 7719 6002 7793 6033
rect 6748 5925 7254 5971
rect 7486 5987 7793 6002
rect 7839 5987 7912 6033
rect 7486 5941 7912 5987
rect 5279 5811 5867 5857
rect 6748 5856 6868 5925
rect 6972 5856 7092 5925
rect 7486 5856 7606 5941
rect 5279 5765 5788 5811
rect 5834 5765 5867 5811
rect 5279 5734 5867 5765
rect 5055 5674 5175 5718
rect 5279 5674 5399 5734
rect 5055 5358 5175 5402
rect 5279 5358 5399 5402
rect 5055 5329 5174 5358
rect 5279 5329 5398 5358
rect 6748 5358 6868 5402
rect 6972 5358 7092 5402
rect 6748 5329 6867 5358
rect 6972 5329 7091 5358
rect 7486 5329 7606 5402
rect 9526 5095 9646 5293
rect 9526 4955 9568 5095
rect 9614 4955 9646 5095
rect 9526 4798 9646 4955
rect 9750 5095 9870 5293
rect 9750 4955 9791 5095
rect 9837 4955 9870 5095
rect 9750 4798 9870 4955
rect 9974 5095 10094 5293
rect 9974 4955 10015 5095
rect 10061 4955 10094 5095
rect 9974 4798 10094 4955
rect 8114 4437 8233 4467
rect 8114 4393 8234 4437
rect 5157 3892 5397 3936
rect 6235 3892 6475 3936
rect 6954 3897 7154 3941
rect 7600 3940 7720 3984
rect 5157 3603 5397 3772
rect 5157 3557 5623 3603
rect 6235 3602 6475 3772
rect 6954 3602 7154 3777
rect 7600 3602 7720 3790
rect 8114 3603 8234 3789
rect 8114 3602 8458 3603
rect 5157 3511 5345 3557
rect 5391 3511 5503 3557
rect 5549 3511 5623 3557
rect 5157 3465 5623 3511
rect 6109 3557 6475 3602
rect 6109 3511 6183 3557
rect 6229 3511 6475 3557
rect 6109 3465 6475 3511
rect 6833 3557 7154 3602
rect 6833 3511 6907 3557
rect 6953 3511 7154 3557
rect 6833 3465 7154 3511
rect 7473 3557 7720 3602
rect 7473 3511 7547 3557
rect 7593 3511 7720 3557
rect 7473 3465 7720 3511
rect 7991 3557 8458 3602
rect 7991 3511 8065 3557
rect 8111 3511 8458 3557
rect 7991 3465 8458 3511
rect 5157 3260 5397 3465
rect 6235 3260 6475 3465
rect 6954 3260 7154 3465
rect 7600 3260 7720 3465
rect 8114 3260 8234 3465
rect 8338 3260 8458 3465
rect 5157 3036 5397 3080
rect 6235 3036 6475 3080
rect 6954 3036 7154 3080
rect 7600 2838 7720 2882
rect 7600 2810 7719 2838
rect 8114 2462 8234 2506
rect 8338 2462 8458 2506
rect 8114 2434 8233 2462
rect 8338 2434 8457 2462
rect 10725 4537 10845 4659
rect 10725 4491 10763 4537
rect 10809 4491 10845 4537
rect 10725 4113 10845 4491
rect 10949 4338 11069 4659
rect 11173 4338 11293 4659
rect 10949 4319 11293 4338
rect 10949 4273 11049 4319
rect 11189 4273 11293 4319
rect 10949 4254 11293 4273
rect 10949 4113 11069 4254
rect 11173 4113 11293 4254
rect 11397 4537 11517 4659
rect 11397 4491 11434 4537
rect 11480 4491 11517 4537
rect 11397 4113 11517 4491
rect 12010 4288 12130 4659
rect 12234 4525 12354 4659
rect 12458 4525 12578 4659
rect 12010 4242 12046 4288
rect 12092 4242 12130 4288
rect 12010 4113 12130 4242
rect 12233 4506 12578 4525
rect 12233 4460 12294 4506
rect 12528 4460 12578 4506
rect 12233 4441 12578 4460
rect 12233 4113 12353 4441
rect 12458 4113 12578 4441
rect 12682 4307 12802 4659
rect 12681 4288 12802 4307
rect 12681 4242 12718 4288
rect 12764 4242 12802 4288
rect 12681 4223 12802 4242
rect 12681 4113 12801 4223
rect 12010 3132 12130 3205
rect 12233 3132 12353 3205
rect 12458 3132 12578 3205
rect 12681 3132 12801 3205
rect 10725 412 10845 484
rect 10949 412 11069 484
rect 11173 412 11293 484
rect 11397 412 11517 484
rect 9526 190 9646 262
rect 9750 190 9870 262
rect 9974 190 10094 262
<< polycontact >>
rect 6474 13336 8494 13382
rect 9003 12158 13279 12204
rect 8924 11392 13294 11438
rect 6766 11114 7658 11160
rect 7828 7939 7874 7985
rect 7828 7775 7874 7821
rect 6240 7345 6286 7391
rect 6398 7345 6444 7391
rect 7604 7386 7650 7432
rect 5256 7032 5302 7078
rect 5054 5978 5100 6024
rect 7134 5971 7180 6017
rect 7793 5987 7839 6033
rect 5788 5765 5834 5811
rect 9568 4955 9614 5095
rect 9791 4955 9837 5095
rect 10015 4955 10061 5095
rect 5345 3511 5391 3557
rect 5503 3511 5549 3557
rect 6183 3511 6229 3557
rect 6907 3511 6953 3557
rect 7547 3511 7593 3557
rect 8065 3511 8111 3557
rect 10763 4491 10809 4537
rect 11049 4273 11189 4319
rect 11434 4491 11480 4537
rect 12046 4242 12092 4288
rect 12294 4460 12528 4506
rect 12718 4242 12764 4288
<< metal1 >>
rect 6003 16273 13713 16310
rect 6003 16227 6192 16273
rect 6238 16238 6350 16273
rect 6238 16227 6329 16238
rect 6396 16227 6508 16273
rect 6554 16227 6666 16273
rect 6712 16238 6824 16273
rect 6712 16227 6777 16238
rect 6870 16227 6982 16273
rect 7028 16227 7140 16273
rect 7186 16238 7298 16273
rect 7186 16227 7225 16238
rect 6003 16186 6329 16227
rect 6381 16190 6777 16227
rect 6381 16186 6419 16190
rect 6003 16092 6419 16186
rect 6003 16046 6038 16092
rect 6084 16046 6419 16092
rect 6003 16020 6419 16046
rect 6003 15968 6329 16020
rect 6381 15968 6419 16020
rect 6003 15944 6419 15968
rect 6740 16186 6777 16190
rect 6829 16190 7225 16227
rect 6829 16186 6867 16190
rect 6740 16020 6867 16186
rect 6740 15968 6777 16020
rect 6829 15968 6867 16020
rect 6003 15928 6333 15944
rect 6003 15882 6038 15928
rect 6084 15882 6333 15928
rect 6003 15803 6333 15882
rect 6379 15803 6419 15944
rect 6003 15765 6329 15803
rect 6003 15719 6038 15765
rect 6084 15751 6329 15765
rect 6381 15751 6419 15803
rect 6084 15719 6333 15751
rect 6003 15602 6333 15719
rect 6003 15556 6038 15602
rect 6084 15585 6333 15602
rect 6379 15585 6419 15751
rect 6084 15556 6329 15585
rect 6003 15533 6329 15556
rect 6381 15533 6419 15585
rect 6003 15439 6333 15533
rect 6003 15393 6038 15439
rect 6084 15393 6333 15439
rect 6003 15367 6333 15393
rect 6379 15367 6419 15533
rect 6003 15315 6329 15367
rect 6381 15315 6419 15367
rect 6003 15275 6333 15315
rect 6003 15229 6038 15275
rect 6084 15229 6333 15275
rect 6003 15149 6333 15229
rect 6379 15149 6419 15315
rect 6003 15112 6329 15149
rect 6003 15066 6038 15112
rect 6084 15097 6329 15112
rect 6381 15097 6419 15149
rect 6084 15066 6333 15097
rect 6003 14949 6333 15066
rect 6003 14903 6038 14949
rect 6084 14932 6333 14949
rect 6379 14932 6419 15097
rect 6084 14903 6329 14932
rect 6003 14880 6329 14903
rect 6381 14880 6419 14932
rect 6003 14786 6333 14880
rect 6003 14740 6038 14786
rect 6084 14740 6333 14786
rect 6003 14714 6333 14740
rect 6379 14714 6419 14880
rect 6003 14662 6329 14714
rect 6381 14662 6419 14714
rect 6003 14622 6333 14662
rect 6003 14576 6038 14622
rect 6084 14576 6333 14622
rect 6003 14459 6333 14576
rect 6003 14413 6038 14459
rect 6084 14413 6333 14459
rect 6003 14296 6333 14413
rect 6003 14250 6038 14296
rect 6084 14250 6333 14296
rect 6003 14133 6333 14250
rect 6003 14087 6038 14133
rect 6084 14087 6333 14133
rect 6003 13970 6333 14087
rect 6003 13924 6038 13970
rect 6084 13924 6333 13970
rect 6003 13806 6333 13924
rect 6003 13760 6038 13806
rect 6084 13760 6333 13806
rect 6003 13643 6333 13760
rect 6003 13597 6038 13643
rect 6084 13597 6333 13643
rect 6003 13480 6333 13597
rect 6003 13434 6038 13480
rect 6084 13474 6333 13480
rect 6379 14622 6419 14662
rect 6557 15944 6603 15957
rect 6379 13474 6413 14622
rect 6084 13470 6413 13474
rect 6513 14433 6557 14474
rect 6740 15944 6867 15968
rect 7188 16186 7225 16190
rect 7277 16227 7298 16238
rect 7344 16227 7457 16273
rect 7503 16227 7615 16273
rect 7661 16238 7773 16273
rect 7661 16227 7673 16238
rect 7277 16190 7673 16227
rect 7277 16186 7315 16190
rect 7188 16020 7315 16186
rect 7188 15968 7225 16020
rect 7277 15968 7315 16020
rect 6740 15803 6781 15944
rect 6827 15803 6867 15944
rect 6740 15751 6777 15803
rect 6829 15751 6867 15803
rect 6740 15585 6781 15751
rect 6827 15585 6867 15751
rect 6740 15533 6777 15585
rect 6829 15533 6867 15585
rect 6740 15367 6781 15533
rect 6827 15367 6867 15533
rect 6740 15315 6777 15367
rect 6829 15315 6867 15367
rect 6740 15149 6781 15315
rect 6827 15149 6867 15315
rect 6740 15097 6777 15149
rect 6829 15097 6867 15149
rect 6740 14932 6781 15097
rect 6827 14932 6867 15097
rect 6740 14880 6777 14932
rect 6829 14880 6867 14932
rect 6740 14714 6781 14880
rect 6827 14714 6867 14880
rect 6740 14662 6777 14714
rect 6829 14662 6867 14714
rect 6740 14622 6781 14662
rect 6513 14381 6551 14433
rect 6513 14216 6557 14381
rect 6513 14164 6551 14216
rect 6513 13998 6557 14164
rect 6513 13946 6551 13998
rect 6513 13780 6557 13946
rect 6513 13728 6551 13780
rect 6513 13563 6557 13728
rect 6513 13511 6551 13563
rect 6513 13474 6557 13511
rect 6603 13474 6640 14474
rect 6513 13470 6640 13474
rect 6827 14622 6867 14662
rect 7005 15944 7051 15957
rect 6084 13434 6119 13470
rect 6333 13461 6379 13470
rect 6557 13461 6603 13470
rect 6781 13461 6827 13474
rect 6961 14433 7005 14474
rect 7188 15944 7315 15968
rect 7636 16186 7673 16190
rect 7725 16227 7773 16238
rect 7819 16227 7931 16273
rect 7977 16227 8089 16273
rect 8135 16238 8247 16273
rect 8173 16227 8247 16238
rect 8293 16227 8405 16273
rect 8451 16227 8563 16273
rect 8609 16238 8721 16273
rect 8621 16227 8721 16238
rect 8767 16238 8880 16273
rect 8767 16227 8859 16238
rect 8926 16227 9038 16273
rect 9084 16227 9196 16273
rect 9242 16238 9354 16273
rect 9242 16227 9307 16238
rect 9400 16227 9512 16273
rect 9558 16227 9670 16273
rect 9716 16238 9828 16273
rect 9716 16227 9755 16238
rect 7725 16190 8121 16227
rect 7725 16186 7763 16190
rect 7636 16020 7763 16186
rect 7636 15968 7673 16020
rect 7725 15968 7763 16020
rect 7188 15803 7229 15944
rect 7275 15803 7315 15944
rect 7188 15751 7225 15803
rect 7277 15751 7315 15803
rect 7188 15585 7229 15751
rect 7275 15585 7315 15751
rect 7188 15533 7225 15585
rect 7277 15533 7315 15585
rect 7188 15367 7229 15533
rect 7275 15367 7315 15533
rect 7188 15315 7225 15367
rect 7277 15315 7315 15367
rect 7188 15149 7229 15315
rect 7275 15149 7315 15315
rect 7188 15097 7225 15149
rect 7277 15097 7315 15149
rect 7188 14932 7229 15097
rect 7275 14932 7315 15097
rect 7188 14880 7225 14932
rect 7277 14880 7315 14932
rect 7188 14714 7229 14880
rect 7275 14714 7315 14880
rect 7188 14662 7225 14714
rect 7277 14662 7315 14714
rect 7188 14622 7229 14662
rect 6961 14381 6999 14433
rect 6961 14216 7005 14381
rect 6961 14164 6999 14216
rect 6961 13998 7005 14164
rect 6961 13946 6999 13998
rect 6961 13780 7005 13946
rect 6961 13728 6999 13780
rect 6961 13563 7005 13728
rect 6961 13511 6999 13563
rect 6961 13474 7005 13511
rect 7051 13474 7088 14474
rect 6961 13470 7088 13474
rect 7275 14622 7315 14662
rect 7453 15944 7499 15957
rect 7005 13461 7051 13470
rect 7229 13461 7275 13474
rect 7409 14433 7453 14474
rect 7636 15944 7763 15968
rect 8084 16186 8121 16190
rect 8173 16190 8569 16227
rect 8173 16186 8211 16190
rect 8084 16020 8211 16186
rect 8084 15968 8121 16020
rect 8173 15968 8211 16020
rect 7636 15803 7677 15944
rect 7723 15803 7763 15944
rect 7636 15751 7673 15803
rect 7725 15751 7763 15803
rect 7636 15585 7677 15751
rect 7723 15585 7763 15751
rect 7636 15533 7673 15585
rect 7725 15533 7763 15585
rect 7636 15367 7677 15533
rect 7723 15367 7763 15533
rect 7636 15315 7673 15367
rect 7725 15315 7763 15367
rect 7636 15149 7677 15315
rect 7723 15149 7763 15315
rect 7636 15097 7673 15149
rect 7725 15097 7763 15149
rect 7636 14932 7677 15097
rect 7723 14932 7763 15097
rect 7636 14880 7673 14932
rect 7725 14880 7763 14932
rect 7636 14714 7677 14880
rect 7723 14714 7763 14880
rect 7636 14662 7673 14714
rect 7725 14662 7763 14714
rect 7636 14622 7677 14662
rect 7409 14381 7447 14433
rect 7409 14216 7453 14381
rect 7409 14164 7447 14216
rect 7409 13998 7453 14164
rect 7409 13946 7447 13998
rect 7409 13780 7453 13946
rect 7409 13728 7447 13780
rect 7409 13563 7453 13728
rect 7409 13511 7447 13563
rect 7409 13474 7453 13511
rect 7499 13474 7536 14474
rect 7409 13470 7536 13474
rect 7723 14622 7763 14662
rect 7901 15944 7947 15957
rect 7453 13461 7499 13470
rect 7677 13461 7723 13474
rect 7857 14433 7901 14474
rect 8084 15944 8211 15968
rect 8532 16186 8569 16190
rect 8621 16190 8859 16227
rect 8621 16186 8659 16190
rect 8532 16020 8659 16186
rect 8532 15968 8569 16020
rect 8621 15968 8659 16020
rect 8084 15803 8125 15944
rect 8171 15803 8211 15944
rect 8084 15751 8121 15803
rect 8173 15751 8211 15803
rect 8084 15585 8125 15751
rect 8171 15585 8211 15751
rect 8084 15533 8121 15585
rect 8173 15533 8211 15585
rect 8084 15367 8125 15533
rect 8171 15367 8211 15533
rect 8084 15315 8121 15367
rect 8173 15315 8211 15367
rect 8084 15149 8125 15315
rect 8171 15149 8211 15315
rect 8084 15097 8121 15149
rect 8173 15097 8211 15149
rect 8084 14932 8125 15097
rect 8171 14932 8211 15097
rect 8084 14880 8121 14932
rect 8173 14880 8211 14932
rect 8084 14714 8125 14880
rect 8171 14714 8211 14880
rect 8084 14662 8121 14714
rect 8173 14662 8211 14714
rect 8084 14622 8125 14662
rect 7857 14381 7895 14433
rect 7857 14216 7901 14381
rect 7857 14164 7895 14216
rect 7857 13998 7901 14164
rect 7857 13946 7895 13998
rect 7857 13780 7901 13946
rect 7857 13728 7895 13780
rect 7857 13563 7901 13728
rect 7857 13511 7895 13563
rect 7857 13474 7901 13511
rect 7947 13474 7984 14474
rect 7857 13470 7984 13474
rect 8171 14622 8211 14662
rect 8349 15944 8395 15957
rect 7901 13461 7947 13470
rect 8125 13461 8171 13474
rect 8305 14433 8349 14474
rect 8532 15944 8659 15968
rect 8532 15803 8573 15944
rect 8619 15803 8659 15944
rect 8532 15751 8569 15803
rect 8621 15751 8659 15803
rect 8532 15585 8573 15751
rect 8619 15585 8659 15751
rect 8532 15533 8569 15585
rect 8621 15533 8659 15585
rect 8532 15367 8573 15533
rect 8619 15367 8659 15533
rect 8532 15315 8569 15367
rect 8621 15315 8659 15367
rect 8532 15149 8573 15315
rect 8619 15149 8659 15315
rect 8532 15097 8569 15149
rect 8621 15097 8659 15149
rect 8532 14932 8573 15097
rect 8619 14932 8659 15097
rect 8532 14880 8569 14932
rect 8621 14880 8659 14932
rect 8532 14714 8573 14880
rect 8619 14714 8659 14880
rect 8532 14662 8569 14714
rect 8621 14662 8659 14714
rect 8532 14622 8573 14662
rect 8305 14381 8343 14433
rect 8305 14216 8349 14381
rect 8305 14164 8343 14216
rect 8305 13998 8349 14164
rect 8305 13946 8343 13998
rect 8305 13780 8349 13946
rect 8305 13728 8343 13780
rect 8305 13563 8349 13728
rect 8305 13511 8343 13563
rect 8305 13474 8349 13511
rect 8395 13474 8432 14474
rect 8305 13470 8432 13474
rect 8619 14622 8659 14662
rect 8822 16186 8859 16190
rect 8911 16190 9307 16227
rect 8911 16186 8949 16190
rect 8822 16020 8949 16186
rect 8822 15968 8859 16020
rect 8911 15968 8949 16020
rect 8822 15944 8949 15968
rect 9270 16186 9307 16190
rect 9359 16190 9755 16227
rect 9359 16186 9397 16190
rect 9270 16020 9397 16186
rect 9270 15968 9307 16020
rect 9359 15968 9397 16020
rect 8822 15803 8862 15944
rect 8908 15803 8949 15944
rect 8822 15751 8859 15803
rect 8911 15751 8949 15803
rect 8822 15585 8862 15751
rect 8908 15585 8949 15751
rect 8822 15533 8859 15585
rect 8911 15533 8949 15585
rect 8822 15367 8862 15533
rect 8908 15367 8949 15533
rect 8822 15315 8859 15367
rect 8911 15315 8949 15367
rect 8822 15149 8862 15315
rect 8908 15149 8949 15315
rect 8822 15097 8859 15149
rect 8911 15097 8949 15149
rect 8822 14932 8862 15097
rect 8908 14932 8949 15097
rect 8822 14880 8859 14932
rect 8911 14880 8949 14932
rect 8822 14714 8862 14880
rect 8908 14714 8949 14880
rect 8822 14662 8859 14714
rect 8911 14662 8949 14714
rect 8822 14622 8862 14662
rect 8349 13461 8395 13470
rect 8573 13461 8619 13474
rect 6003 13317 6119 13434
rect 6463 13382 8505 13393
rect 6463 13336 6474 13382
rect 8494 13336 8505 13382
rect 6463 13325 6577 13336
rect 6003 13271 6038 13317
rect 6084 13271 6119 13317
rect 6003 13153 6119 13271
rect 6539 13284 6577 13325
rect 6629 13284 6788 13336
rect 6840 13284 7000 13336
rect 7052 13284 7211 13336
rect 7263 13325 8505 13336
rect 7263 13284 7301 13325
rect 6539 13243 7301 13284
rect 6003 13107 6038 13153
rect 6084 13141 6119 13153
rect 6084 13107 8645 13141
rect 6003 13104 8645 13107
rect 6003 13058 6349 13104
rect 6395 13058 6507 13104
rect 6553 13058 6665 13104
rect 6711 13058 6823 13104
rect 6869 13058 6982 13104
rect 7028 13058 7140 13104
rect 7186 13058 7298 13104
rect 7344 13058 7456 13104
rect 7502 13058 7614 13104
rect 7660 13058 7772 13104
rect 7818 13058 7930 13104
rect 7976 13058 8089 13104
rect 8135 13058 8247 13104
rect 8293 13058 8405 13104
rect 8451 13058 8563 13104
rect 8609 13058 8645 13104
rect 6003 12990 8645 13058
rect 6003 12944 6038 12990
rect 6084 12944 8645 12990
rect 6003 12941 8645 12944
rect 6003 12895 6349 12941
rect 6395 12895 6507 12941
rect 6553 12895 6665 12941
rect 6711 12895 6823 12941
rect 6869 12895 6982 12941
rect 7028 12895 7140 12941
rect 7186 12895 7298 12941
rect 7344 12895 7456 12941
rect 7502 12895 7614 12941
rect 7660 12895 7772 12941
rect 7818 12895 7930 12941
rect 7976 12895 8089 12941
rect 8135 12895 8247 12941
rect 8293 12895 8405 12941
rect 8451 12895 8563 12941
rect 8609 12895 8645 12941
rect 6003 12827 8645 12895
rect 6003 12781 6038 12827
rect 6084 12781 8645 12827
rect 6003 12777 8645 12781
rect 6003 12731 6349 12777
rect 6395 12731 6507 12777
rect 6553 12731 6665 12777
rect 6711 12731 6823 12777
rect 6869 12731 6982 12777
rect 7028 12731 7140 12777
rect 7186 12731 7298 12777
rect 7344 12731 7456 12777
rect 7502 12731 7614 12777
rect 7660 12731 7772 12777
rect 7818 12731 7930 12777
rect 7976 12731 8089 12777
rect 8135 12731 8247 12777
rect 8293 12731 8405 12777
rect 8451 12731 8563 12777
rect 8609 12731 8645 12777
rect 6003 12664 8645 12731
rect 6003 12618 6038 12664
rect 6084 12618 8645 12664
rect 6003 12614 8645 12618
rect 6003 12568 6349 12614
rect 6395 12568 6507 12614
rect 6553 12568 6665 12614
rect 6711 12568 6823 12614
rect 6869 12568 6982 12614
rect 7028 12568 7140 12614
rect 7186 12568 7298 12614
rect 7344 12568 7456 12614
rect 7502 12568 7614 12614
rect 7660 12568 7772 12614
rect 7818 12568 7930 12614
rect 7976 12568 8089 12614
rect 8135 12568 8247 12614
rect 8293 12568 8405 12614
rect 8451 12568 8563 12614
rect 8609 12568 8645 12614
rect 6003 12501 8645 12568
rect 6003 12455 6038 12501
rect 6084 12455 8645 12501
rect 6003 12451 8645 12455
rect 6003 12405 6349 12451
rect 6395 12405 6507 12451
rect 6553 12405 6665 12451
rect 6711 12405 6823 12451
rect 6869 12405 6982 12451
rect 7028 12405 7140 12451
rect 7186 12405 7298 12451
rect 7344 12405 7456 12451
rect 7502 12405 7614 12451
rect 7660 12405 7772 12451
rect 7818 12405 7930 12451
rect 7976 12405 8089 12451
rect 8135 12405 8247 12451
rect 8293 12405 8405 12451
rect 8451 12405 8563 12451
rect 8609 12405 8645 12451
rect 6003 12337 8645 12405
rect 6003 12291 6038 12337
rect 6084 12291 8645 12337
rect 6003 12287 8645 12291
rect 6003 12241 6349 12287
rect 6395 12241 6507 12287
rect 6553 12241 6665 12287
rect 6711 12241 6823 12287
rect 6869 12241 6982 12287
rect 7028 12241 7140 12287
rect 7186 12241 7298 12287
rect 7344 12241 7456 12287
rect 7502 12241 7614 12287
rect 7660 12241 7772 12287
rect 7818 12241 7930 12287
rect 7976 12241 8089 12287
rect 8135 12241 8247 12287
rect 8293 12241 8405 12287
rect 8451 12241 8563 12287
rect 8609 12241 8645 12287
rect 8908 14622 8949 14662
rect 9086 15944 9132 15957
rect 9045 14336 9086 14376
rect 9270 15944 9397 15968
rect 9718 16186 9755 16190
rect 9807 16227 9828 16238
rect 9874 16227 9986 16273
rect 10032 16227 10144 16273
rect 10190 16238 10303 16273
rect 10190 16227 10203 16238
rect 9807 16190 10203 16227
rect 9807 16186 9845 16190
rect 9718 16020 9845 16186
rect 9718 15968 9755 16020
rect 9807 15968 9845 16020
rect 9270 15803 9310 15944
rect 9356 15803 9397 15944
rect 9270 15751 9307 15803
rect 9359 15751 9397 15803
rect 9270 15585 9310 15751
rect 9356 15585 9397 15751
rect 9270 15533 9307 15585
rect 9359 15533 9397 15585
rect 9270 15367 9310 15533
rect 9356 15367 9397 15533
rect 9270 15315 9307 15367
rect 9359 15315 9397 15367
rect 9270 15149 9310 15315
rect 9356 15149 9397 15315
rect 9270 15097 9307 15149
rect 9359 15097 9397 15149
rect 9270 14932 9310 15097
rect 9356 14932 9397 15097
rect 9270 14880 9307 14932
rect 9359 14880 9397 14932
rect 9270 14714 9310 14880
rect 9356 14714 9397 14880
rect 9270 14662 9307 14714
rect 9359 14662 9397 14714
rect 9270 14622 9310 14662
rect 9132 14336 9174 14376
rect 9045 14284 9083 14336
rect 9135 14284 9174 14336
rect 9045 14118 9086 14284
rect 9132 14118 9174 14284
rect 9045 14066 9083 14118
rect 9135 14066 9174 14118
rect 9045 13900 9086 14066
rect 9132 13900 9174 14066
rect 9045 13848 9083 13900
rect 9135 13848 9174 13900
rect 9045 13683 9086 13848
rect 9132 13683 9174 13848
rect 9045 13631 9083 13683
rect 9135 13631 9174 13683
rect 9045 13465 9086 13631
rect 9132 13465 9174 13631
rect 9045 13413 9083 13465
rect 9135 13413 9174 13465
rect 9045 13247 9086 13413
rect 9132 13247 9174 13413
rect 9045 13195 9083 13247
rect 9135 13195 9174 13247
rect 9045 13030 9086 13195
rect 9132 13030 9174 13195
rect 9045 12978 9083 13030
rect 9135 12978 9174 13030
rect 9045 12812 9086 12978
rect 9132 12812 9174 12978
rect 9045 12760 9083 12812
rect 9135 12760 9174 12812
rect 9045 12594 9086 12760
rect 9132 12594 9174 12760
rect 9045 12542 9083 12594
rect 9135 12542 9174 12594
rect 9045 12502 9086 12542
rect 8862 12283 8908 12296
rect 9132 12502 9174 12542
rect 9086 12283 9132 12296
rect 9356 14622 9397 14662
rect 9534 15944 9580 15957
rect 9493 14336 9534 14376
rect 9718 15944 9845 15968
rect 10166 16186 10203 16190
rect 10255 16227 10303 16238
rect 10349 16227 10461 16273
rect 10507 16227 10619 16273
rect 10665 16238 10777 16273
rect 10703 16227 10777 16238
rect 10823 16227 10935 16273
rect 10981 16227 11093 16273
rect 11139 16238 11251 16273
rect 11151 16227 11251 16238
rect 11297 16227 11409 16273
rect 11455 16238 11567 16273
rect 11455 16227 11547 16238
rect 11613 16227 11726 16273
rect 11772 16227 11884 16273
rect 11930 16238 12042 16273
rect 11930 16227 11995 16238
rect 12088 16227 12200 16273
rect 12246 16227 12358 16273
rect 12404 16238 12516 16273
rect 12404 16227 12443 16238
rect 10255 16190 10651 16227
rect 10255 16186 10293 16190
rect 10166 16020 10293 16186
rect 10166 15968 10203 16020
rect 10255 15968 10293 16020
rect 9718 15803 9758 15944
rect 9804 15803 9845 15944
rect 9718 15751 9755 15803
rect 9807 15751 9845 15803
rect 9718 15585 9758 15751
rect 9804 15585 9845 15751
rect 9718 15533 9755 15585
rect 9807 15533 9845 15585
rect 9718 15367 9758 15533
rect 9804 15367 9845 15533
rect 9718 15315 9755 15367
rect 9807 15315 9845 15367
rect 9718 15149 9758 15315
rect 9804 15149 9845 15315
rect 9718 15097 9755 15149
rect 9807 15097 9845 15149
rect 9718 14932 9758 15097
rect 9804 14932 9845 15097
rect 9718 14880 9755 14932
rect 9807 14880 9845 14932
rect 9718 14714 9758 14880
rect 9804 14714 9845 14880
rect 9718 14662 9755 14714
rect 9807 14662 9845 14714
rect 9718 14622 9758 14662
rect 9580 14336 9622 14376
rect 9493 14284 9531 14336
rect 9583 14284 9622 14336
rect 9493 14118 9534 14284
rect 9580 14118 9622 14284
rect 9493 14066 9531 14118
rect 9583 14066 9622 14118
rect 9493 13900 9534 14066
rect 9580 13900 9622 14066
rect 9493 13848 9531 13900
rect 9583 13848 9622 13900
rect 9493 13683 9534 13848
rect 9580 13683 9622 13848
rect 9493 13631 9531 13683
rect 9583 13631 9622 13683
rect 9493 13465 9534 13631
rect 9580 13465 9622 13631
rect 9493 13413 9531 13465
rect 9583 13413 9622 13465
rect 9493 13247 9534 13413
rect 9580 13247 9622 13413
rect 9493 13195 9531 13247
rect 9583 13195 9622 13247
rect 9493 13030 9534 13195
rect 9580 13030 9622 13195
rect 9493 12978 9531 13030
rect 9583 12978 9622 13030
rect 9493 12812 9534 12978
rect 9580 12812 9622 12978
rect 9493 12760 9531 12812
rect 9583 12760 9622 12812
rect 9493 12594 9534 12760
rect 9580 12594 9622 12760
rect 9493 12542 9531 12594
rect 9583 12542 9622 12594
rect 9493 12502 9534 12542
rect 9310 12283 9356 12296
rect 9580 12502 9622 12542
rect 9534 12283 9580 12296
rect 9804 14622 9845 14662
rect 9982 15944 10028 15957
rect 9941 14336 9982 14376
rect 10166 15944 10293 15968
rect 10614 16186 10651 16190
rect 10703 16190 11099 16227
rect 10703 16186 10741 16190
rect 10614 16020 10741 16186
rect 10614 15968 10651 16020
rect 10703 15968 10741 16020
rect 10166 15803 10206 15944
rect 10252 15803 10293 15944
rect 10166 15751 10203 15803
rect 10255 15751 10293 15803
rect 10166 15585 10206 15751
rect 10252 15585 10293 15751
rect 10166 15533 10203 15585
rect 10255 15533 10293 15585
rect 10166 15367 10206 15533
rect 10252 15367 10293 15533
rect 10166 15315 10203 15367
rect 10255 15315 10293 15367
rect 10166 15149 10206 15315
rect 10252 15149 10293 15315
rect 10166 15097 10203 15149
rect 10255 15097 10293 15149
rect 10166 14932 10206 15097
rect 10252 14932 10293 15097
rect 10166 14880 10203 14932
rect 10255 14880 10293 14932
rect 10166 14714 10206 14880
rect 10252 14714 10293 14880
rect 10166 14662 10203 14714
rect 10255 14662 10293 14714
rect 10166 14622 10206 14662
rect 10028 14336 10070 14376
rect 9941 14284 9979 14336
rect 10031 14284 10070 14336
rect 9941 14118 9982 14284
rect 10028 14118 10070 14284
rect 9941 14066 9979 14118
rect 10031 14066 10070 14118
rect 9941 13900 9982 14066
rect 10028 13900 10070 14066
rect 9941 13848 9979 13900
rect 10031 13848 10070 13900
rect 9941 13683 9982 13848
rect 10028 13683 10070 13848
rect 9941 13631 9979 13683
rect 10031 13631 10070 13683
rect 9941 13465 9982 13631
rect 10028 13465 10070 13631
rect 9941 13413 9979 13465
rect 10031 13413 10070 13465
rect 9941 13247 9982 13413
rect 10028 13247 10070 13413
rect 9941 13195 9979 13247
rect 10031 13195 10070 13247
rect 9941 13030 9982 13195
rect 10028 13030 10070 13195
rect 9941 12978 9979 13030
rect 10031 12978 10070 13030
rect 9941 12812 9982 12978
rect 10028 12812 10070 12978
rect 9941 12760 9979 12812
rect 10031 12760 10070 12812
rect 9941 12594 9982 12760
rect 10028 12594 10070 12760
rect 9941 12542 9979 12594
rect 10031 12542 10070 12594
rect 9941 12502 9982 12542
rect 9758 12283 9804 12296
rect 10028 12502 10070 12542
rect 9982 12283 10028 12296
rect 10252 14622 10293 14662
rect 10430 15944 10476 15957
rect 10389 14336 10430 14376
rect 10614 15944 10741 15968
rect 11062 16186 11099 16190
rect 11151 16190 11547 16227
rect 11151 16186 11189 16190
rect 11062 16020 11189 16186
rect 11062 15968 11099 16020
rect 11151 15968 11189 16020
rect 10614 15803 10654 15944
rect 10700 15803 10741 15944
rect 10614 15751 10651 15803
rect 10703 15751 10741 15803
rect 10614 15585 10654 15751
rect 10700 15585 10741 15751
rect 10614 15533 10651 15585
rect 10703 15533 10741 15585
rect 10614 15367 10654 15533
rect 10700 15367 10741 15533
rect 10614 15315 10651 15367
rect 10703 15315 10741 15367
rect 10614 15149 10654 15315
rect 10700 15149 10741 15315
rect 10614 15097 10651 15149
rect 10703 15097 10741 15149
rect 10614 14932 10654 15097
rect 10700 14932 10741 15097
rect 10614 14880 10651 14932
rect 10703 14880 10741 14932
rect 10614 14714 10654 14880
rect 10700 14714 10741 14880
rect 10614 14662 10651 14714
rect 10703 14662 10741 14714
rect 10614 14622 10654 14662
rect 10476 14336 10518 14376
rect 10389 14284 10427 14336
rect 10479 14284 10518 14336
rect 10389 14118 10430 14284
rect 10476 14118 10518 14284
rect 10389 14066 10427 14118
rect 10479 14066 10518 14118
rect 10389 13900 10430 14066
rect 10476 13900 10518 14066
rect 10389 13848 10427 13900
rect 10479 13848 10518 13900
rect 10389 13683 10430 13848
rect 10476 13683 10518 13848
rect 10389 13631 10427 13683
rect 10479 13631 10518 13683
rect 10389 13465 10430 13631
rect 10476 13465 10518 13631
rect 10389 13413 10427 13465
rect 10479 13413 10518 13465
rect 10389 13247 10430 13413
rect 10476 13247 10518 13413
rect 10389 13195 10427 13247
rect 10479 13195 10518 13247
rect 10389 13030 10430 13195
rect 10476 13030 10518 13195
rect 10389 12978 10427 13030
rect 10479 12978 10518 13030
rect 10389 12812 10430 12978
rect 10476 12812 10518 12978
rect 10389 12760 10427 12812
rect 10479 12760 10518 12812
rect 10389 12594 10430 12760
rect 10476 12594 10518 12760
rect 10389 12542 10427 12594
rect 10479 12542 10518 12594
rect 10389 12502 10430 12542
rect 10206 12283 10252 12296
rect 10476 12502 10518 12542
rect 10430 12283 10476 12296
rect 10700 14622 10741 14662
rect 10878 15944 10924 15957
rect 10837 14336 10878 14376
rect 11062 15944 11189 15968
rect 11510 16186 11547 16190
rect 11599 16190 11995 16227
rect 11599 16186 11637 16190
rect 11510 16020 11637 16186
rect 11510 15968 11547 16020
rect 11599 15968 11637 16020
rect 11062 15803 11102 15944
rect 11148 15803 11189 15944
rect 11062 15751 11099 15803
rect 11151 15751 11189 15803
rect 11062 15585 11102 15751
rect 11148 15585 11189 15751
rect 11062 15533 11099 15585
rect 11151 15533 11189 15585
rect 11062 15367 11102 15533
rect 11148 15367 11189 15533
rect 11062 15315 11099 15367
rect 11151 15315 11189 15367
rect 11062 15149 11102 15315
rect 11148 15149 11189 15315
rect 11062 15097 11099 15149
rect 11151 15097 11189 15149
rect 11062 14932 11102 15097
rect 11148 14932 11189 15097
rect 11062 14880 11099 14932
rect 11151 14880 11189 14932
rect 11062 14714 11102 14880
rect 11148 14714 11189 14880
rect 11062 14662 11099 14714
rect 11151 14662 11189 14714
rect 11062 14622 11102 14662
rect 10924 14336 10966 14376
rect 10837 14284 10875 14336
rect 10927 14284 10966 14336
rect 10837 14118 10878 14284
rect 10924 14118 10966 14284
rect 10837 14066 10875 14118
rect 10927 14066 10966 14118
rect 10837 13900 10878 14066
rect 10924 13900 10966 14066
rect 10837 13848 10875 13900
rect 10927 13848 10966 13900
rect 10837 13683 10878 13848
rect 10924 13683 10966 13848
rect 10837 13631 10875 13683
rect 10927 13631 10966 13683
rect 10837 13465 10878 13631
rect 10924 13465 10966 13631
rect 10837 13413 10875 13465
rect 10927 13413 10966 13465
rect 10837 13247 10878 13413
rect 10924 13247 10966 13413
rect 10837 13195 10875 13247
rect 10927 13195 10966 13247
rect 10837 13030 10878 13195
rect 10924 13030 10966 13195
rect 10837 12978 10875 13030
rect 10927 12978 10966 13030
rect 10837 12812 10878 12978
rect 10924 12812 10966 12978
rect 10837 12760 10875 12812
rect 10927 12760 10966 12812
rect 10837 12594 10878 12760
rect 10924 12594 10966 12760
rect 10837 12542 10875 12594
rect 10927 12542 10966 12594
rect 10837 12502 10878 12542
rect 10654 12283 10700 12296
rect 10924 12502 10966 12542
rect 10878 12283 10924 12296
rect 11148 14622 11189 14662
rect 11326 15944 11372 15957
rect 11285 14336 11326 14376
rect 11510 15944 11637 15968
rect 11958 16186 11995 16190
rect 12047 16190 12443 16227
rect 12047 16186 12085 16190
rect 11958 16020 12085 16186
rect 11958 15968 11995 16020
rect 12047 15968 12085 16020
rect 11510 15803 11550 15944
rect 11596 15803 11637 15944
rect 11510 15751 11547 15803
rect 11599 15751 11637 15803
rect 11510 15585 11550 15751
rect 11596 15585 11637 15751
rect 11510 15533 11547 15585
rect 11599 15533 11637 15585
rect 11510 15367 11550 15533
rect 11596 15367 11637 15533
rect 11510 15315 11547 15367
rect 11599 15315 11637 15367
rect 11510 15149 11550 15315
rect 11596 15149 11637 15315
rect 11510 15097 11547 15149
rect 11599 15097 11637 15149
rect 11510 14932 11550 15097
rect 11596 14932 11637 15097
rect 11510 14880 11547 14932
rect 11599 14880 11637 14932
rect 11510 14714 11550 14880
rect 11596 14714 11637 14880
rect 11510 14662 11547 14714
rect 11599 14662 11637 14714
rect 11510 14622 11550 14662
rect 11372 14336 11414 14376
rect 11285 14284 11323 14336
rect 11375 14284 11414 14336
rect 11285 14118 11326 14284
rect 11372 14118 11414 14284
rect 11285 14066 11323 14118
rect 11375 14066 11414 14118
rect 11285 13900 11326 14066
rect 11372 13900 11414 14066
rect 11285 13848 11323 13900
rect 11375 13848 11414 13900
rect 11285 13683 11326 13848
rect 11372 13683 11414 13848
rect 11285 13631 11323 13683
rect 11375 13631 11414 13683
rect 11285 13465 11326 13631
rect 11372 13465 11414 13631
rect 11285 13413 11323 13465
rect 11375 13413 11414 13465
rect 11285 13247 11326 13413
rect 11372 13247 11414 13413
rect 11285 13195 11323 13247
rect 11375 13195 11414 13247
rect 11285 13030 11326 13195
rect 11372 13030 11414 13195
rect 11285 12978 11323 13030
rect 11375 12978 11414 13030
rect 11285 12812 11326 12978
rect 11372 12812 11414 12978
rect 11285 12760 11323 12812
rect 11375 12760 11414 12812
rect 11285 12594 11326 12760
rect 11372 12594 11414 12760
rect 11285 12542 11323 12594
rect 11375 12542 11414 12594
rect 11285 12502 11326 12542
rect 11102 12283 11148 12296
rect 11372 12502 11414 12542
rect 11326 12283 11372 12296
rect 11596 14622 11637 14662
rect 11774 15944 11820 15957
rect 11733 14336 11774 14376
rect 11958 15944 12085 15968
rect 12406 16186 12443 16190
rect 12495 16227 12516 16238
rect 12562 16227 12674 16273
rect 12720 16227 12832 16273
rect 12878 16238 12990 16273
rect 12878 16227 12891 16238
rect 12495 16190 12891 16227
rect 12495 16186 12533 16190
rect 12406 16020 12533 16186
rect 12406 15968 12443 16020
rect 12495 15968 12533 16020
rect 11958 15803 11998 15944
rect 12044 15803 12085 15944
rect 11958 15751 11995 15803
rect 12047 15751 12085 15803
rect 11958 15585 11998 15751
rect 12044 15585 12085 15751
rect 11958 15533 11995 15585
rect 12047 15533 12085 15585
rect 11958 15367 11998 15533
rect 12044 15367 12085 15533
rect 11958 15315 11995 15367
rect 12047 15315 12085 15367
rect 11958 15149 11998 15315
rect 12044 15149 12085 15315
rect 11958 15097 11995 15149
rect 12047 15097 12085 15149
rect 11958 14932 11998 15097
rect 12044 14932 12085 15097
rect 11958 14880 11995 14932
rect 12047 14880 12085 14932
rect 11958 14714 11998 14880
rect 12044 14714 12085 14880
rect 11958 14662 11995 14714
rect 12047 14662 12085 14714
rect 11958 14622 11998 14662
rect 11820 14336 11862 14376
rect 11733 14284 11771 14336
rect 11823 14284 11862 14336
rect 11733 14118 11774 14284
rect 11820 14118 11862 14284
rect 11733 14066 11771 14118
rect 11823 14066 11862 14118
rect 11733 13900 11774 14066
rect 11820 13900 11862 14066
rect 11733 13848 11771 13900
rect 11823 13848 11862 13900
rect 11733 13683 11774 13848
rect 11820 13683 11862 13848
rect 11733 13631 11771 13683
rect 11823 13631 11862 13683
rect 11733 13465 11774 13631
rect 11820 13465 11862 13631
rect 11733 13413 11771 13465
rect 11823 13413 11862 13465
rect 11733 13247 11774 13413
rect 11820 13247 11862 13413
rect 11733 13195 11771 13247
rect 11823 13195 11862 13247
rect 11733 13030 11774 13195
rect 11820 13030 11862 13195
rect 11733 12978 11771 13030
rect 11823 12978 11862 13030
rect 11733 12812 11774 12978
rect 11820 12812 11862 12978
rect 11733 12760 11771 12812
rect 11823 12760 11862 12812
rect 11733 12594 11774 12760
rect 11820 12594 11862 12760
rect 11733 12542 11771 12594
rect 11823 12542 11862 12594
rect 11733 12502 11774 12542
rect 11550 12283 11596 12296
rect 11820 12502 11862 12542
rect 11774 12283 11820 12296
rect 12044 14622 12085 14662
rect 12222 15944 12268 15957
rect 12181 14336 12222 14376
rect 12406 15944 12533 15968
rect 12854 16186 12891 16190
rect 12943 16227 12990 16238
rect 13036 16227 13149 16273
rect 13195 16227 13307 16273
rect 13353 16238 13465 16273
rect 13391 16227 13465 16238
rect 13511 16227 13713 16273
rect 12943 16190 13339 16227
rect 12943 16186 12981 16190
rect 12854 16020 12981 16186
rect 12854 15968 12891 16020
rect 12943 15968 12981 16020
rect 12406 15803 12446 15944
rect 12492 15803 12533 15944
rect 12406 15751 12443 15803
rect 12495 15751 12533 15803
rect 12406 15585 12446 15751
rect 12492 15585 12533 15751
rect 12406 15533 12443 15585
rect 12495 15533 12533 15585
rect 12406 15367 12446 15533
rect 12492 15367 12533 15533
rect 12406 15315 12443 15367
rect 12495 15315 12533 15367
rect 12406 15149 12446 15315
rect 12492 15149 12533 15315
rect 12406 15097 12443 15149
rect 12495 15097 12533 15149
rect 12406 14932 12446 15097
rect 12492 14932 12533 15097
rect 12406 14880 12443 14932
rect 12495 14880 12533 14932
rect 12406 14714 12446 14880
rect 12492 14714 12533 14880
rect 12406 14662 12443 14714
rect 12495 14662 12533 14714
rect 12406 14622 12446 14662
rect 12268 14336 12310 14376
rect 12181 14284 12219 14336
rect 12271 14284 12310 14336
rect 12181 14118 12222 14284
rect 12268 14118 12310 14284
rect 12181 14066 12219 14118
rect 12271 14066 12310 14118
rect 12181 13900 12222 14066
rect 12268 13900 12310 14066
rect 12181 13848 12219 13900
rect 12271 13848 12310 13900
rect 12181 13683 12222 13848
rect 12268 13683 12310 13848
rect 12181 13631 12219 13683
rect 12271 13631 12310 13683
rect 12181 13465 12222 13631
rect 12268 13465 12310 13631
rect 12181 13413 12219 13465
rect 12271 13413 12310 13465
rect 12181 13247 12222 13413
rect 12268 13247 12310 13413
rect 12181 13195 12219 13247
rect 12271 13195 12310 13247
rect 12181 13030 12222 13195
rect 12268 13030 12310 13195
rect 12181 12978 12219 13030
rect 12271 12978 12310 13030
rect 12181 12812 12222 12978
rect 12268 12812 12310 12978
rect 12181 12760 12219 12812
rect 12271 12760 12310 12812
rect 12181 12594 12222 12760
rect 12268 12594 12310 12760
rect 12181 12542 12219 12594
rect 12271 12542 12310 12594
rect 12181 12502 12222 12542
rect 11998 12283 12044 12296
rect 12268 12502 12310 12542
rect 12222 12283 12268 12296
rect 12492 14622 12533 14662
rect 12670 15944 12716 15957
rect 12629 14336 12670 14376
rect 12854 15944 12981 15968
rect 13301 16186 13339 16190
rect 13391 16186 13713 16227
rect 13301 16092 13713 16186
rect 13301 16046 13632 16092
rect 13678 16046 13713 16092
rect 13301 16020 13713 16046
rect 13301 15968 13339 16020
rect 13391 15968 13713 16020
rect 12854 15803 12894 15944
rect 12940 15803 12981 15944
rect 12854 15751 12891 15803
rect 12943 15751 12981 15803
rect 12854 15585 12894 15751
rect 12940 15585 12981 15751
rect 12854 15533 12891 15585
rect 12943 15533 12981 15585
rect 12854 15367 12894 15533
rect 12940 15367 12981 15533
rect 12854 15315 12891 15367
rect 12943 15315 12981 15367
rect 12854 15149 12894 15315
rect 12940 15149 12981 15315
rect 12854 15097 12891 15149
rect 12943 15097 12981 15149
rect 12854 14932 12894 15097
rect 12940 14932 12981 15097
rect 12854 14880 12891 14932
rect 12943 14880 12981 14932
rect 12854 14714 12894 14880
rect 12940 14714 12981 14880
rect 12854 14662 12891 14714
rect 12943 14662 12981 14714
rect 12854 14622 12894 14662
rect 12716 14336 12758 14376
rect 12629 14284 12667 14336
rect 12719 14284 12758 14336
rect 12629 14118 12670 14284
rect 12716 14118 12758 14284
rect 12629 14066 12667 14118
rect 12719 14066 12758 14118
rect 12629 13900 12670 14066
rect 12716 13900 12758 14066
rect 12629 13848 12667 13900
rect 12719 13848 12758 13900
rect 12629 13683 12670 13848
rect 12716 13683 12758 13848
rect 12629 13631 12667 13683
rect 12719 13631 12758 13683
rect 12629 13465 12670 13631
rect 12716 13465 12758 13631
rect 12629 13413 12667 13465
rect 12719 13413 12758 13465
rect 12629 13247 12670 13413
rect 12716 13247 12758 13413
rect 12629 13195 12667 13247
rect 12719 13195 12758 13247
rect 12629 13030 12670 13195
rect 12716 13030 12758 13195
rect 12629 12978 12667 13030
rect 12719 12978 12758 13030
rect 12629 12812 12670 12978
rect 12716 12812 12758 12978
rect 12629 12760 12667 12812
rect 12719 12760 12758 12812
rect 12629 12594 12670 12760
rect 12716 12594 12758 12760
rect 12629 12542 12667 12594
rect 12719 12542 12758 12594
rect 12629 12502 12670 12542
rect 12446 12283 12492 12296
rect 12716 12502 12758 12542
rect 12670 12283 12716 12296
rect 12940 14622 12981 14662
rect 13118 15944 13164 15957
rect 13077 14336 13118 14376
rect 13301 15944 13713 15968
rect 13301 15803 13342 15944
rect 13388 15928 13713 15944
rect 13388 15882 13632 15928
rect 13678 15882 13713 15928
rect 13388 15803 13713 15882
rect 13301 15751 13339 15803
rect 13391 15765 13713 15803
rect 13391 15751 13632 15765
rect 13301 15585 13342 15751
rect 13388 15719 13632 15751
rect 13678 15719 13713 15765
rect 13388 15602 13713 15719
rect 13388 15585 13632 15602
rect 13301 15533 13339 15585
rect 13391 15556 13632 15585
rect 13678 15556 13713 15602
rect 13391 15533 13713 15556
rect 13301 15367 13342 15533
rect 13388 15439 13713 15533
rect 13388 15393 13632 15439
rect 13678 15393 13713 15439
rect 13388 15367 13713 15393
rect 13301 15315 13339 15367
rect 13391 15315 13713 15367
rect 13301 15149 13342 15315
rect 13388 15275 13713 15315
rect 13388 15229 13632 15275
rect 13678 15229 13713 15275
rect 13388 15149 13713 15229
rect 13301 15097 13339 15149
rect 13391 15112 13713 15149
rect 13391 15097 13632 15112
rect 13301 14932 13342 15097
rect 13388 15066 13632 15097
rect 13678 15066 13713 15112
rect 13388 14949 13713 15066
rect 13388 14932 13632 14949
rect 13301 14880 13339 14932
rect 13391 14903 13632 14932
rect 13678 14903 13713 14949
rect 13391 14880 13713 14903
rect 13301 14714 13342 14880
rect 13388 14786 13713 14880
rect 13388 14740 13632 14786
rect 13678 14740 13713 14786
rect 13388 14714 13713 14740
rect 13301 14662 13339 14714
rect 13391 14662 13713 14714
rect 13164 14336 13206 14376
rect 13077 14284 13115 14336
rect 13167 14284 13206 14336
rect 13077 14118 13118 14284
rect 13164 14118 13206 14284
rect 13077 14066 13115 14118
rect 13167 14066 13206 14118
rect 13077 13900 13118 14066
rect 13164 13900 13206 14066
rect 13077 13848 13115 13900
rect 13167 13848 13206 13900
rect 13077 13683 13118 13848
rect 13164 13683 13206 13848
rect 13077 13631 13115 13683
rect 13167 13631 13206 13683
rect 13077 13465 13118 13631
rect 13164 13465 13206 13631
rect 13077 13413 13115 13465
rect 13167 13413 13206 13465
rect 13077 13247 13118 13413
rect 13164 13247 13206 13413
rect 13077 13195 13115 13247
rect 13167 13195 13206 13247
rect 13077 13030 13118 13195
rect 13164 13030 13206 13195
rect 13077 12978 13115 13030
rect 13167 12978 13206 13030
rect 13077 12812 13118 12978
rect 13164 12812 13206 12978
rect 13077 12760 13115 12812
rect 13167 12760 13206 12812
rect 13077 12594 13118 12760
rect 13164 12594 13206 12760
rect 13077 12542 13115 12594
rect 13167 12542 13206 12594
rect 13077 12502 13118 12542
rect 12894 12283 12940 12296
rect 13164 12502 13206 12542
rect 13118 12283 13164 12296
rect 13301 12296 13342 14662
rect 13388 14622 13713 14662
rect 13388 14576 13632 14622
rect 13678 14576 13713 14622
rect 13388 14459 13713 14576
rect 13388 14413 13632 14459
rect 13678 14413 13713 14459
rect 13388 14296 13713 14413
rect 13388 14250 13632 14296
rect 13678 14250 13713 14296
rect 13388 14133 13713 14250
rect 13388 14087 13632 14133
rect 13678 14087 13713 14133
rect 13388 13970 13713 14087
rect 13388 13924 13632 13970
rect 13678 13924 13713 13970
rect 13388 13806 13713 13924
rect 13388 13760 13632 13806
rect 13678 13760 13713 13806
rect 13388 13643 13713 13760
rect 13388 13597 13632 13643
rect 13678 13597 13713 13643
rect 13388 13480 13713 13597
rect 13388 13434 13632 13480
rect 13678 13434 13713 13480
rect 13388 13317 13713 13434
rect 13388 13271 13632 13317
rect 13678 13271 13713 13317
rect 13388 13153 13713 13271
rect 13388 13107 13632 13153
rect 13678 13107 13713 13153
rect 13388 12990 13713 13107
rect 13388 12944 13632 12990
rect 13678 12944 13713 12990
rect 13388 12827 13713 12944
rect 13388 12781 13632 12827
rect 13678 12781 13713 12827
rect 13388 12664 13713 12781
rect 13388 12618 13632 12664
rect 13678 12618 13713 12664
rect 13388 12501 13713 12618
rect 13388 12455 13632 12501
rect 13678 12455 13713 12501
rect 13388 12337 13713 12455
rect 13388 12296 13632 12337
rect 13301 12291 13632 12296
rect 13678 12291 13713 12337
rect 13342 12283 13388 12291
rect 6003 12174 8645 12241
rect 6003 12128 6038 12174
rect 6084 12128 8645 12174
rect 8992 12204 13290 12215
rect 8992 12158 9003 12204
rect 13279 12158 13290 12204
rect 8992 12147 9142 12158
rect 6003 12124 8645 12128
rect 6003 12078 6349 12124
rect 6395 12078 6507 12124
rect 6553 12078 6665 12124
rect 6711 12078 6823 12124
rect 6869 12078 6982 12124
rect 7028 12078 7140 12124
rect 7186 12078 7298 12124
rect 7344 12078 7456 12124
rect 7502 12078 7614 12124
rect 7660 12078 7772 12124
rect 7818 12078 7930 12124
rect 7976 12078 8089 12124
rect 8135 12078 8247 12124
rect 8293 12078 8405 12124
rect 8451 12078 8563 12124
rect 8609 12078 8645 12124
rect 9104 12118 9142 12147
rect 9194 12118 9353 12158
rect 9405 12118 9564 12158
rect 9616 12118 9774 12158
rect 9826 12118 9985 12158
rect 10037 12118 10197 12158
rect 10249 12118 10408 12158
rect 10460 12118 10618 12158
rect 10670 12118 10829 12158
rect 10881 12118 11040 12158
rect 11092 12147 13290 12158
rect 13597 12174 13713 12291
rect 11092 12118 11130 12147
rect 9104 12078 11130 12118
rect 13597 12128 13632 12174
rect 13678 12128 13713 12174
rect 6003 12011 8645 12078
rect 6003 11965 6038 12011
rect 6084 11998 8645 12011
rect 13597 12011 13713 12128
rect 13597 11998 13632 12011
rect 6084 11965 13632 11998
rect 13678 11965 13713 12011
rect 6003 11961 13713 11965
rect 6003 11915 6192 11961
rect 6238 11915 6350 11961
rect 6396 11915 6508 11961
rect 6554 11915 6666 11961
rect 6712 11915 6824 11961
rect 6870 11915 6982 11961
rect 7028 11915 7140 11961
rect 7186 11915 7298 11961
rect 7344 11915 7457 11961
rect 7503 11915 7615 11961
rect 7661 11915 7773 11961
rect 7819 11915 7931 11961
rect 7977 11915 8089 11961
rect 8135 11915 8247 11961
rect 8293 11915 8405 11961
rect 8451 11915 8563 11961
rect 8609 11915 8721 11961
rect 8767 11915 8880 11961
rect 8926 11915 9038 11961
rect 9084 11915 9196 11961
rect 9242 11915 9354 11961
rect 9400 11915 9512 11961
rect 9558 11915 9670 11961
rect 9716 11915 9828 11961
rect 9874 11915 9986 11961
rect 10032 11915 10144 11961
rect 10190 11915 10303 11961
rect 10349 11915 10461 11961
rect 10507 11915 10619 11961
rect 10665 11915 10777 11961
rect 10823 11915 10935 11961
rect 10981 11915 11093 11961
rect 11139 11915 11251 11961
rect 11297 11915 11409 11961
rect 11455 11915 11567 11961
rect 11613 11915 11726 11961
rect 11772 11915 11884 11961
rect 11930 11915 12042 11961
rect 12088 11915 12200 11961
rect 12246 11915 12358 11961
rect 12404 11915 12516 11961
rect 12562 11915 12674 11961
rect 12720 11915 12832 11961
rect 12878 11915 12990 11961
rect 13036 11915 13149 11961
rect 13195 11915 13307 11961
rect 13353 11915 13465 11961
rect 13511 11915 13713 11961
rect 6003 11878 13713 11915
rect 13608 11596 13724 11633
rect 13608 11550 13643 11596
rect 13689 11550 13724 11596
rect 6289 11478 8284 11515
rect 6289 11432 6323 11478
rect 6369 11432 6481 11478
rect 6527 11432 6639 11478
rect 6685 11432 6798 11478
rect 6844 11432 6956 11478
rect 7002 11432 7114 11478
rect 7160 11432 7272 11478
rect 7318 11432 7430 11478
rect 7476 11432 7588 11478
rect 7634 11432 7747 11478
rect 7793 11432 7905 11478
rect 7951 11432 8063 11478
rect 8109 11432 8284 11478
rect 9104 11477 11130 11517
rect 9104 11449 9142 11477
rect 6289 11395 8284 11432
rect 6289 11334 6404 11395
rect 6283 11333 6404 11334
rect 6276 11315 6404 11333
rect 6276 11293 6323 11315
rect 6276 11241 6314 11293
rect 6369 11269 6404 11315
rect 6366 11241 6404 11269
rect 6276 11152 6404 11241
rect 8010 11243 8284 11395
rect 8913 11438 9142 11449
rect 9194 11438 9353 11477
rect 9405 11438 9564 11477
rect 9616 11438 9774 11477
rect 9826 11438 9985 11477
rect 10037 11438 10197 11477
rect 10249 11438 10408 11477
rect 10460 11438 10618 11477
rect 10670 11438 10829 11477
rect 10881 11438 11040 11477
rect 11092 11449 11130 11477
rect 11092 11438 13305 11449
rect 8913 11392 8924 11438
rect 13294 11392 13305 11438
rect 8913 11381 13305 11392
rect 13608 11433 13724 11550
rect 13608 11387 13643 11433
rect 13689 11387 13724 11433
rect 6276 11106 6323 11152
rect 6369 11106 6404 11152
rect 6569 11200 7331 11240
rect 6569 11148 6607 11200
rect 6659 11160 6818 11200
rect 6870 11160 7030 11200
rect 7082 11160 7241 11200
rect 7293 11171 7331 11200
rect 8010 11197 8045 11243
rect 8091 11197 8203 11243
rect 8249 11197 8284 11243
rect 7293 11160 7669 11171
rect 6659 11148 6766 11160
rect 6569 11114 6766 11148
rect 7658 11114 7669 11160
rect 6569 11107 7669 11114
rect 6276 11075 6404 11106
rect 6755 11103 7669 11107
rect 6276 11023 6314 11075
rect 6366 11025 6404 11075
rect 8010 11080 8284 11197
rect 6625 11025 6671 11035
rect 6366 11023 6705 11025
rect 6276 11022 6705 11023
rect 6276 10988 6625 11022
rect 6276 10942 6323 10988
rect 6369 10942 6625 10988
rect 6276 10858 6625 10942
rect 6276 10806 6314 10858
rect 6366 10825 6625 10858
rect 6276 10779 6323 10806
rect 6369 10779 6625 10825
rect 6276 10662 6625 10779
rect 6276 10640 6323 10662
rect 6276 10588 6314 10640
rect 6369 10616 6625 10662
rect 6366 10588 6625 10616
rect 6276 10499 6625 10588
rect 6276 10453 6323 10499
rect 6369 10453 6625 10499
rect 6276 10422 6625 10453
rect 6276 10370 6314 10422
rect 6366 10370 6625 10422
rect 6276 10335 6625 10370
rect 6276 10289 6323 10335
rect 6369 10289 6625 10335
rect 6276 10205 6625 10289
rect 6276 10153 6314 10205
rect 6366 10172 6625 10205
rect 6276 10126 6323 10153
rect 6369 10126 6625 10172
rect 6276 10009 6625 10126
rect 6276 9987 6323 10009
rect 6276 9935 6314 9987
rect 6369 9963 6625 10009
rect 6366 9935 6625 9963
rect 6276 9895 6625 9935
rect 6289 9845 6625 9895
rect 6289 9799 6323 9845
rect 6369 9799 6625 9845
rect 6289 9682 6625 9799
rect 6289 9636 6323 9682
rect 6369 9636 6625 9682
rect 6289 9519 6625 9636
rect 6289 9473 6323 9519
rect 6369 9473 6625 9519
rect 6289 9356 6625 9473
rect 6289 9310 6323 9356
rect 6369 9310 6625 9356
rect 6289 9192 6625 9310
rect 6289 9146 6323 9192
rect 6369 9146 6625 9192
rect 6289 9052 6625 9146
rect 6671 9052 6705 11022
rect 6849 11022 6895 11035
rect 6815 10955 6849 10956
rect 6808 10915 6849 10955
rect 7073 11022 7119 11035
rect 6895 10955 6929 10956
rect 6895 10954 6933 10955
rect 6895 10915 6936 10954
rect 6808 10863 6846 10915
rect 6898 10863 6936 10915
rect 6808 10697 6849 10863
rect 6895 10697 6936 10863
rect 6808 10645 6846 10697
rect 6898 10645 6936 10697
rect 6808 10480 6849 10645
rect 6895 10480 6936 10645
rect 6808 10428 6846 10480
rect 6898 10428 6936 10480
rect 6808 10262 6849 10428
rect 6895 10262 6936 10428
rect 6808 10210 6846 10262
rect 6898 10210 6936 10262
rect 6808 10044 6849 10210
rect 6895 10044 6936 10210
rect 6808 9992 6846 10044
rect 6898 9992 6936 10044
rect 6808 9827 6849 9992
rect 6895 9827 6936 9992
rect 6808 9775 6846 9827
rect 6898 9775 6936 9827
rect 6808 9609 6849 9775
rect 6895 9609 6936 9775
rect 6808 9557 6846 9609
rect 6898 9557 6936 9609
rect 6808 9517 6849 9557
rect 6821 9516 6849 9517
rect 6289 9047 6705 9052
rect 6895 9516 6936 9557
rect 7032 10262 7073 10302
rect 7297 11022 7343 11035
rect 7262 10955 7297 10956
rect 7255 10915 7297 10955
rect 7521 11022 7567 11035
rect 7343 10955 7376 10956
rect 7343 10954 7380 10955
rect 7343 10915 7383 10954
rect 7255 10863 7293 10915
rect 7345 10863 7383 10915
rect 7255 10697 7297 10863
rect 7343 10697 7383 10863
rect 7255 10645 7293 10697
rect 7345 10645 7383 10697
rect 7255 10480 7297 10645
rect 7343 10480 7383 10645
rect 7255 10428 7293 10480
rect 7345 10428 7383 10480
rect 7119 10262 7160 10302
rect 7032 10210 7070 10262
rect 7122 10210 7160 10262
rect 7032 10044 7073 10210
rect 7119 10044 7160 10210
rect 7032 9992 7070 10044
rect 7122 9992 7160 10044
rect 7032 9826 7073 9992
rect 7119 9826 7160 9992
rect 7032 9774 7070 9826
rect 7122 9774 7160 9826
rect 7032 9608 7073 9774
rect 7119 9608 7160 9774
rect 7032 9556 7070 9608
rect 7122 9556 7160 9608
rect 7032 9516 7073 9556
rect 6289 9029 6404 9047
rect 6625 9039 6671 9047
rect 6849 9039 6895 9052
rect 7119 9516 7160 9556
rect 7255 10262 7297 10428
rect 7343 10262 7383 10428
rect 7255 10210 7293 10262
rect 7345 10210 7383 10262
rect 7255 10044 7297 10210
rect 7343 10044 7383 10210
rect 7255 9992 7293 10044
rect 7345 9992 7383 10044
rect 7255 9827 7297 9992
rect 7343 9827 7383 9992
rect 7255 9775 7293 9827
rect 7345 9775 7383 9827
rect 7255 9609 7297 9775
rect 7343 9609 7383 9775
rect 7255 9557 7293 9609
rect 7345 9557 7383 9609
rect 7255 9517 7297 9557
rect 7268 9516 7297 9517
rect 7073 9039 7119 9052
rect 7343 9516 7383 9557
rect 7479 10262 7521 10302
rect 7745 11022 7791 11035
rect 7710 10955 7745 10956
rect 7703 10915 7745 10955
rect 8010 11034 8045 11080
rect 8091 11034 8203 11080
rect 8249 11034 8284 11080
rect 7791 10955 7824 10956
rect 7791 10954 7828 10955
rect 7791 10915 7831 10954
rect 7703 10863 7741 10915
rect 7793 10863 7831 10915
rect 7703 10697 7745 10863
rect 7791 10697 7831 10863
rect 7703 10645 7741 10697
rect 7793 10645 7831 10697
rect 7703 10480 7745 10645
rect 7791 10480 7831 10645
rect 8010 10917 8284 11034
rect 8010 10871 8045 10917
rect 8091 10871 8203 10917
rect 8249 10871 8284 10917
rect 8010 10753 8284 10871
rect 8010 10707 8045 10753
rect 8091 10707 8203 10753
rect 8249 10707 8284 10753
rect 8010 10590 8284 10707
rect 8862 11300 8908 11313
rect 8010 10544 8045 10590
rect 8091 10544 8203 10590
rect 8249 10544 8284 10590
rect 8010 10515 8284 10544
rect 8823 10593 8862 10633
rect 9086 11300 9132 11313
rect 9045 11195 9086 11236
rect 9310 11300 9356 11313
rect 9132 11195 9173 11236
rect 9045 11143 9083 11195
rect 9135 11143 9173 11195
rect 9045 10978 9086 11143
rect 9132 10978 9173 11143
rect 9045 10926 9083 10978
rect 9135 10926 9173 10978
rect 9045 10760 9086 10926
rect 9132 10760 9173 10926
rect 9045 10708 9083 10760
rect 9135 10708 9173 10760
rect 8908 10593 8951 10633
rect 8823 10541 8861 10593
rect 8913 10541 8951 10593
rect 7703 10428 7741 10480
rect 7793 10428 7831 10480
rect 7567 10262 7607 10302
rect 7479 10210 7517 10262
rect 7569 10210 7607 10262
rect 7479 10044 7521 10210
rect 7567 10044 7607 10210
rect 7479 9992 7517 10044
rect 7569 9992 7607 10044
rect 7479 9826 7521 9992
rect 7567 9826 7607 9992
rect 7479 9774 7517 9826
rect 7569 9774 7607 9826
rect 7479 9608 7521 9774
rect 7567 9608 7607 9774
rect 7479 9556 7517 9608
rect 7569 9556 7607 9608
rect 7479 9516 7521 9556
rect 7297 9039 7343 9052
rect 7567 9516 7607 9556
rect 7703 10262 7745 10428
rect 7791 10262 7831 10428
rect 7703 10210 7741 10262
rect 7793 10210 7831 10262
rect 7703 10044 7745 10210
rect 7791 10044 7831 10210
rect 7703 9992 7741 10044
rect 7793 9992 7831 10044
rect 7703 9827 7745 9992
rect 7791 9827 7831 9992
rect 7703 9775 7741 9827
rect 7793 9775 7831 9827
rect 7703 9609 7745 9775
rect 7791 9609 7831 9775
rect 7703 9557 7741 9609
rect 7793 9557 7831 9609
rect 7703 9517 7745 9557
rect 7716 9516 7745 9517
rect 7521 9039 7567 9052
rect 7791 9516 7831 9557
rect 7980 10474 8319 10515
rect 7980 10422 8017 10474
rect 8069 10427 8229 10474
rect 7980 10381 8045 10422
rect 8091 10381 8203 10427
rect 8281 10422 8319 10474
rect 8249 10381 8319 10422
rect 7980 10264 8319 10381
rect 7980 10257 8045 10264
rect 7980 10205 8017 10257
rect 8091 10218 8203 10264
rect 8249 10257 8319 10264
rect 8069 10205 8229 10218
rect 8281 10205 8319 10257
rect 7980 10100 8319 10205
rect 7980 10054 8045 10100
rect 8091 10054 8203 10100
rect 8249 10054 8319 10100
rect 7980 10039 8319 10054
rect 7980 9987 8017 10039
rect 8069 9987 8229 10039
rect 8281 9987 8319 10039
rect 7980 9937 8319 9987
rect 7980 9891 8045 9937
rect 8091 9891 8203 9937
rect 8249 9891 8319 9937
rect 7980 9821 8319 9891
rect 8823 10375 8862 10541
rect 8908 10375 8951 10541
rect 8823 10323 8861 10375
rect 8913 10323 8951 10375
rect 8823 10157 8862 10323
rect 8908 10157 8951 10323
rect 8823 10105 8861 10157
rect 8913 10105 8951 10157
rect 8823 9939 8862 10105
rect 8908 9939 8951 10105
rect 9045 10542 9086 10708
rect 9132 10542 9173 10708
rect 9045 10490 9083 10542
rect 9135 10490 9173 10542
rect 9045 10324 9086 10490
rect 9132 10324 9173 10490
rect 9045 10272 9083 10324
rect 9135 10272 9173 10324
rect 9045 10107 9086 10272
rect 9132 10107 9173 10272
rect 9045 10055 9083 10107
rect 9135 10055 9173 10107
rect 9045 10015 9086 10055
rect 9051 10014 9086 10015
rect 8823 9887 8861 9939
rect 8913 9887 8951 9939
rect 8823 9852 8862 9887
rect 8908 9852 8951 9887
rect 8823 9847 8951 9852
rect 9132 10015 9173 10055
rect 9271 10593 9310 10633
rect 9534 11300 9580 11313
rect 9493 11195 9534 11236
rect 9758 11300 9804 11313
rect 9580 11195 9621 11236
rect 9493 11143 9531 11195
rect 9583 11143 9621 11195
rect 9493 10978 9534 11143
rect 9580 10978 9621 11143
rect 9493 10926 9531 10978
rect 9583 10926 9621 10978
rect 9493 10760 9534 10926
rect 9580 10760 9621 10926
rect 9493 10708 9531 10760
rect 9583 10708 9621 10760
rect 9356 10593 9399 10633
rect 9271 10541 9309 10593
rect 9361 10541 9399 10593
rect 9271 10375 9310 10541
rect 9356 10375 9399 10541
rect 9271 10323 9309 10375
rect 9361 10323 9399 10375
rect 9271 10157 9310 10323
rect 9356 10157 9399 10323
rect 9271 10105 9309 10157
rect 9361 10105 9399 10157
rect 9132 10014 9167 10015
rect 8862 9839 8908 9847
rect 9086 9839 9132 9852
rect 9271 9939 9310 10105
rect 9356 9939 9399 10105
rect 9493 10542 9534 10708
rect 9580 10542 9621 10708
rect 9493 10490 9531 10542
rect 9583 10490 9621 10542
rect 9493 10324 9534 10490
rect 9580 10324 9621 10490
rect 9493 10272 9531 10324
rect 9583 10272 9621 10324
rect 9493 10107 9534 10272
rect 9580 10107 9621 10272
rect 9493 10055 9531 10107
rect 9583 10055 9621 10107
rect 9493 10015 9534 10055
rect 9499 10014 9534 10015
rect 9271 9887 9309 9939
rect 9361 9887 9399 9939
rect 9271 9852 9310 9887
rect 9356 9852 9399 9887
rect 9271 9847 9399 9852
rect 9580 10015 9621 10055
rect 9719 10593 9758 10633
rect 9982 11300 10028 11313
rect 9941 11195 9982 11236
rect 10206 11300 10252 11313
rect 10028 11195 10069 11236
rect 9941 11143 9979 11195
rect 10031 11143 10069 11195
rect 9941 10978 9982 11143
rect 10028 10978 10069 11143
rect 9941 10926 9979 10978
rect 10031 10926 10069 10978
rect 9941 10760 9982 10926
rect 10028 10760 10069 10926
rect 9941 10708 9979 10760
rect 10031 10708 10069 10760
rect 9804 10593 9847 10633
rect 9719 10541 9757 10593
rect 9809 10541 9847 10593
rect 9719 10375 9758 10541
rect 9804 10375 9847 10541
rect 9719 10323 9757 10375
rect 9809 10323 9847 10375
rect 9719 10157 9758 10323
rect 9804 10157 9847 10323
rect 9719 10105 9757 10157
rect 9809 10105 9847 10157
rect 9580 10014 9615 10015
rect 9310 9839 9356 9847
rect 9534 9839 9580 9852
rect 9719 9939 9758 10105
rect 9804 9939 9847 10105
rect 9941 10542 9982 10708
rect 10028 10542 10069 10708
rect 9941 10490 9979 10542
rect 10031 10490 10069 10542
rect 9941 10324 9982 10490
rect 10028 10324 10069 10490
rect 9941 10272 9979 10324
rect 10031 10272 10069 10324
rect 9941 10107 9982 10272
rect 10028 10107 10069 10272
rect 9941 10055 9979 10107
rect 10031 10055 10069 10107
rect 9941 10015 9982 10055
rect 9947 10014 9982 10015
rect 9719 9887 9757 9939
rect 9809 9887 9847 9939
rect 9719 9852 9758 9887
rect 9804 9852 9847 9887
rect 9719 9847 9847 9852
rect 10028 10015 10069 10055
rect 10167 10593 10206 10633
rect 10430 11300 10476 11313
rect 10389 11195 10430 11236
rect 10654 11300 10700 11313
rect 10476 11195 10517 11236
rect 10389 11143 10427 11195
rect 10479 11143 10517 11195
rect 10389 10978 10430 11143
rect 10476 10978 10517 11143
rect 10389 10926 10427 10978
rect 10479 10926 10517 10978
rect 10389 10760 10430 10926
rect 10476 10760 10517 10926
rect 10389 10708 10427 10760
rect 10479 10708 10517 10760
rect 10252 10593 10295 10633
rect 10167 10541 10205 10593
rect 10257 10541 10295 10593
rect 10167 10375 10206 10541
rect 10252 10375 10295 10541
rect 10167 10323 10205 10375
rect 10257 10323 10295 10375
rect 10167 10157 10206 10323
rect 10252 10157 10295 10323
rect 10167 10105 10205 10157
rect 10257 10105 10295 10157
rect 10028 10014 10063 10015
rect 9758 9839 9804 9847
rect 9982 9839 10028 9852
rect 10167 9939 10206 10105
rect 10252 9939 10295 10105
rect 10389 10542 10430 10708
rect 10476 10542 10517 10708
rect 10389 10490 10427 10542
rect 10479 10490 10517 10542
rect 10389 10324 10430 10490
rect 10476 10324 10517 10490
rect 10389 10272 10427 10324
rect 10479 10272 10517 10324
rect 10389 10107 10430 10272
rect 10476 10107 10517 10272
rect 10389 10055 10427 10107
rect 10479 10055 10517 10107
rect 10389 10015 10430 10055
rect 10395 10014 10430 10015
rect 10167 9887 10205 9939
rect 10257 9887 10295 9939
rect 10167 9852 10206 9887
rect 10252 9852 10295 9887
rect 10167 9847 10295 9852
rect 10476 10015 10517 10055
rect 10615 10593 10654 10633
rect 10878 11300 10924 11313
rect 10837 11195 10878 11236
rect 11102 11300 11148 11313
rect 10924 11195 10965 11236
rect 10837 11143 10875 11195
rect 10927 11143 10965 11195
rect 10837 10978 10878 11143
rect 10924 10978 10965 11143
rect 10837 10926 10875 10978
rect 10927 10926 10965 10978
rect 10837 10760 10878 10926
rect 10924 10760 10965 10926
rect 10837 10708 10875 10760
rect 10927 10708 10965 10760
rect 10700 10593 10743 10633
rect 10615 10541 10653 10593
rect 10705 10541 10743 10593
rect 10615 10375 10654 10541
rect 10700 10375 10743 10541
rect 10615 10323 10653 10375
rect 10705 10323 10743 10375
rect 10615 10157 10654 10323
rect 10700 10157 10743 10323
rect 10615 10105 10653 10157
rect 10705 10105 10743 10157
rect 10476 10014 10511 10015
rect 10206 9839 10252 9847
rect 10430 9839 10476 9852
rect 10615 9939 10654 10105
rect 10700 9939 10743 10105
rect 10837 10542 10878 10708
rect 10924 10542 10965 10708
rect 10837 10490 10875 10542
rect 10927 10490 10965 10542
rect 10837 10324 10878 10490
rect 10924 10324 10965 10490
rect 10837 10272 10875 10324
rect 10927 10272 10965 10324
rect 10837 10107 10878 10272
rect 10924 10107 10965 10272
rect 10837 10055 10875 10107
rect 10927 10055 10965 10107
rect 10837 10015 10878 10055
rect 10843 10014 10878 10015
rect 10615 9887 10653 9939
rect 10705 9887 10743 9939
rect 10615 9852 10654 9887
rect 10700 9852 10743 9887
rect 10615 9847 10743 9852
rect 10924 10015 10965 10055
rect 11063 10593 11102 10633
rect 11326 11300 11372 11313
rect 11285 11195 11326 11236
rect 11550 11300 11596 11313
rect 11372 11195 11413 11236
rect 11285 11143 11323 11195
rect 11375 11143 11413 11195
rect 11285 10978 11326 11143
rect 11372 10978 11413 11143
rect 11285 10926 11323 10978
rect 11375 10926 11413 10978
rect 11285 10760 11326 10926
rect 11372 10760 11413 10926
rect 11285 10708 11323 10760
rect 11375 10708 11413 10760
rect 11148 10593 11191 10633
rect 11063 10541 11101 10593
rect 11153 10541 11191 10593
rect 11063 10375 11102 10541
rect 11148 10375 11191 10541
rect 11063 10323 11101 10375
rect 11153 10323 11191 10375
rect 11063 10157 11102 10323
rect 11148 10157 11191 10323
rect 11063 10105 11101 10157
rect 11153 10105 11191 10157
rect 10924 10014 10959 10015
rect 10654 9839 10700 9847
rect 10878 9839 10924 9852
rect 11063 9939 11102 10105
rect 11148 9939 11191 10105
rect 11285 10542 11326 10708
rect 11372 10542 11413 10708
rect 11285 10490 11323 10542
rect 11375 10490 11413 10542
rect 11285 10324 11326 10490
rect 11372 10324 11413 10490
rect 11285 10272 11323 10324
rect 11375 10272 11413 10324
rect 11285 10107 11326 10272
rect 11372 10107 11413 10272
rect 11285 10055 11323 10107
rect 11375 10055 11413 10107
rect 11285 10015 11326 10055
rect 11291 10014 11326 10015
rect 11063 9887 11101 9939
rect 11153 9887 11191 9939
rect 11063 9852 11102 9887
rect 11148 9852 11191 9887
rect 11063 9847 11191 9852
rect 11372 10015 11413 10055
rect 11511 10593 11550 10633
rect 11774 11300 11820 11313
rect 11733 11195 11774 11236
rect 11998 11300 12044 11313
rect 11820 11195 11861 11236
rect 11733 11143 11771 11195
rect 11823 11143 11861 11195
rect 11733 10978 11774 11143
rect 11820 10978 11861 11143
rect 11733 10926 11771 10978
rect 11823 10926 11861 10978
rect 11733 10760 11774 10926
rect 11820 10760 11861 10926
rect 11733 10708 11771 10760
rect 11823 10708 11861 10760
rect 11596 10593 11639 10633
rect 11511 10541 11549 10593
rect 11601 10541 11639 10593
rect 11511 10375 11550 10541
rect 11596 10375 11639 10541
rect 11511 10323 11549 10375
rect 11601 10323 11639 10375
rect 11511 10157 11550 10323
rect 11596 10157 11639 10323
rect 11511 10105 11549 10157
rect 11601 10105 11639 10157
rect 11372 10014 11407 10015
rect 11102 9839 11148 9847
rect 11326 9839 11372 9852
rect 11511 9939 11550 10105
rect 11596 9939 11639 10105
rect 11733 10542 11774 10708
rect 11820 10542 11861 10708
rect 11733 10490 11771 10542
rect 11823 10490 11861 10542
rect 11733 10324 11774 10490
rect 11820 10324 11861 10490
rect 11733 10272 11771 10324
rect 11823 10272 11861 10324
rect 11733 10107 11774 10272
rect 11820 10107 11861 10272
rect 11733 10055 11771 10107
rect 11823 10055 11861 10107
rect 11733 10015 11774 10055
rect 11739 10014 11774 10015
rect 11511 9887 11549 9939
rect 11601 9887 11639 9939
rect 11511 9852 11550 9887
rect 11596 9852 11639 9887
rect 11511 9847 11639 9852
rect 11820 10015 11861 10055
rect 11959 10593 11998 10633
rect 12222 11300 12268 11313
rect 12181 11195 12222 11236
rect 12446 11300 12492 11313
rect 12268 11195 12309 11236
rect 12181 11143 12219 11195
rect 12271 11143 12309 11195
rect 12181 10978 12222 11143
rect 12268 10978 12309 11143
rect 12181 10926 12219 10978
rect 12271 10926 12309 10978
rect 12181 10760 12222 10926
rect 12268 10760 12309 10926
rect 12181 10708 12219 10760
rect 12271 10708 12309 10760
rect 12044 10593 12087 10633
rect 11959 10541 11997 10593
rect 12049 10541 12087 10593
rect 11959 10375 11998 10541
rect 12044 10375 12087 10541
rect 11959 10323 11997 10375
rect 12049 10323 12087 10375
rect 11959 10157 11998 10323
rect 12044 10157 12087 10323
rect 11959 10105 11997 10157
rect 12049 10105 12087 10157
rect 11820 10014 11855 10015
rect 11550 9839 11596 9847
rect 11774 9839 11820 9852
rect 11959 9939 11998 10105
rect 12044 9939 12087 10105
rect 12181 10542 12222 10708
rect 12268 10542 12309 10708
rect 12181 10490 12219 10542
rect 12271 10490 12309 10542
rect 12181 10324 12222 10490
rect 12268 10324 12309 10490
rect 12181 10272 12219 10324
rect 12271 10272 12309 10324
rect 12181 10107 12222 10272
rect 12268 10107 12309 10272
rect 12181 10055 12219 10107
rect 12271 10055 12309 10107
rect 12181 10015 12222 10055
rect 12187 10014 12222 10015
rect 11959 9887 11997 9939
rect 12049 9887 12087 9939
rect 11959 9852 11998 9887
rect 12044 9852 12087 9887
rect 11959 9847 12087 9852
rect 12268 10015 12309 10055
rect 12407 10593 12446 10633
rect 12670 11300 12716 11313
rect 12629 11195 12670 11236
rect 12894 11300 12940 11313
rect 12716 11195 12757 11236
rect 12629 11143 12667 11195
rect 12719 11143 12757 11195
rect 12629 10978 12670 11143
rect 12716 10978 12757 11143
rect 12629 10926 12667 10978
rect 12719 10926 12757 10978
rect 12629 10760 12670 10926
rect 12716 10760 12757 10926
rect 12629 10708 12667 10760
rect 12719 10708 12757 10760
rect 12492 10593 12535 10633
rect 12407 10541 12445 10593
rect 12497 10541 12535 10593
rect 12407 10375 12446 10541
rect 12492 10375 12535 10541
rect 12407 10323 12445 10375
rect 12497 10323 12535 10375
rect 12407 10157 12446 10323
rect 12492 10157 12535 10323
rect 12407 10105 12445 10157
rect 12497 10105 12535 10157
rect 12268 10014 12303 10015
rect 11998 9839 12044 9847
rect 12222 9839 12268 9852
rect 12407 9939 12446 10105
rect 12492 9939 12535 10105
rect 12629 10542 12670 10708
rect 12716 10542 12757 10708
rect 12629 10490 12667 10542
rect 12719 10490 12757 10542
rect 12629 10324 12670 10490
rect 12716 10324 12757 10490
rect 12629 10272 12667 10324
rect 12719 10272 12757 10324
rect 12629 10107 12670 10272
rect 12716 10107 12757 10272
rect 12629 10055 12667 10107
rect 12719 10055 12757 10107
rect 12629 10015 12670 10055
rect 12635 10014 12670 10015
rect 12407 9887 12445 9939
rect 12497 9887 12535 9939
rect 12407 9852 12446 9887
rect 12492 9852 12535 9887
rect 12407 9847 12535 9852
rect 12716 10015 12757 10055
rect 12855 10593 12894 10633
rect 13118 11300 13164 11313
rect 13342 11304 13388 11313
rect 13608 11304 13724 11387
rect 13077 11195 13118 11236
rect 13301 11300 13724 11304
rect 13164 11195 13205 11236
rect 13077 11143 13115 11195
rect 13167 11143 13205 11195
rect 13077 10978 13118 11143
rect 13164 10978 13205 11143
rect 13077 10926 13115 10978
rect 13167 10926 13205 10978
rect 13077 10760 13118 10926
rect 13164 10760 13205 10926
rect 13077 10708 13115 10760
rect 13167 10708 13205 10760
rect 12940 10593 12983 10633
rect 12855 10541 12893 10593
rect 12945 10541 12983 10593
rect 12855 10375 12894 10541
rect 12940 10375 12983 10541
rect 12855 10323 12893 10375
rect 12945 10323 12983 10375
rect 12855 10157 12894 10323
rect 12940 10157 12983 10323
rect 12855 10105 12893 10157
rect 12945 10105 12983 10157
rect 12716 10014 12751 10015
rect 12446 9839 12492 9847
rect 12670 9839 12716 9852
rect 12855 9939 12894 10105
rect 12940 9939 12983 10105
rect 13077 10542 13118 10708
rect 13164 10542 13205 10708
rect 13077 10490 13115 10542
rect 13167 10490 13205 10542
rect 13077 10324 13118 10490
rect 13164 10324 13205 10490
rect 13077 10272 13115 10324
rect 13167 10272 13205 10324
rect 13077 10107 13118 10272
rect 13164 10107 13205 10272
rect 13077 10055 13115 10107
rect 13167 10055 13205 10107
rect 13077 10015 13118 10055
rect 13083 10014 13118 10015
rect 12855 9887 12893 9939
rect 12945 9887 12983 9939
rect 12855 9852 12894 9887
rect 12940 9852 12983 9887
rect 12855 9847 12983 9852
rect 13164 10015 13205 10055
rect 13301 10593 13342 11300
rect 13388 11270 13724 11300
rect 13388 11224 13643 11270
rect 13689 11224 13724 11270
rect 13388 11107 13724 11224
rect 13388 11061 13643 11107
rect 13689 11061 13724 11107
rect 13388 10943 13724 11061
rect 13388 10897 13643 10943
rect 13689 10897 13724 10943
rect 13388 10780 13724 10897
rect 13388 10734 13643 10780
rect 13689 10734 13724 10780
rect 13388 10667 13724 10734
rect 13388 10627 13730 10667
rect 13388 10593 13640 10627
rect 13301 10541 13339 10593
rect 13391 10575 13640 10593
rect 13692 10575 13730 10627
rect 13391 10571 13643 10575
rect 13689 10571 13730 10575
rect 13391 10541 13730 10571
rect 13301 10375 13342 10541
rect 13388 10453 13730 10541
rect 13388 10409 13643 10453
rect 13689 10409 13730 10453
rect 13388 10375 13640 10409
rect 13301 10323 13339 10375
rect 13391 10357 13640 10375
rect 13692 10357 13730 10409
rect 13391 10323 13730 10357
rect 13301 10157 13342 10323
rect 13388 10290 13730 10323
rect 13388 10244 13643 10290
rect 13689 10244 13730 10290
rect 13388 10191 13730 10244
rect 13388 10157 13640 10191
rect 13301 10105 13339 10157
rect 13391 10139 13640 10157
rect 13692 10139 13730 10191
rect 13391 10127 13730 10139
rect 13391 10105 13643 10127
rect 13164 10014 13199 10015
rect 12894 9839 12940 9847
rect 13118 9839 13164 9852
rect 13301 9939 13342 10105
rect 13388 10081 13643 10105
rect 13689 10081 13730 10127
rect 13388 9973 13730 10081
rect 13388 9939 13640 9973
rect 13301 9887 13339 9939
rect 13391 9921 13640 9939
rect 13692 9921 13730 9973
rect 13391 9918 13643 9921
rect 13689 9918 13730 9921
rect 13391 9887 13730 9918
rect 13301 9852 13342 9887
rect 13388 9881 13730 9887
rect 13388 9852 13724 9881
rect 13301 9847 13724 9852
rect 13342 9839 13388 9847
rect 7980 9769 8017 9821
rect 8069 9774 8229 9821
rect 7980 9728 8045 9769
rect 8091 9728 8203 9774
rect 8281 9769 8319 9821
rect 8249 9728 8319 9769
rect 7980 9610 8319 9728
rect 7980 9604 8045 9610
rect 7980 9552 8017 9604
rect 8091 9564 8203 9610
rect 8249 9604 8319 9610
rect 8069 9552 8229 9564
rect 8281 9552 8319 9604
rect 7980 9511 8319 9552
rect 7745 9039 7791 9052
rect 8010 9447 8284 9511
rect 8010 9401 8045 9447
rect 8091 9401 8203 9447
rect 8249 9401 8284 9447
rect 8010 9284 8284 9401
rect 8010 9238 8045 9284
rect 8091 9238 8203 9284
rect 8249 9238 8284 9284
rect 8010 9121 8284 9238
rect 8010 9075 8045 9121
rect 8091 9075 8203 9121
rect 8249 9075 8284 9121
rect 6289 8983 6323 9029
rect 6369 8983 6404 9029
rect 6289 8915 6404 8983
rect 8010 8957 8284 9075
rect 6289 8866 6405 8915
rect 6289 8820 6323 8866
rect 6369 8820 6405 8866
rect 6289 8668 6405 8820
rect 8010 8911 8045 8957
rect 8091 8911 8203 8957
rect 8249 8911 8284 8957
rect 8010 8794 8284 8911
rect 8010 8748 8045 8794
rect 8091 8748 8203 8794
rect 8249 8748 8284 8794
rect 8010 8668 8284 8748
rect 355 8631 8284 8668
rect 355 8585 400 8631
rect 446 8585 558 8631
rect 604 8585 716 8631
rect 762 8585 875 8631
rect 921 8585 1033 8631
rect 1079 8585 1191 8631
rect 1237 8585 1349 8631
rect 1395 8585 1507 8631
rect 1553 8585 1665 8631
rect 1711 8585 1823 8631
rect 1869 8585 1981 8631
rect 2027 8585 2139 8631
rect 2185 8585 2298 8631
rect 2344 8585 2456 8631
rect 2502 8585 2614 8631
rect 2660 8585 2772 8631
rect 2818 8585 2930 8631
rect 2976 8585 3088 8631
rect 3134 8585 3246 8631
rect 3292 8585 3404 8631
rect 3450 8585 3562 8631
rect 3608 8585 3721 8631
rect 3767 8585 3879 8631
rect 3925 8585 4037 8631
rect 4083 8585 4195 8631
rect 4241 8585 4353 8631
rect 4399 8585 4511 8631
rect 4557 8585 4670 8631
rect 4716 8585 4828 8631
rect 4874 8585 4986 8631
rect 5032 8585 5144 8631
rect 5190 8585 5302 8631
rect 5348 8585 5460 8631
rect 5506 8585 5618 8631
rect 5664 8585 5776 8631
rect 5822 8585 5934 8631
rect 5980 8585 6093 8631
rect 6139 8585 6251 8631
rect 6297 8585 6409 8631
rect 6455 8585 6567 8631
rect 6613 8585 6725 8631
rect 6771 8585 6883 8631
rect 6929 8585 7041 8631
rect 7087 8585 7199 8631
rect 7245 8585 7357 8631
rect 7403 8585 7516 8631
rect 7562 8585 7674 8631
rect 7720 8585 7832 8631
rect 7878 8585 8045 8631
rect 8091 8585 8203 8631
rect 8249 8585 8284 8631
rect 355 8548 8284 8585
rect 8947 9495 13491 9532
rect 8947 9449 8982 9495
rect 9028 9449 9140 9495
rect 9186 9449 9299 9495
rect 9345 9449 9457 9495
rect 9503 9449 9615 9495
rect 9661 9449 9773 9495
rect 9819 9449 9931 9495
rect 9977 9449 10089 9495
rect 10135 9449 10247 9495
rect 10293 9449 10405 9495
rect 10451 9449 10563 9495
rect 10609 9449 10722 9495
rect 10768 9449 10880 9495
rect 10926 9449 11038 9495
rect 11084 9449 11196 9495
rect 11242 9449 11354 9495
rect 11400 9449 11512 9495
rect 11558 9449 11671 9495
rect 11717 9449 11829 9495
rect 11875 9449 11987 9495
rect 12033 9449 12145 9495
rect 12191 9449 12303 9495
rect 12349 9449 12461 9495
rect 12507 9449 12619 9495
rect 12665 9449 12777 9495
rect 12823 9449 12935 9495
rect 12981 9449 13094 9495
rect 13140 9449 13252 9495
rect 13298 9449 13410 9495
rect 13456 9449 13491 9495
rect 8947 9412 13491 9449
rect 8947 9332 9532 9412
rect 8947 9286 8982 9332
rect 9028 9286 9140 9332
rect 9186 9286 9532 9332
rect 8947 9180 9532 9286
rect 8947 9169 9451 9180
rect 8947 9123 8982 9169
rect 9028 9123 9140 9169
rect 9186 9123 9451 9169
rect 8947 9006 9451 9123
rect 8947 8960 8982 9006
rect 9028 8960 9140 9006
rect 9186 8960 9451 9006
rect 8947 8842 9451 8960
rect 8947 8796 8982 8842
rect 9028 8796 9140 8842
rect 9186 8796 9451 8842
rect 8947 8679 9451 8796
rect 8947 8633 8982 8679
rect 9028 8633 9140 8679
rect 9186 8633 9451 8679
rect 355 8306 4292 8548
rect 4944 8543 5061 8548
rect 355 8260 403 8306
rect 449 8260 561 8306
rect 607 8260 719 8306
rect 765 8260 877 8306
rect 923 8260 1035 8306
rect 1081 8260 1193 8306
rect 1239 8260 1351 8306
rect 1397 8260 1509 8306
rect 1555 8260 1667 8306
rect 1713 8260 1826 8306
rect 1872 8260 1984 8306
rect 2030 8260 2142 8306
rect 2188 8260 2300 8306
rect 2346 8260 2458 8306
rect 2504 8260 2616 8306
rect 2662 8260 2774 8306
rect 2820 8260 2933 8306
rect 2979 8260 3091 8306
rect 3137 8260 3249 8306
rect 3295 8260 3407 8306
rect 3453 8260 3565 8306
rect 3611 8260 3723 8306
rect 3769 8260 3881 8306
rect 3927 8260 4039 8306
rect 4085 8260 4197 8306
rect 4243 8260 4292 8306
rect 355 8258 4292 8260
rect 355 8206 457 8258
rect 509 8206 668 8258
rect 720 8206 878 8258
rect 930 8206 1089 8258
rect 1141 8206 1300 8258
rect 1352 8206 1511 8258
rect 1563 8206 1722 8258
rect 1774 8206 1932 8258
rect 1984 8206 2143 8258
rect 2195 8206 2355 8258
rect 2407 8206 2566 8258
rect 2618 8206 2776 8258
rect 2828 8206 2987 8258
rect 3039 8206 3198 8258
rect 3250 8206 3409 8258
rect 3461 8206 3620 8258
rect 3672 8206 3830 8258
rect 3882 8206 4041 8258
rect 4093 8206 4292 8258
rect 355 8143 4292 8206
rect 355 8097 403 8143
rect 449 8097 561 8143
rect 607 8097 719 8143
rect 765 8097 877 8143
rect 923 8097 1035 8143
rect 1081 8097 1193 8143
rect 1239 8097 1351 8143
rect 1397 8097 1509 8143
rect 1555 8097 1667 8143
rect 1713 8097 1826 8143
rect 1872 8097 1984 8143
rect 2030 8097 2142 8143
rect 2188 8097 2300 8143
rect 2346 8097 2458 8143
rect 2504 8097 2616 8143
rect 2662 8097 2774 8143
rect 2820 8097 2933 8143
rect 2979 8097 3091 8143
rect 3137 8097 3249 8143
rect 3295 8097 3407 8143
rect 3453 8097 3565 8143
rect 3611 8097 3723 8143
rect 3769 8097 3881 8143
rect 3927 8097 4039 8143
rect 4085 8097 4197 8143
rect 4243 8097 4292 8143
rect 355 8040 4292 8097
rect 355 7988 457 8040
rect 509 7988 668 8040
rect 720 7988 878 8040
rect 930 7988 1089 8040
rect 1141 7988 1300 8040
rect 1352 7988 1511 8040
rect 1563 7988 1722 8040
rect 1774 7988 1932 8040
rect 1984 7988 2143 8040
rect 2195 7988 2355 8040
rect 2407 7988 2566 8040
rect 2618 7988 2776 8040
rect 2828 7988 2987 8040
rect 3039 7988 3198 8040
rect 3250 7988 3409 8040
rect 3461 7988 3620 8040
rect 3672 7988 3830 8040
rect 3882 7988 4041 8040
rect 4093 7988 4292 8040
rect 355 7980 4292 7988
rect 355 7934 403 7980
rect 449 7934 561 7980
rect 607 7934 719 7980
rect 765 7934 877 7980
rect 923 7934 1035 7980
rect 1081 7934 1193 7980
rect 1239 7934 1351 7980
rect 1397 7934 1509 7980
rect 1555 7934 1667 7980
rect 1713 7934 1826 7980
rect 1872 7934 1984 7980
rect 2030 7934 2142 7980
rect 2188 7934 2300 7980
rect 2346 7934 2458 7980
rect 2504 7934 2616 7980
rect 2662 7934 2774 7980
rect 2820 7934 2933 7980
rect 2979 7934 3091 7980
rect 3137 7934 3249 7980
rect 3295 7934 3407 7980
rect 3453 7934 3565 7980
rect 3611 7934 3723 7980
rect 3769 7934 3881 7980
rect 3927 7934 4039 7980
rect 4085 7934 4197 7980
rect 4243 7934 4292 7980
rect 4945 8120 5061 8543
rect 8947 8516 9451 8633
rect 8947 8470 8982 8516
rect 9028 8470 9140 8516
rect 9186 8470 9451 8516
rect 8947 8436 9451 8470
rect 8939 8395 9451 8436
rect 9497 8435 9532 9180
rect 9675 9180 9721 9193
rect 9636 8990 9675 9030
rect 9864 9180 9980 9412
rect 9864 9126 9899 9180
rect 9721 8990 9760 9030
rect 9636 8938 9672 8990
rect 9724 8938 9760 8990
rect 9636 8772 9675 8938
rect 9721 8772 9760 8938
rect 9636 8720 9672 8772
rect 9724 8720 9760 8772
rect 9636 8680 9675 8720
rect 9497 8395 9538 8435
rect 6862 8287 7702 8391
rect 6862 8200 6978 8287
rect 6862 8154 6897 8200
rect 6943 8154 6978 8200
rect 7121 8200 7167 8213
rect 5204 8124 5250 8133
rect 4945 8074 4980 8120
rect 5026 8074 5061 8120
rect 4945 8000 5061 8074
rect 4945 7954 4980 8000
rect 5026 7954 5061 8000
rect 4945 7949 5061 7954
rect 5169 8120 5285 8124
rect 5169 8074 5204 8120
rect 5250 8074 5285 8120
rect 5169 8000 5285 8074
rect 5169 7954 5204 8000
rect 5250 7970 5285 8000
rect 6862 8080 6978 8154
rect 6862 8034 6897 8080
rect 6943 8034 6978 8080
rect 5250 7954 5713 7970
rect 4980 7941 5026 7949
rect 355 7822 4292 7934
rect 355 7770 457 7822
rect 509 7770 668 7822
rect 720 7770 878 7822
rect 930 7770 1089 7822
rect 1141 7770 1300 7822
rect 1352 7770 1511 7822
rect 1563 7770 1722 7822
rect 1774 7770 1932 7822
rect 1984 7770 2143 7822
rect 2195 7770 2355 7822
rect 2407 7770 2566 7822
rect 2618 7770 2776 7822
rect 2828 7770 2987 7822
rect 3039 7770 3198 7822
rect 3250 7770 3409 7822
rect 3461 7770 3620 7822
rect 3672 7770 3830 7822
rect 3882 7770 4041 7822
rect 4093 7770 4292 7822
rect 355 7730 4292 7770
rect 5169 7913 5713 7954
rect 5169 7861 5411 7913
rect 5463 7861 5623 7913
rect 5675 7861 5713 7913
rect 5169 7786 5713 7861
rect 4980 7641 5026 7649
rect 4945 7636 5061 7641
rect 4945 7590 4980 7636
rect 5026 7590 5061 7636
rect 4945 7509 5061 7590
rect 4945 7463 4980 7509
rect 5026 7463 5061 7509
rect 4945 7382 5061 7463
rect 4945 7336 4980 7382
rect 5026 7336 5061 7382
rect 4945 7254 5061 7336
rect 4945 7208 4980 7254
rect 5026 7208 5061 7254
rect 4945 7106 5061 7208
rect 5169 7636 5285 7786
rect 5169 7590 5204 7636
rect 5250 7590 5285 7636
rect 6673 7729 6719 7742
rect 6673 7616 6719 7683
rect 6862 7729 6978 8034
rect 7082 8154 7121 8193
rect 7411 8200 7457 8213
rect 7167 8154 7206 8193
rect 7082 8153 7206 8154
rect 7082 8101 7118 8153
rect 7170 8101 7206 8153
rect 7082 8080 7206 8101
rect 7082 8034 7121 8080
rect 7167 8034 7206 8080
rect 7411 8080 7457 8154
rect 7082 7935 7206 8034
rect 7082 7883 7118 7935
rect 7170 7883 7206 7935
rect 7082 7843 7206 7883
rect 7376 8034 7411 8051
rect 7600 8200 7702 8287
rect 7600 8154 7635 8200
rect 7681 8154 7702 8200
rect 7600 8080 7702 8154
rect 8939 8343 8977 8395
rect 9029 8353 9189 8395
rect 9029 8343 9140 8353
rect 8939 8307 8982 8343
rect 9028 8307 9140 8343
rect 9186 8343 9189 8353
rect 9241 8343 9448 8395
rect 9500 8343 9538 8395
rect 9186 8307 9451 8343
rect 8939 8190 9451 8307
rect 8939 8178 8982 8190
rect 9028 8178 9140 8190
rect 8939 8126 8977 8178
rect 9029 8144 9140 8178
rect 9186 8178 9451 8190
rect 9497 8178 9538 8343
rect 9186 8144 9189 8178
rect 9029 8126 9189 8144
rect 9241 8126 9448 8178
rect 9500 8126 9538 8178
rect 7457 8034 7492 8051
rect 6862 7683 6897 7729
rect 6943 7683 6978 7729
rect 5169 7509 5285 7590
rect 5169 7463 5204 7509
rect 5250 7463 5285 7509
rect 5169 7382 5285 7463
rect 6638 7573 6754 7616
rect 6638 7527 6673 7573
rect 6719 7527 6754 7573
rect 6862 7573 6978 7683
rect 7121 7729 7167 7742
rect 7121 7616 7167 7683
rect 7376 7729 7492 8034
rect 7376 7683 7411 7729
rect 7457 7683 7492 7729
rect 6862 7548 6897 7573
rect 6638 7444 6754 7527
rect 6943 7548 6978 7573
rect 7086 7573 7202 7616
rect 6897 7514 6943 7527
rect 7086 7527 7121 7573
rect 7167 7527 7202 7573
rect 7086 7444 7202 7527
rect 5169 7336 5204 7382
rect 5250 7336 5285 7382
rect 5169 7254 5285 7336
rect 6154 7391 6494 7432
rect 6154 7339 6192 7391
rect 6286 7345 6398 7391
rect 6244 7339 6404 7345
rect 6456 7339 6494 7391
rect 6638 7342 7202 7444
rect 6154 7298 6494 7339
rect 5169 7208 5204 7254
rect 5250 7208 5285 7254
rect 5169 7204 5285 7208
rect 6673 7258 6719 7271
rect 6897 7262 6943 7271
rect 5204 7195 5250 7204
rect 6673 7152 6719 7212
rect 4944 7104 5061 7106
rect 4938 7065 5066 7104
rect 4938 7013 4976 7065
rect 5028 7013 5066 7065
rect 704 6914 4456 6951
rect 704 6868 739 6914
rect 785 6868 897 6914
rect 943 6868 1055 6914
rect 1101 6868 1213 6914
rect 1259 6868 1371 6914
rect 1417 6868 1529 6914
rect 1575 6868 1687 6914
rect 1733 6868 1845 6914
rect 1891 6868 2003 6914
rect 2049 6868 2162 6914
rect 2208 6868 2320 6914
rect 2366 6868 2478 6914
rect 2524 6868 2636 6914
rect 2682 6868 2794 6914
rect 2840 6868 2952 6914
rect 2998 6868 3111 6914
rect 3157 6868 3269 6914
rect 3315 6868 3427 6914
rect 3473 6868 3585 6914
rect 3631 6868 3743 6914
rect 3789 6868 3901 6914
rect 3947 6868 4059 6914
rect 4105 6868 4217 6914
rect 4263 6868 4375 6914
rect 4421 6868 4456 6914
rect 704 6861 4456 6868
rect 704 6809 743 6861
rect 795 6809 954 6861
rect 1006 6809 1164 6861
rect 1216 6809 1375 6861
rect 1427 6809 1586 6861
rect 1638 6809 1797 6861
rect 1849 6809 2008 6861
rect 2060 6809 2218 6861
rect 2270 6809 2429 6861
rect 2481 6809 2641 6861
rect 2693 6809 2852 6861
rect 2904 6809 3062 6861
rect 3114 6809 3273 6861
rect 3325 6809 3484 6861
rect 3536 6809 3695 6861
rect 3747 6809 3906 6861
rect 3958 6809 4116 6861
rect 4168 6809 4327 6861
rect 4379 6809 4456 6861
rect 704 6751 4456 6809
rect 704 6705 739 6751
rect 785 6705 897 6751
rect 943 6705 1055 6751
rect 1101 6705 1213 6751
rect 1259 6705 1371 6751
rect 1417 6705 1529 6751
rect 1575 6705 1687 6751
rect 1733 6705 1845 6751
rect 1891 6705 2003 6751
rect 2049 6705 2162 6751
rect 2208 6705 2320 6751
rect 2366 6705 2478 6751
rect 2524 6705 2636 6751
rect 2682 6705 2794 6751
rect 2840 6705 2952 6751
rect 2998 6705 3111 6751
rect 3157 6705 3269 6751
rect 3315 6705 3427 6751
rect 3473 6705 3585 6751
rect 3631 6705 3743 6751
rect 3789 6705 3901 6751
rect 3947 6705 4059 6751
rect 4105 6705 4217 6751
rect 4263 6705 4375 6751
rect 4421 6705 4456 6751
rect 704 6643 4456 6705
rect 704 6591 743 6643
rect 795 6591 954 6643
rect 1006 6591 1164 6643
rect 1216 6591 1375 6643
rect 1427 6591 1586 6643
rect 1638 6591 1797 6643
rect 1849 6591 2008 6643
rect 2060 6591 2218 6643
rect 2270 6591 2429 6643
rect 2481 6591 2641 6643
rect 2693 6591 2852 6643
rect 2904 6591 3062 6643
rect 3114 6591 3273 6643
rect 3325 6591 3484 6643
rect 3536 6591 3695 6643
rect 3747 6591 3906 6643
rect 3958 6591 4116 6643
rect 4168 6591 4327 6643
rect 4379 6591 4456 6643
rect 704 6588 4456 6591
rect 704 6542 739 6588
rect 785 6542 897 6588
rect 943 6542 1055 6588
rect 1101 6542 1213 6588
rect 1259 6542 1371 6588
rect 1417 6542 1529 6588
rect 1575 6542 1687 6588
rect 1733 6542 1845 6588
rect 1891 6542 2003 6588
rect 2049 6542 2162 6588
rect 2208 6542 2320 6588
rect 2366 6542 2478 6588
rect 2524 6542 2636 6588
rect 2682 6542 2794 6588
rect 2840 6542 2952 6588
rect 2998 6542 3111 6588
rect 3157 6542 3269 6588
rect 3315 6542 3427 6588
rect 3473 6542 3585 6588
rect 3631 6542 3743 6588
rect 3789 6542 3901 6588
rect 3947 6542 4059 6588
rect 4105 6542 4217 6588
rect 4263 6542 4375 6588
rect 4421 6542 4456 6588
rect 704 6505 4456 6542
rect 4938 6847 5066 7013
rect 5221 7078 5509 7115
rect 5221 7032 5256 7078
rect 5302 7032 5509 7078
rect 6673 7046 6719 7106
rect 5221 6993 5509 7032
rect 4938 6795 4976 6847
rect 5028 6795 5066 6847
rect 4938 6629 5066 6795
rect 4938 6577 4976 6629
rect 5028 6577 5066 6629
rect 4938 6537 5066 6577
rect 5393 6770 5509 6993
rect 6348 7000 6673 7036
rect 6858 7258 6982 7262
rect 6858 7222 6897 7258
rect 6943 7222 6982 7258
rect 6858 7170 6894 7222
rect 6946 7170 6982 7222
rect 6858 7152 6982 7170
rect 6858 7106 6897 7152
rect 6943 7106 6982 7152
rect 7086 7258 7202 7342
rect 7086 7212 7121 7258
rect 7167 7212 7202 7258
rect 7086 7152 7202 7212
rect 7086 7115 7121 7152
rect 6858 7046 6982 7106
rect 6719 7000 6754 7036
rect 6348 6969 6754 7000
rect 6348 6923 6383 6969
rect 6429 6940 6754 6969
rect 6429 6923 6673 6940
rect 6348 6894 6673 6923
rect 6719 6894 6754 6940
rect 6858 7004 6897 7046
rect 6943 7004 6982 7046
rect 6858 6952 6894 7004
rect 6946 6952 6982 7004
rect 6858 6940 6982 6952
rect 6858 6912 6897 6940
rect 6348 6857 6754 6894
rect 6348 6805 6386 6857
rect 6438 6834 6754 6857
rect 6438 6805 6673 6834
rect 6348 6788 6673 6805
rect 6719 6788 6754 6834
rect 6348 6777 6754 6788
rect 5393 6730 5519 6770
rect 5393 6678 5431 6730
rect 5483 6678 5519 6730
rect 4945 6405 5061 6537
rect 4945 6359 4980 6405
rect 5026 6359 5061 6405
rect 4945 6224 5061 6359
rect 4945 6178 4980 6224
rect 5026 6178 5061 6224
rect 4945 6140 5061 6178
rect 5393 6512 5519 6678
rect 5393 6460 5431 6512
rect 5483 6460 5519 6512
rect 5393 6420 5519 6460
rect 6348 6731 6383 6777
rect 6429 6731 6754 6777
rect 6348 6728 6754 6731
rect 6348 6682 6673 6728
rect 6719 6682 6754 6728
rect 6348 6639 6754 6682
rect 6348 6587 6386 6639
rect 6438 6622 6754 6639
rect 6438 6587 6673 6622
rect 6348 6584 6673 6587
rect 6348 6538 6383 6584
rect 6429 6576 6673 6584
rect 6719 6576 6754 6622
rect 6429 6538 6754 6576
rect 6348 6516 6754 6538
rect 6348 6470 6673 6516
rect 6719 6470 6754 6516
rect 6348 6421 6754 6470
rect 5393 6405 5509 6420
rect 5393 6359 5428 6405
rect 5474 6359 5509 6405
rect 5393 6224 5509 6359
rect 5393 6178 5428 6224
rect 5474 6178 5509 6224
rect 4802 6024 5142 6061
rect 4802 6020 5054 6024
rect 5100 6020 5142 6024
rect 4802 5968 4840 6020
rect 4892 5968 5052 6020
rect 5104 5968 5142 6020
rect 704 5931 4456 5968
rect 704 5885 739 5931
rect 785 5885 897 5931
rect 943 5885 1055 5931
rect 1101 5885 1213 5931
rect 1259 5885 1371 5931
rect 1417 5885 1529 5931
rect 1575 5885 1687 5931
rect 1733 5885 1845 5931
rect 1891 5885 2003 5931
rect 2049 5885 2162 5931
rect 2208 5885 2320 5931
rect 2366 5885 2478 5931
rect 2524 5885 2636 5931
rect 2682 5885 2794 5931
rect 2840 5885 2952 5931
rect 2998 5885 3111 5931
rect 3157 5885 3269 5931
rect 3315 5885 3427 5931
rect 3473 5885 3585 5931
rect 3631 5885 3743 5931
rect 3789 5885 3901 5931
rect 3947 5885 4059 5931
rect 4105 5885 4217 5931
rect 4263 5885 4375 5931
rect 4421 5885 4456 5931
rect 4802 5928 5142 5968
rect 704 5877 4456 5885
rect 704 5825 743 5877
rect 795 5825 954 5877
rect 1006 5825 1164 5877
rect 1216 5825 1375 5877
rect 1427 5825 1586 5877
rect 1638 5825 1797 5877
rect 1849 5825 2008 5877
rect 2060 5825 2218 5877
rect 2270 5825 2429 5877
rect 2481 5825 2641 5877
rect 2693 5825 2852 5877
rect 2904 5825 3062 5877
rect 3114 5825 3273 5877
rect 3325 5825 3484 5877
rect 3536 5825 3695 5877
rect 3747 5825 3906 5877
rect 3958 5825 4116 5877
rect 4168 5825 4327 5877
rect 4379 5825 4456 5877
rect 5393 5848 5509 6178
rect 6348 6375 6383 6421
rect 6438 6410 6754 6421
rect 6348 6369 6386 6375
rect 6438 6369 6673 6410
rect 6348 6364 6673 6369
rect 6719 6364 6754 6410
rect 6348 6303 6754 6364
rect 6348 6257 6673 6303
rect 6719 6257 6754 6303
rect 6348 6196 6754 6257
rect 6348 6150 6673 6196
rect 6719 6150 6754 6196
rect 6862 6894 6897 6912
rect 6943 6912 6982 6940
rect 7080 7106 7121 7115
rect 7167 7115 7202 7152
rect 7376 7609 7492 7683
rect 7600 8034 7635 8080
rect 7681 8034 7702 8080
rect 7600 7729 7702 8034
rect 7795 8083 7919 8123
rect 7795 8031 7831 8083
rect 7883 8031 7919 8083
rect 7795 7985 7919 8031
rect 7795 7939 7828 7985
rect 7874 7939 7919 7985
rect 7795 7865 7919 7939
rect 7795 7821 7831 7865
rect 7795 7775 7828 7821
rect 7883 7813 7919 7865
rect 7874 7775 7919 7813
rect 7795 7773 7919 7775
rect 8939 8026 9451 8126
rect 8939 7980 8982 8026
rect 9028 7980 9140 8026
rect 9186 7980 9451 8026
rect 8939 7960 9451 7980
rect 9497 7960 9538 8126
rect 8939 7908 8977 7960
rect 9029 7908 9189 7960
rect 9241 7908 9448 7960
rect 9500 7908 9538 7960
rect 8939 7863 9451 7908
rect 8939 7817 8982 7863
rect 9028 7817 9140 7863
rect 9186 7817 9451 7863
rect 7795 7738 7907 7773
rect 8939 7743 9451 7817
rect 9497 7743 9538 7908
rect 7600 7683 7635 7729
rect 7681 7683 7702 7729
rect 7600 7614 7702 7683
rect 8939 7691 8977 7743
rect 9029 7700 9189 7743
rect 9029 7691 9140 7700
rect 8939 7654 8982 7691
rect 9028 7654 9140 7691
rect 9186 7691 9189 7700
rect 9241 7691 9448 7743
rect 9500 7691 9538 7743
rect 9186 7654 9451 7691
rect 7376 7563 7411 7609
rect 7457 7563 7492 7609
rect 7167 7106 7208 7115
rect 7080 7075 7208 7106
rect 7080 7023 7118 7075
rect 7170 7023 7208 7075
rect 7080 7000 7121 7023
rect 7167 7000 7208 7023
rect 7080 6940 7208 7000
rect 6943 6894 6978 6912
rect 6862 6834 6978 6894
rect 6862 6788 6897 6834
rect 6943 6788 6978 6834
rect 6862 6728 6978 6788
rect 6862 6682 6897 6728
rect 6943 6682 6978 6728
rect 6862 6622 6978 6682
rect 6862 6576 6897 6622
rect 6943 6576 6978 6622
rect 6862 6516 6978 6576
rect 6862 6470 6897 6516
rect 6943 6470 6978 6516
rect 6862 6410 6978 6470
rect 6862 6364 6897 6410
rect 6943 6364 6978 6410
rect 6862 6303 6978 6364
rect 7080 6894 7121 6940
rect 7167 6894 7208 6940
rect 7080 6857 7208 6894
rect 7080 6805 7118 6857
rect 7170 6805 7208 6857
rect 7080 6788 7121 6805
rect 7167 6788 7208 6805
rect 7080 6728 7208 6788
rect 7080 6682 7121 6728
rect 7167 6682 7208 6728
rect 7080 6639 7208 6682
rect 7080 6587 7118 6639
rect 7170 6587 7208 6639
rect 7080 6576 7121 6587
rect 7167 6576 7208 6587
rect 7080 6516 7208 6576
rect 7080 6470 7121 6516
rect 7167 6470 7208 6516
rect 7080 6421 7208 6470
rect 7080 6369 7118 6421
rect 7170 6369 7208 6421
rect 7080 6364 7121 6369
rect 7167 6364 7208 6369
rect 7080 6329 7208 6364
rect 7376 6818 7492 7563
rect 7635 7609 7681 7614
rect 7635 7550 7681 7563
rect 8939 7536 9451 7654
rect 8939 7525 8982 7536
rect 9028 7525 9140 7536
rect 8939 7473 8977 7525
rect 9029 7490 9140 7525
rect 9186 7525 9451 7536
rect 9497 7525 9538 7691
rect 9186 7490 9189 7525
rect 9029 7473 9189 7490
rect 9241 7473 9448 7525
rect 9500 7473 9538 7525
rect 7569 7468 7874 7469
rect 7569 7432 7919 7468
rect 7569 7386 7604 7432
rect 7650 7428 7919 7432
rect 7650 7386 7831 7428
rect 7569 7376 7831 7386
rect 7883 7376 7919 7428
rect 7569 7349 7919 7376
rect 7793 7210 7919 7349
rect 7793 7158 7831 7210
rect 7883 7158 7919 7210
rect 7793 7118 7919 7158
rect 8939 7373 9451 7473
rect 8939 7327 8982 7373
rect 9028 7327 9140 7373
rect 9186 7327 9451 7373
rect 8939 7307 9451 7327
rect 9497 7307 9538 7473
rect 8939 7255 8977 7307
rect 9029 7255 9189 7307
rect 9241 7255 9448 7307
rect 9500 7255 9538 7307
rect 8939 7210 9451 7255
rect 8939 7164 8982 7210
rect 9028 7164 9140 7210
rect 9186 7164 9451 7210
rect 7376 6772 7411 6818
rect 7457 6772 7492 6818
rect 7376 6691 7492 6772
rect 7376 6645 7411 6691
rect 7457 6645 7492 6691
rect 7376 6564 7492 6645
rect 7376 6518 7411 6564
rect 7457 6518 7492 6564
rect 7376 6436 7492 6518
rect 7376 6390 7411 6436
rect 7457 6390 7492 6436
rect 6862 6257 6897 6303
rect 6943 6257 6978 6303
rect 6862 6196 6978 6257
rect 6862 6158 6897 6196
rect 6348 6145 6754 6150
rect 6855 6150 6897 6158
rect 6943 6158 6978 6196
rect 7121 6303 7167 6329
rect 7121 6196 7167 6257
rect 6943 6150 6985 6158
rect 6673 6137 6719 6145
rect 6855 6118 6985 6150
rect 7121 6137 7167 6150
rect 6855 6066 6894 6118
rect 6946 6066 6985 6118
rect 6350 5970 6474 6010
rect 6350 5918 6386 5970
rect 6438 5918 6474 5970
rect 6350 5848 6474 5918
rect 6855 5900 6985 6066
rect 7376 6054 7492 6390
rect 7099 6017 7492 6054
rect 7099 5971 7134 6017
rect 7180 5971 7492 6017
rect 7099 5934 7492 5971
rect 6673 5848 6719 5856
rect 6855 5848 6894 5900
rect 6946 5848 6985 5900
rect 704 5768 4456 5825
rect 704 5722 739 5768
rect 785 5722 897 5768
rect 943 5722 1055 5768
rect 1101 5722 1213 5768
rect 1259 5722 1371 5768
rect 1417 5722 1529 5768
rect 1575 5722 1687 5768
rect 1733 5722 1845 5768
rect 1891 5722 2003 5768
rect 2049 5722 2162 5768
rect 2208 5722 2320 5768
rect 2366 5722 2478 5768
rect 2524 5722 2636 5768
rect 2682 5722 2794 5768
rect 2840 5722 2952 5768
rect 2998 5722 3111 5768
rect 3157 5722 3269 5768
rect 3315 5722 3427 5768
rect 3473 5722 3585 5768
rect 3631 5722 3743 5768
rect 3789 5722 3901 5768
rect 3947 5722 4059 5768
rect 4105 5722 4217 5768
rect 4263 5722 4375 5768
rect 4421 5722 4456 5768
rect 704 5659 4456 5722
rect 704 5607 743 5659
rect 795 5607 954 5659
rect 1006 5607 1164 5659
rect 1216 5607 1375 5659
rect 1427 5607 1586 5659
rect 1638 5607 1797 5659
rect 1849 5607 2008 5659
rect 2060 5607 2218 5659
rect 2270 5607 2429 5659
rect 2481 5607 2641 5659
rect 2693 5607 2852 5659
rect 2904 5607 3062 5659
rect 3114 5607 3273 5659
rect 3325 5607 3484 5659
rect 3536 5607 3695 5659
rect 3747 5607 3906 5659
rect 3958 5607 4116 5659
rect 4168 5607 4327 5659
rect 4379 5607 4456 5659
rect 4945 5746 5509 5848
rect 4945 5661 5061 5746
rect 5204 5666 5250 5674
rect 4945 5639 4980 5661
rect 704 5605 4456 5607
rect 704 5559 739 5605
rect 785 5559 897 5605
rect 943 5559 1055 5605
rect 1101 5559 1213 5605
rect 1259 5559 1371 5605
rect 1417 5559 1529 5605
rect 1575 5559 1687 5605
rect 1733 5559 1845 5605
rect 1891 5559 2003 5605
rect 2049 5559 2162 5605
rect 2208 5559 2320 5605
rect 2366 5559 2478 5605
rect 2524 5559 2636 5605
rect 2682 5559 2794 5605
rect 2840 5559 2952 5605
rect 2998 5559 3111 5605
rect 3157 5559 3269 5605
rect 3315 5559 3427 5605
rect 3473 5559 3585 5605
rect 3631 5559 3743 5605
rect 3789 5559 3901 5605
rect 3947 5559 4059 5605
rect 4105 5559 4217 5605
rect 4263 5559 4375 5605
rect 4421 5559 4456 5605
rect 704 5522 4456 5559
rect 5026 5639 5061 5661
rect 5164 5661 5288 5666
rect 4980 5402 5026 5415
rect 5164 5626 5204 5661
rect 5250 5626 5288 5661
rect 5164 5574 5200 5626
rect 5252 5574 5288 5626
rect 5393 5661 5509 5746
rect 5393 5621 5428 5661
rect 5164 5415 5204 5574
rect 5250 5415 5288 5574
rect 5164 5408 5288 5415
rect 5164 5356 5200 5408
rect 5252 5356 5288 5408
rect 5474 5621 5509 5661
rect 5751 5811 5880 5848
rect 5751 5765 5788 5811
rect 5834 5807 5880 5811
rect 5751 5755 5789 5765
rect 5841 5755 5880 5807
rect 5751 5589 5880 5755
rect 5751 5537 5789 5589
rect 5841 5537 5880 5589
rect 5751 5497 5880 5537
rect 6348 5843 6754 5848
rect 6348 5797 6673 5843
rect 6719 5797 6754 5843
rect 6855 5843 6985 5848
rect 6855 5807 6897 5843
rect 6348 5752 6754 5797
rect 6348 5707 6386 5752
rect 6438 5716 6754 5752
rect 6862 5797 6897 5807
rect 6943 5807 6985 5843
rect 7121 5843 7167 5856
rect 6943 5797 6978 5807
rect 6862 5737 6978 5797
rect 7121 5757 7167 5797
rect 7376 5843 7492 5934
rect 7376 5797 7411 5843
rect 7457 5797 7492 5843
rect 7376 5759 7492 5797
rect 7569 6818 7681 6831
rect 7569 6772 7635 6818
rect 7569 6691 7681 6772
rect 7569 6645 7635 6691
rect 7569 6564 7681 6645
rect 7569 6518 7635 6564
rect 7569 6436 7681 6518
rect 7569 6390 7635 6436
rect 7569 6377 7681 6390
rect 7569 5856 7680 6377
rect 7793 6069 7874 7118
rect 8939 7089 9451 7164
rect 9497 7089 9538 7255
rect 8939 7037 8977 7089
rect 9029 7046 9189 7089
rect 9029 7037 9140 7046
rect 8939 7000 8982 7037
rect 9028 7000 9140 7037
rect 9186 7037 9189 7046
rect 9241 7037 9448 7089
rect 9500 7037 9538 7089
rect 9186 7000 9451 7037
rect 8939 6883 9451 7000
rect 8939 6872 8982 6883
rect 9028 6872 9140 6883
rect 8939 6820 8977 6872
rect 9029 6837 9140 6872
rect 9186 6872 9451 6883
rect 9497 6872 9538 7037
rect 9186 6837 9189 6872
rect 9029 6820 9189 6837
rect 9241 6820 9448 6872
rect 9500 6820 9538 6872
rect 8939 6720 9451 6820
rect 8939 6674 8982 6720
rect 9028 6674 9140 6720
rect 9186 6674 9451 6720
rect 8939 6654 9451 6674
rect 9497 6654 9538 6820
rect 8939 6602 8977 6654
rect 9029 6602 9189 6654
rect 9241 6602 9448 6654
rect 9500 6602 9538 6654
rect 8939 6557 9451 6602
rect 8939 6511 8982 6557
rect 9028 6511 9140 6557
rect 9186 6511 9451 6557
rect 8939 6437 9451 6511
rect 9497 6437 9538 6602
rect 8939 6385 8977 6437
rect 9029 6394 9189 6437
rect 9029 6385 9140 6394
rect 8939 6348 8982 6385
rect 9028 6348 9140 6385
rect 9186 6385 9189 6394
rect 9241 6385 9448 6437
rect 9500 6385 9538 6437
rect 9186 6348 9451 6385
rect 8939 6344 9451 6348
rect 7758 6033 7874 6069
rect 7758 5987 7793 6033
rect 7839 5987 7874 6033
rect 7758 5950 7874 5987
rect 8947 6230 9451 6344
rect 8947 6184 8982 6230
rect 9028 6184 9140 6230
rect 9186 6184 9451 6230
rect 8947 6067 9451 6184
rect 8947 6021 8982 6067
rect 9028 6021 9140 6067
rect 9186 6021 9451 6067
rect 8947 5904 9451 6021
rect 8947 5858 8982 5904
rect 9028 5858 9140 5904
rect 9186 5858 9451 5904
rect 7569 5843 7681 5856
rect 7569 5797 7635 5843
rect 6348 5661 6383 5707
rect 6438 5700 6673 5716
rect 6429 5670 6673 5700
rect 6719 5670 6754 5716
rect 6429 5661 6754 5670
rect 6348 5589 6754 5661
rect 6348 5543 6673 5589
rect 6719 5543 6754 5589
rect 6348 5497 6383 5543
rect 6429 5501 6754 5543
rect 6897 5716 6943 5737
rect 6897 5589 6943 5670
rect 6429 5497 6464 5501
rect 5428 5402 5474 5415
rect 5164 5316 5288 5356
rect 5168 5315 5285 5316
rect 5169 5165 5285 5315
rect 6348 5165 6464 5497
rect 6673 5461 6719 5501
rect 6673 5402 6719 5415
rect 6897 5461 6943 5543
rect 6897 5402 6943 5415
rect 7086 5716 7202 5757
rect 7086 5670 7121 5716
rect 7167 5670 7202 5716
rect 7086 5589 7202 5670
rect 7086 5543 7121 5589
rect 7167 5543 7202 5589
rect 7086 5461 7202 5543
rect 7086 5415 7121 5461
rect 7167 5415 7202 5461
rect 7086 5165 7202 5415
rect 7411 5716 7457 5759
rect 7411 5589 7457 5670
rect 7411 5461 7457 5543
rect 7411 5402 7457 5415
rect 7569 5716 7681 5797
rect 8947 5741 9451 5858
rect 7569 5670 7635 5716
rect 7681 5670 8811 5716
rect 7569 5596 8811 5670
rect 8947 5695 8982 5741
rect 9028 5695 9140 5741
rect 9186 5695 9451 5741
rect 8947 5659 9451 5695
rect 8948 5658 9451 5659
rect 9416 5657 9451 5658
rect 7569 5589 7681 5596
rect 7569 5543 7635 5589
rect 7569 5461 7681 5543
rect 7569 5415 7635 5461
rect 7569 5410 7681 5415
rect 7635 5402 7681 5410
rect 8696 5249 8811 5596
rect 9497 6344 9538 6385
rect 9497 5657 9532 6344
rect 9451 5293 9497 5306
rect 9721 8680 9760 8720
rect 9858 8395 9899 8436
rect 9945 9126 9980 9180
rect 10123 9180 10300 9193
rect 10086 8990 10123 9030
rect 10169 8990 10300 9180
rect 10650 9182 10696 9195
rect 10086 8938 10122 8990
rect 10174 8938 10300 8990
rect 10086 8772 10123 8938
rect 10169 8772 10300 8938
rect 10086 8720 10122 8772
rect 10174 8720 10300 8772
rect 10086 8680 10123 8720
rect 9945 8435 9977 8436
rect 9945 8395 9986 8435
rect 9858 8343 9896 8395
rect 9948 8343 9986 8395
rect 9858 8178 9899 8343
rect 9945 8178 9986 8343
rect 9858 8126 9896 8178
rect 9948 8126 9986 8178
rect 9858 7960 9899 8126
rect 9945 7960 9986 8126
rect 9858 7908 9896 7960
rect 9948 7908 9986 7960
rect 9858 7743 9899 7908
rect 9945 7743 9986 7908
rect 9858 7691 9896 7743
rect 9948 7691 9986 7743
rect 9858 7525 9899 7691
rect 9945 7525 9986 7691
rect 9858 7473 9896 7525
rect 9948 7473 9986 7525
rect 9858 7307 9899 7473
rect 9945 7307 9986 7473
rect 9858 7255 9896 7307
rect 9948 7255 9986 7307
rect 9858 7089 9899 7255
rect 9945 7089 9986 7255
rect 9858 7037 9896 7089
rect 9948 7037 9986 7089
rect 9858 6872 9899 7037
rect 9945 6872 9986 7037
rect 9858 6820 9896 6872
rect 9948 6820 9986 6872
rect 9858 6654 9899 6820
rect 9945 6654 9986 6820
rect 9858 6602 9896 6654
rect 9948 6602 9986 6654
rect 9858 6437 9899 6602
rect 9945 6437 9986 6602
rect 9858 6385 9896 6437
rect 9948 6385 9986 6437
rect 9858 6344 9899 6385
rect 9675 5293 9721 5306
rect 9945 6344 9986 6385
rect 9899 5293 9945 5306
rect 10169 5306 10300 8720
rect 10123 5293 10300 5306
rect 8585 5208 8925 5249
rect 67 4997 8120 5165
rect 8585 5156 8623 5208
rect 8675 5156 8835 5208
rect 8887 5156 8925 5208
rect 9752 5201 9868 5202
rect 9978 5201 10094 5202
rect 8585 5115 8925 5156
rect 9745 5161 9875 5201
rect 9745 5109 9784 5161
rect 9836 5109 9875 5161
rect 9557 5095 9625 5106
rect 9557 5002 9568 5095
rect 67 4937 314 4997
rect 67 4885 255 4937
rect 307 4885 314 4937
rect 67 4719 314 4885
rect 67 4667 255 4719
rect 307 4667 314 4719
rect 67 4501 314 4667
rect 67 4449 255 4501
rect 307 4449 314 4501
rect 67 4351 314 4449
rect 7760 4380 8120 4997
rect 7760 4351 8039 4380
rect 67 4334 8039 4351
rect 8085 4334 8120 4380
rect 67 4283 8120 4334
rect 67 4231 255 4283
rect 307 4231 466 4283
rect 518 4231 677 4283
rect 729 4231 887 4283
rect 939 4231 1098 4283
rect 1150 4231 1309 4283
rect 1361 4231 1520 4283
rect 1572 4231 1731 4283
rect 1783 4231 1941 4283
rect 1993 4231 2152 4283
rect 2204 4231 2363 4283
rect 2415 4231 2574 4283
rect 2626 4231 2785 4283
rect 2837 4231 2996 4283
rect 3048 4231 3207 4283
rect 3259 4231 3418 4283
rect 3470 4231 3629 4283
rect 3681 4231 3839 4283
rect 3891 4231 4050 4283
rect 4102 4231 4261 4283
rect 4313 4231 4472 4283
rect 4524 4231 4683 4283
rect 4735 4231 4893 4283
rect 4945 4231 5104 4283
rect 5156 4231 5315 4283
rect 5367 4273 8120 4283
rect 8228 4955 9568 5002
rect 9614 4955 9625 5095
rect 8228 4882 9625 4955
rect 9745 5095 9875 5109
rect 9745 4955 9791 5095
rect 9837 4955 9875 5095
rect 9745 4943 9875 4955
rect 9745 4891 9784 4943
rect 9836 4891 9875 4943
rect 8228 4380 8344 4882
rect 9745 4850 9875 4891
rect 9971 5161 10101 5201
rect 9971 5109 10010 5161
rect 10062 5109 10101 5161
rect 9971 5095 10101 5109
rect 9971 4955 10015 5095
rect 10061 4955 10101 5095
rect 9971 4943 10101 4955
rect 9971 4891 10010 4943
rect 10062 4891 10101 4943
rect 9971 4850 10101 4891
rect 8228 4334 8263 4380
rect 8309 4334 8344 4380
rect 8228 4281 8344 4334
rect 8878 4775 9532 4789
rect 8878 4752 9545 4775
rect 8878 4720 9451 4752
rect 9497 4734 9545 4752
rect 8878 4674 8926 4720
rect 8972 4701 9084 4720
rect 8972 4674 8981 4701
rect 8878 4649 8981 4674
rect 9033 4674 9084 4701
rect 9130 4706 9451 4720
rect 9130 4701 9454 4706
rect 9130 4674 9193 4701
rect 9033 4649 9193 4674
rect 9245 4682 9454 4701
rect 9506 4682 9545 4734
rect 10184 4696 10300 5293
rect 10608 9097 10650 9137
rect 10839 9182 10955 9412
rect 10696 9097 10738 9137
rect 10839 9126 10874 9182
rect 10608 9045 10647 9097
rect 10699 9045 10738 9097
rect 10608 8879 10650 9045
rect 10696 8879 10738 9045
rect 10608 8827 10647 8879
rect 10699 8827 10738 8879
rect 10608 8661 10650 8827
rect 10696 8661 10738 8827
rect 10608 8609 10647 8661
rect 10699 8609 10738 8661
rect 10608 8444 10650 8609
rect 10696 8444 10738 8609
rect 10608 8392 10647 8444
rect 10699 8392 10738 8444
rect 10608 8226 10650 8392
rect 10696 8226 10738 8392
rect 10608 8174 10647 8226
rect 10699 8174 10738 8226
rect 10608 8008 10650 8174
rect 10696 8008 10738 8174
rect 10608 7956 10647 8008
rect 10699 7956 10738 8008
rect 10608 7791 10650 7956
rect 10696 7791 10738 7956
rect 10608 7739 10647 7791
rect 10699 7739 10738 7791
rect 10608 7573 10650 7739
rect 10696 7573 10738 7739
rect 10608 7521 10647 7573
rect 10699 7521 10738 7573
rect 10608 7356 10650 7521
rect 10696 7356 10738 7521
rect 10608 7304 10647 7356
rect 10699 7304 10738 7356
rect 10608 7138 10650 7304
rect 10696 7138 10738 7304
rect 10608 7086 10647 7138
rect 10699 7086 10738 7138
rect 10608 6920 10650 7086
rect 10696 6920 10738 7086
rect 10608 6868 10647 6920
rect 10699 6868 10738 6920
rect 10608 6702 10650 6868
rect 10696 6702 10738 6868
rect 10608 6650 10647 6702
rect 10699 6650 10738 6702
rect 10608 6485 10650 6650
rect 10696 6485 10738 6650
rect 10608 6433 10647 6485
rect 10699 6433 10738 6485
rect 10608 6267 10650 6433
rect 10696 6267 10738 6433
rect 10833 8386 10874 8427
rect 10920 9126 10955 9182
rect 11098 9182 11144 9195
rect 11056 9097 11098 9137
rect 11287 9182 11403 9412
rect 11144 9097 11186 9137
rect 11287 9126 11322 9182
rect 11056 9045 11095 9097
rect 11147 9045 11186 9097
rect 11056 8879 11098 9045
rect 11144 8879 11186 9045
rect 11056 8827 11095 8879
rect 11147 8827 11186 8879
rect 11056 8661 11098 8827
rect 11144 8661 11186 8827
rect 11056 8609 11095 8661
rect 11147 8609 11186 8661
rect 11056 8444 11098 8609
rect 11144 8444 11186 8609
rect 10920 8426 10952 8427
rect 10920 8386 10961 8426
rect 10833 8334 10871 8386
rect 10923 8334 10961 8386
rect 10833 8169 10874 8334
rect 10920 8169 10961 8334
rect 10833 8117 10871 8169
rect 10923 8117 10961 8169
rect 10833 7951 10874 8117
rect 10920 7951 10961 8117
rect 10833 7899 10871 7951
rect 10923 7899 10961 7951
rect 10833 7734 10874 7899
rect 10920 7734 10961 7899
rect 10833 7682 10871 7734
rect 10923 7682 10961 7734
rect 10833 7516 10874 7682
rect 10920 7516 10961 7682
rect 10833 7464 10871 7516
rect 10923 7464 10961 7516
rect 10833 7298 10874 7464
rect 10920 7298 10961 7464
rect 10833 7246 10871 7298
rect 10923 7246 10961 7298
rect 10833 7080 10874 7246
rect 10920 7080 10961 7246
rect 10833 7028 10871 7080
rect 10923 7028 10961 7080
rect 10833 6863 10874 7028
rect 10920 6863 10961 7028
rect 10833 6811 10871 6863
rect 10923 6811 10961 6863
rect 10833 6645 10874 6811
rect 10920 6645 10961 6811
rect 10833 6593 10871 6645
rect 10923 6593 10961 6645
rect 10833 6428 10874 6593
rect 10920 6428 10961 6593
rect 10833 6376 10871 6428
rect 10923 6376 10961 6428
rect 10833 6335 10874 6376
rect 10608 6215 10647 6267
rect 10699 6215 10738 6267
rect 10608 6050 10650 6215
rect 10696 6050 10738 6215
rect 10608 5998 10647 6050
rect 10699 5998 10738 6050
rect 10608 5832 10650 5998
rect 10696 5832 10738 5998
rect 10608 5780 10647 5832
rect 10699 5780 10738 5832
rect 10608 5614 10650 5780
rect 10696 5614 10738 5780
rect 10608 5562 10647 5614
rect 10699 5562 10738 5614
rect 10608 5397 10650 5562
rect 10696 5397 10738 5562
rect 10608 5345 10647 5397
rect 10699 5345 10738 5397
rect 10608 5179 10650 5345
rect 10696 5179 10738 5345
rect 10608 5127 10647 5179
rect 10699 5127 10738 5179
rect 10608 4961 10650 5127
rect 10696 4961 10738 5127
rect 10608 4909 10647 4961
rect 10699 4909 10738 4961
rect 10608 4869 10650 4909
rect 9245 4649 9545 4682
rect 8878 4584 9545 4649
rect 8878 4557 9451 4584
rect 8878 4511 8926 4557
rect 8972 4511 9084 4557
rect 9130 4538 9451 4557
rect 9497 4538 9545 4584
rect 9130 4517 9545 4538
rect 9130 4511 9454 4517
rect 8878 4483 9454 4511
rect 8878 4431 8981 4483
rect 9033 4431 9193 4483
rect 9245 4465 9454 4483
rect 9506 4465 9545 4517
rect 9245 4431 9545 4465
rect 8878 4417 9545 4431
rect 8878 4394 9451 4417
rect 8878 4348 8926 4394
rect 8972 4348 9084 4394
rect 9130 4371 9451 4394
rect 9497 4371 9545 4417
rect 9130 4348 9545 4371
rect 8878 4299 9545 4348
rect 5367 4231 8039 4273
rect 67 4227 8039 4231
rect 8085 4227 8120 4273
rect 67 4191 8120 4227
rect 5082 3855 5128 4191
rect 5082 3772 5128 3809
rect 5386 3855 5859 3892
rect 5386 3809 5426 3855
rect 5472 3809 5859 3855
rect 5386 3772 5859 3809
rect 6127 3855 6242 4191
rect 6127 3809 6160 3855
rect 6206 3809 6242 3855
rect 6127 3772 6242 3809
rect 6504 3855 6619 3918
rect 6550 3809 6619 3855
rect 5324 3594 5664 3599
rect 5310 3558 5664 3594
rect 5310 3557 5362 3558
rect 5414 3557 5574 3558
rect 5310 3511 5345 3557
rect 5414 3511 5503 3557
rect 5549 3511 5574 3557
rect 5310 3506 5362 3511
rect 5414 3506 5574 3511
rect 5626 3506 5664 3558
rect 5310 3474 5664 3506
rect 5324 3466 5664 3474
rect 5743 3594 5859 3772
rect 6504 3594 6619 3809
rect 6848 3860 6925 4191
rect 6848 3814 6879 3860
rect 6848 3777 6925 3814
rect 7183 3860 7299 3918
rect 7229 3814 7299 3860
rect 7183 3594 7299 3814
rect 7490 3888 7606 4191
rect 8004 4166 8120 4191
rect 8004 4120 8039 4166
rect 8085 4120 8120 4166
rect 8004 4060 8120 4120
rect 8004 4014 8039 4060
rect 8085 4014 8120 4060
rect 8004 3954 8120 4014
rect 7490 3842 7525 3888
rect 7571 3842 7606 3888
rect 7490 3789 7606 3842
rect 7749 3888 7795 3941
rect 7749 3594 7795 3842
rect 8004 3908 8039 3954
rect 8085 3908 8120 3954
rect 8004 3848 8120 3908
rect 8004 3802 8039 3848
rect 8085 3802 8120 3848
rect 8004 3789 8120 3802
rect 8263 4273 8309 4281
rect 8263 4166 8309 4227
rect 8263 4060 8309 4120
rect 8263 3954 8309 4014
rect 8263 3848 8309 3908
rect 5743 3557 6264 3594
rect 5743 3511 6183 3557
rect 6229 3511 6264 3557
rect 5743 3474 6264 3511
rect 6504 3557 6987 3594
rect 6504 3511 6907 3557
rect 6953 3511 6987 3557
rect 6504 3474 6987 3511
rect 7183 3593 7598 3594
rect 7183 3557 7627 3593
rect 7183 3511 7547 3557
rect 7593 3511 7627 3557
rect 7183 3474 7627 3511
rect 7749 3557 8146 3594
rect 7749 3511 8065 3557
rect 8111 3511 8146 3557
rect 7749 3474 8146 3511
rect 5743 3260 5859 3474
rect 5082 3247 5128 3260
rect 5082 3139 5128 3201
rect 5082 2742 5128 3093
rect 5426 3247 5859 3260
rect 5472 3201 5859 3247
rect 5426 3139 5859 3201
rect 5472 3093 5859 3139
rect 5426 3080 5859 3093
rect 6117 3247 6233 3260
rect 6504 3252 6619 3474
rect 6117 3201 6160 3247
rect 6206 3201 6233 3247
rect 6117 3139 6233 3201
rect 6117 3093 6160 3139
rect 6206 3093 6233 3139
rect 6117 2742 6233 3093
rect 6503 3247 6619 3252
rect 6503 3201 6504 3247
rect 6550 3201 6619 3247
rect 6503 3139 6619 3201
rect 6503 3093 6504 3139
rect 6550 3093 6619 3139
rect 6503 3050 6619 3093
rect 6841 3247 6957 3260
rect 6841 3201 6879 3247
rect 6925 3201 6957 3247
rect 6841 3139 6957 3201
rect 6841 3093 6879 3139
rect 6925 3093 6957 3139
rect 6841 2742 6957 3093
rect 7183 3247 7299 3474
rect 7229 3201 7299 3247
rect 7183 3139 7299 3201
rect 7229 3093 7299 3139
rect 7183 3080 7299 3093
rect 7490 3247 7606 3260
rect 7490 2895 7525 3247
rect 7571 2895 7606 3247
rect 7490 2751 7606 2895
rect 7749 3247 7795 3474
rect 7749 2882 7795 2895
rect 8004 3247 8120 3260
rect 8004 3201 8039 3247
rect 8085 3201 8120 3247
rect 8004 3133 8120 3201
rect 8004 3087 8039 3133
rect 8085 3087 8120 3133
rect 8004 3063 8120 3087
rect 7003 2742 7606 2751
rect 2514 2730 7606 2742
rect 2514 2678 2526 2730
rect 2578 2678 2658 2730
rect 2710 2678 2790 2730
rect 2842 2678 2922 2730
rect 2974 2678 3054 2730
rect 3106 2678 3186 2730
rect 3238 2678 3318 2730
rect 3370 2678 3450 2730
rect 3502 2678 3582 2730
rect 3634 2678 3714 2730
rect 3766 2719 3846 2730
rect 3898 2719 3978 2730
rect 4030 2719 4110 2730
rect 4162 2719 4242 2730
rect 4294 2719 4374 2730
rect 4426 2719 4506 2730
rect 4558 2719 4638 2730
rect 4690 2719 4770 2730
rect 4822 2719 4902 2730
rect 4954 2719 5034 2730
rect 5086 2719 5166 2730
rect 5218 2719 5298 2730
rect 5350 2719 5430 2730
rect 3766 2678 3772 2719
rect 2514 2673 3772 2678
rect 3818 2678 3846 2719
rect 3942 2678 3978 2719
rect 4066 2678 4110 2719
rect 4190 2678 4242 2719
rect 4314 2678 4374 2719
rect 4438 2678 4506 2719
rect 4562 2678 4638 2719
rect 4690 2678 4764 2719
rect 4822 2678 4888 2719
rect 4954 2678 5012 2719
rect 5086 2678 5136 2719
rect 5218 2678 5260 2719
rect 5350 2678 5384 2719
rect 3818 2673 3896 2678
rect 3942 2673 4020 2678
rect 4066 2673 4144 2678
rect 4190 2673 4268 2678
rect 4314 2673 4392 2678
rect 4438 2673 4516 2678
rect 4562 2673 4640 2678
rect 4686 2673 4764 2678
rect 4810 2673 4888 2678
rect 4934 2673 5012 2678
rect 5058 2673 5136 2678
rect 5182 2673 5260 2678
rect 5306 2673 5384 2678
rect 5482 2719 5562 2730
rect 5482 2678 5508 2719
rect 5430 2673 5508 2678
rect 5554 2678 5562 2719
rect 5614 2719 5694 2730
rect 5614 2678 5632 2719
rect 5554 2673 5632 2678
rect 5678 2678 5694 2719
rect 5746 2719 5826 2730
rect 5746 2678 5756 2719
rect 5678 2673 5756 2678
rect 5802 2678 5826 2719
rect 5878 2719 5958 2730
rect 6010 2719 6090 2730
rect 6142 2719 6222 2730
rect 6274 2719 6354 2730
rect 6406 2719 6486 2730
rect 6538 2719 6618 2730
rect 6670 2719 6750 2730
rect 6802 2719 6882 2730
rect 6934 2719 7014 2730
rect 7066 2719 7146 2730
rect 7198 2719 7278 2730
rect 7330 2719 7410 2730
rect 5878 2678 5880 2719
rect 5802 2673 5880 2678
rect 5926 2678 5958 2719
rect 6050 2678 6090 2719
rect 6174 2678 6222 2719
rect 6298 2678 6354 2719
rect 6422 2678 6486 2719
rect 6546 2678 6618 2719
rect 5926 2673 6004 2678
rect 6050 2673 6128 2678
rect 6174 2673 6252 2678
rect 6298 2673 6376 2678
rect 6422 2673 6500 2678
rect 6546 2673 6624 2678
rect 6670 2673 6748 2719
rect 6802 2678 6872 2719
rect 6934 2678 6996 2719
rect 7066 2678 7120 2719
rect 7198 2678 7244 2719
rect 7330 2678 7368 2719
rect 7462 2678 7542 2730
rect 7594 2678 7606 2730
rect 6794 2673 6872 2678
rect 6918 2673 6996 2678
rect 7042 2673 7120 2678
rect 7166 2673 7244 2678
rect 7290 2673 7368 2678
rect 7414 2673 7606 2678
rect 2514 2598 7606 2673
rect 2514 2546 2526 2598
rect 2578 2546 2658 2598
rect 2710 2546 2790 2598
rect 2842 2546 2922 2598
rect 2974 2546 3054 2598
rect 3106 2546 3186 2598
rect 3238 2546 3318 2598
rect 3370 2546 3450 2598
rect 3502 2546 3582 2598
rect 3634 2546 3714 2598
rect 3766 2595 3846 2598
rect 3898 2595 3978 2598
rect 4030 2595 4110 2598
rect 4162 2595 4242 2598
rect 4294 2595 4374 2598
rect 4426 2595 4506 2598
rect 4558 2595 4638 2598
rect 4690 2595 4770 2598
rect 4822 2595 4902 2598
rect 4954 2595 5034 2598
rect 5086 2595 5166 2598
rect 5218 2595 5298 2598
rect 5350 2595 5430 2598
rect 3766 2549 3772 2595
rect 3818 2549 3846 2595
rect 3942 2549 3978 2595
rect 4066 2549 4110 2595
rect 4190 2549 4242 2595
rect 4314 2549 4374 2595
rect 4438 2549 4506 2595
rect 4562 2549 4638 2595
rect 4690 2549 4764 2595
rect 4822 2549 4888 2595
rect 4954 2549 5012 2595
rect 5086 2549 5136 2595
rect 5218 2549 5260 2595
rect 5350 2549 5384 2595
rect 3766 2546 3846 2549
rect 3898 2546 3978 2549
rect 4030 2546 4110 2549
rect 4162 2546 4242 2549
rect 4294 2546 4374 2549
rect 4426 2546 4506 2549
rect 4558 2546 4638 2549
rect 4690 2546 4770 2549
rect 4822 2546 4902 2549
rect 4954 2546 5034 2549
rect 5086 2546 5166 2549
rect 5218 2546 5298 2549
rect 5350 2546 5430 2549
rect 5482 2595 5562 2598
rect 5482 2549 5508 2595
rect 5554 2549 5562 2595
rect 5482 2546 5562 2549
rect 5614 2595 5694 2598
rect 5614 2549 5632 2595
rect 5678 2549 5694 2595
rect 5614 2546 5694 2549
rect 5746 2595 5826 2598
rect 5746 2549 5756 2595
rect 5802 2549 5826 2595
rect 5746 2546 5826 2549
rect 5878 2595 5958 2598
rect 6010 2595 6090 2598
rect 6142 2595 6222 2598
rect 6274 2595 6354 2598
rect 6406 2595 6486 2598
rect 6538 2595 6618 2598
rect 6670 2595 6750 2598
rect 6802 2595 6882 2598
rect 6934 2595 7014 2598
rect 7066 2595 7146 2598
rect 7198 2595 7278 2598
rect 7330 2595 7410 2598
rect 5878 2549 5880 2595
rect 5926 2549 5958 2595
rect 6050 2549 6090 2595
rect 6174 2549 6222 2595
rect 6298 2549 6354 2595
rect 6422 2549 6486 2595
rect 6546 2549 6618 2595
rect 6670 2549 6748 2595
rect 6802 2549 6872 2595
rect 6934 2549 6996 2595
rect 7066 2549 7120 2595
rect 7198 2549 7244 2595
rect 7330 2549 7368 2595
rect 5878 2546 5958 2549
rect 6010 2546 6090 2549
rect 6142 2546 6222 2549
rect 6274 2546 6354 2549
rect 6406 2546 6486 2549
rect 6538 2546 6618 2549
rect 6670 2546 6750 2549
rect 6802 2546 6882 2549
rect 6934 2546 7014 2549
rect 7066 2546 7146 2549
rect 7198 2546 7278 2549
rect 7330 2546 7410 2549
rect 7462 2546 7542 2598
rect 7594 2546 7606 2598
rect 2514 2471 7606 2546
rect 8004 2699 8036 3063
rect 8088 2699 8120 3063
rect 8004 2678 8120 2699
rect 8004 2632 8039 2678
rect 8085 2632 8120 2678
rect 8004 2565 8120 2632
rect 8004 2543 8039 2565
rect 8085 2543 8120 2565
rect 8263 3247 8309 3802
rect 8878 4265 9454 4299
rect 8878 4230 8981 4265
rect 8878 4184 8926 4230
rect 8972 4213 8981 4230
rect 9033 4230 9193 4265
rect 9033 4213 9084 4230
rect 8972 4184 9084 4213
rect 9130 4213 9193 4230
rect 9245 4249 9454 4265
rect 9245 4213 9451 4249
rect 9506 4247 9545 4299
rect 9130 4203 9451 4213
rect 9497 4203 9545 4247
rect 9130 4184 9545 4203
rect 8878 4081 9545 4184
rect 8878 4067 9451 4081
rect 8878 4021 8926 4067
rect 8972 4047 9084 4067
rect 8972 4021 8981 4047
rect 8878 3995 8981 4021
rect 9033 4021 9084 4047
rect 9130 4047 9451 4067
rect 9130 4021 9193 4047
rect 9033 3995 9193 4021
rect 9245 4035 9451 4047
rect 9245 4029 9454 4035
rect 9506 4029 9545 4081
rect 9245 3995 9545 4029
rect 8878 3913 9545 3995
rect 8878 3904 9451 3913
rect 8878 3858 8926 3904
rect 8972 3858 9084 3904
rect 9130 3867 9451 3904
rect 9497 3867 9545 3913
rect 9130 3864 9545 3867
rect 9130 3858 9454 3864
rect 8878 3812 9454 3858
rect 9506 3812 9545 3864
rect 8878 3746 9545 3812
rect 8878 3741 9451 3746
rect 8878 3695 8926 3741
rect 8972 3695 9084 3741
rect 9130 3700 9451 3741
rect 9497 3700 9545 3746
rect 9130 3695 9545 3700
rect 8878 3646 9545 3695
rect 8878 3594 9454 3646
rect 9506 3594 9545 3646
rect 8878 3578 9545 3594
rect 8878 3577 9451 3578
rect 8878 3531 8926 3577
rect 8972 3531 9084 3577
rect 9130 3532 9451 3577
rect 9497 3532 9545 3578
rect 9130 3531 9545 3532
rect 8878 3429 9545 3531
rect 8878 3414 9454 3429
rect 8878 3368 8926 3414
rect 8972 3368 9084 3414
rect 9130 3410 9454 3414
rect 9130 3368 9451 3410
rect 9506 3377 9545 3429
rect 8878 3364 9451 3368
rect 9497 3364 9545 3377
rect 8263 3133 8309 3201
rect 8263 3019 8309 3087
rect 8263 2905 8309 2973
rect 8263 2791 8309 2859
rect 8263 2678 8309 2745
rect 8263 2565 8309 2632
rect 8039 2506 8085 2519
rect 8452 3247 8568 3260
rect 8452 3201 8487 3247
rect 8533 3201 8568 3247
rect 8452 3133 8568 3201
rect 8452 3087 8487 3133
rect 8533 3087 8568 3133
rect 8452 3063 8568 3087
rect 8452 2699 8484 3063
rect 8536 2699 8568 3063
rect 8452 2678 8568 2699
rect 8452 2632 8487 2678
rect 8533 2632 8568 2678
rect 8452 2565 8568 2632
rect 8452 2543 8487 2565
rect 8263 2506 8309 2519
rect 8533 2543 8568 2565
rect 8878 3251 9545 3364
rect 8878 3205 8926 3251
rect 8972 3205 9084 3251
rect 9130 3242 9545 3251
rect 9130 3205 9451 3242
rect 9497 3211 9545 3242
rect 8878 3196 9451 3205
rect 8878 3159 9454 3196
rect 9506 3159 9545 3211
rect 8878 3088 9545 3159
rect 8878 3042 8926 3088
rect 8972 3042 9084 3088
rect 9130 3075 9545 3088
rect 9130 3042 9451 3075
rect 8878 3029 9451 3042
rect 9497 3029 9545 3075
rect 8878 2993 9545 3029
rect 8878 2941 9454 2993
rect 9506 2941 9545 2993
rect 8878 2925 9545 2941
rect 8878 2879 8926 2925
rect 8972 2879 9084 2925
rect 9130 2905 9545 2925
rect 9130 2879 9451 2905
rect 8878 2859 9451 2879
rect 9497 2859 9545 2905
rect 8878 2776 9545 2859
rect 8878 2761 9454 2776
rect 8878 2715 8926 2761
rect 8972 2715 9084 2761
rect 9130 2735 9454 2761
rect 9130 2715 9451 2735
rect 9506 2724 9545 2776
rect 8878 2689 9451 2715
rect 9497 2689 9545 2724
rect 8878 2598 9545 2689
rect 8878 2552 8926 2598
rect 8972 2552 9084 2598
rect 9130 2565 9545 2598
rect 9130 2552 9451 2565
rect 9497 2558 9545 2565
rect 8487 2506 8533 2519
rect 8878 2519 9451 2552
rect 8878 2506 9454 2519
rect 9506 2506 9545 2558
rect 2514 2466 3772 2471
rect 2514 2414 2526 2466
rect 2578 2414 2658 2466
rect 2710 2414 2790 2466
rect 2842 2414 2922 2466
rect 2974 2414 3054 2466
rect 3106 2414 3186 2466
rect 3238 2414 3318 2466
rect 3370 2414 3450 2466
rect 3502 2414 3582 2466
rect 3634 2414 3714 2466
rect 3766 2425 3772 2466
rect 3818 2466 3896 2471
rect 3942 2466 4020 2471
rect 4066 2466 4144 2471
rect 4190 2466 4268 2471
rect 4314 2466 4392 2471
rect 4438 2466 4516 2471
rect 4562 2466 4640 2471
rect 4686 2466 4764 2471
rect 4810 2466 4888 2471
rect 4934 2466 5012 2471
rect 5058 2466 5136 2471
rect 5182 2466 5260 2471
rect 5306 2466 5384 2471
rect 3818 2425 3846 2466
rect 3942 2425 3978 2466
rect 4066 2425 4110 2466
rect 4190 2425 4242 2466
rect 4314 2425 4374 2466
rect 4438 2425 4506 2466
rect 4562 2425 4638 2466
rect 4690 2425 4764 2466
rect 4822 2425 4888 2466
rect 4954 2425 5012 2466
rect 5086 2425 5136 2466
rect 5218 2425 5260 2466
rect 5350 2425 5384 2466
rect 5430 2466 5508 2471
rect 3766 2414 3846 2425
rect 3898 2414 3978 2425
rect 4030 2414 4110 2425
rect 4162 2414 4242 2425
rect 4294 2414 4374 2425
rect 4426 2414 4506 2425
rect 4558 2414 4638 2425
rect 4690 2414 4770 2425
rect 4822 2414 4902 2425
rect 4954 2414 5034 2425
rect 5086 2414 5166 2425
rect 5218 2414 5298 2425
rect 5350 2414 5430 2425
rect 5482 2425 5508 2466
rect 5554 2466 5632 2471
rect 5554 2425 5562 2466
rect 5482 2414 5562 2425
rect 5614 2425 5632 2466
rect 5678 2466 5756 2471
rect 5678 2425 5694 2466
rect 5614 2414 5694 2425
rect 5746 2425 5756 2466
rect 5802 2466 5880 2471
rect 5802 2425 5826 2466
rect 5746 2414 5826 2425
rect 5878 2425 5880 2466
rect 5926 2466 6004 2471
rect 6050 2466 6128 2471
rect 6174 2466 6252 2471
rect 6298 2466 6376 2471
rect 6422 2466 6500 2471
rect 6546 2466 6624 2471
rect 5926 2425 5958 2466
rect 6050 2425 6090 2466
rect 6174 2425 6222 2466
rect 6298 2425 6354 2466
rect 6422 2425 6486 2466
rect 6546 2425 6618 2466
rect 6670 2425 6748 2471
rect 6794 2466 6872 2471
rect 6918 2466 6996 2471
rect 7042 2466 7120 2471
rect 7166 2466 7244 2471
rect 7290 2466 7368 2471
rect 7414 2466 7606 2471
rect 6802 2425 6872 2466
rect 6934 2425 6996 2466
rect 7066 2425 7120 2466
rect 7198 2425 7244 2466
rect 7330 2425 7368 2466
rect 5878 2414 5958 2425
rect 6010 2414 6090 2425
rect 6142 2414 6222 2425
rect 6274 2414 6354 2425
rect 6406 2414 6486 2425
rect 6538 2414 6618 2425
rect 6670 2414 6750 2425
rect 6802 2414 6882 2425
rect 6934 2414 7014 2425
rect 7066 2414 7146 2425
rect 7198 2414 7278 2425
rect 7330 2414 7410 2425
rect 7462 2414 7542 2466
rect 7594 2414 7606 2466
rect 2514 2347 7606 2414
rect 2514 2334 3772 2347
rect 2514 2282 2526 2334
rect 2578 2282 2658 2334
rect 2710 2282 2790 2334
rect 2842 2282 2922 2334
rect 2974 2282 3054 2334
rect 3106 2282 3186 2334
rect 3238 2282 3318 2334
rect 3370 2282 3450 2334
rect 3502 2282 3582 2334
rect 3634 2282 3714 2334
rect 3766 2301 3772 2334
rect 3818 2334 3896 2347
rect 3942 2334 4020 2347
rect 4066 2334 4144 2347
rect 4190 2334 4268 2347
rect 4314 2334 4392 2347
rect 4438 2334 4516 2347
rect 4562 2334 4640 2347
rect 4686 2334 4764 2347
rect 4810 2334 4888 2347
rect 4934 2334 5012 2347
rect 5058 2334 5136 2347
rect 5182 2334 5260 2347
rect 5306 2334 5384 2347
rect 3818 2301 3846 2334
rect 3942 2301 3978 2334
rect 4066 2301 4110 2334
rect 4190 2301 4242 2334
rect 4314 2301 4374 2334
rect 4438 2301 4506 2334
rect 4562 2301 4638 2334
rect 4690 2301 4764 2334
rect 4822 2301 4888 2334
rect 4954 2301 5012 2334
rect 5086 2301 5136 2334
rect 5218 2301 5260 2334
rect 5350 2301 5384 2334
rect 5430 2334 5508 2347
rect 3766 2282 3846 2301
rect 3898 2282 3978 2301
rect 4030 2282 4110 2301
rect 4162 2282 4242 2301
rect 4294 2282 4374 2301
rect 4426 2282 4506 2301
rect 4558 2282 4638 2301
rect 4690 2282 4770 2301
rect 4822 2282 4902 2301
rect 4954 2282 5034 2301
rect 5086 2282 5166 2301
rect 5218 2282 5298 2301
rect 5350 2282 5430 2301
rect 5482 2301 5508 2334
rect 5554 2334 5632 2347
rect 5554 2301 5562 2334
rect 5482 2282 5562 2301
rect 5614 2301 5632 2334
rect 5678 2334 5756 2347
rect 5678 2301 5694 2334
rect 5614 2282 5694 2301
rect 5746 2301 5756 2334
rect 5802 2334 5880 2347
rect 5802 2301 5826 2334
rect 5746 2282 5826 2301
rect 5878 2301 5880 2334
rect 5926 2334 6004 2347
rect 6050 2334 6128 2347
rect 6174 2334 6252 2347
rect 6298 2334 6376 2347
rect 6422 2334 6500 2347
rect 6546 2334 6624 2347
rect 5926 2301 5958 2334
rect 6050 2301 6090 2334
rect 6174 2301 6222 2334
rect 6298 2301 6354 2334
rect 6422 2301 6486 2334
rect 6546 2301 6618 2334
rect 6670 2301 6748 2347
rect 6794 2334 6872 2347
rect 6918 2334 6996 2347
rect 7042 2334 7120 2347
rect 7166 2334 7244 2347
rect 7290 2334 7368 2347
rect 7414 2334 7606 2347
rect 6802 2301 6872 2334
rect 6934 2301 6996 2334
rect 7066 2301 7120 2334
rect 7198 2301 7244 2334
rect 7330 2301 7368 2334
rect 5878 2282 5958 2301
rect 6010 2282 6090 2301
rect 6142 2282 6222 2301
rect 6274 2282 6354 2301
rect 6406 2282 6486 2301
rect 6538 2282 6618 2301
rect 6670 2282 6750 2301
rect 6802 2282 6882 2301
rect 6934 2282 7014 2301
rect 7066 2282 7146 2301
rect 7198 2282 7278 2301
rect 7330 2282 7410 2301
rect 7462 2282 7542 2334
rect 7594 2282 7606 2334
rect 2514 2270 7606 2282
rect 8878 2435 9545 2506
rect 8878 2389 8926 2435
rect 8972 2389 9084 2435
rect 9130 2395 9545 2435
rect 9130 2389 9451 2395
rect 8878 2349 9451 2389
rect 9497 2349 9545 2395
rect 8878 2340 9545 2349
rect 8878 2288 9454 2340
rect 9506 2288 9545 2340
rect 8878 2271 9545 2288
rect 8878 2225 8926 2271
rect 8972 2225 9084 2271
rect 9130 2225 9545 2271
rect 8878 2179 9451 2225
rect 9497 2179 9545 2225
rect 8878 2123 9545 2179
rect 8878 2108 9454 2123
rect 8878 2062 8926 2108
rect 8972 2062 9084 2108
rect 9130 2071 9454 2108
rect 9506 2071 9545 2123
rect 9130 2062 9545 2071
rect 8878 2055 9545 2062
rect 8878 2009 9451 2055
rect 9497 2009 9545 2055
rect 8878 1945 9545 2009
rect 8878 1899 8926 1945
rect 8972 1899 9084 1945
rect 9130 1905 9545 1945
rect 9130 1899 9454 1905
rect 8878 1884 9454 1899
rect 8878 1838 9451 1884
rect 9506 1853 9545 1905
rect 9497 1838 9545 1853
rect 8878 1781 9545 1838
rect 8878 1735 8926 1781
rect 8972 1735 9084 1781
rect 9130 1735 9545 1781
rect 8878 1714 9545 1735
rect 8878 1668 9451 1714
rect 9497 1687 9545 1714
rect 8878 1635 9454 1668
rect 9506 1635 9545 1687
rect 8878 1618 9545 1635
rect 8878 1572 8926 1618
rect 8972 1572 9084 1618
rect 9130 1572 9545 1618
rect 8878 1544 9545 1572
rect 8878 1498 9451 1544
rect 9497 1498 9545 1544
rect 8878 1470 9545 1498
rect 8878 1455 9454 1470
rect 8878 1409 8926 1455
rect 8972 1409 9084 1455
rect 9130 1418 9454 1455
rect 9506 1418 9545 1470
rect 9130 1409 9545 1418
rect 8878 1374 9545 1409
rect 8878 1328 9451 1374
rect 9497 1328 9545 1374
rect 8878 1292 9545 1328
rect 8878 1246 8926 1292
rect 8972 1246 9084 1292
rect 9130 1252 9545 1292
rect 9130 1246 9454 1252
rect 8878 1204 9454 1246
rect 8878 1158 9451 1204
rect 9506 1200 9545 1252
rect 9497 1158 9545 1200
rect 8878 1129 9545 1158
rect 8878 1083 8926 1129
rect 8972 1083 9084 1129
rect 9130 1083 9545 1129
rect 8878 1035 9545 1083
rect 8878 1034 9454 1035
rect 8878 988 9451 1034
rect 8878 983 9454 988
rect 9506 983 9545 1035
rect 8878 965 9545 983
rect 8878 919 8926 965
rect 8972 919 9084 965
rect 9130 919 9545 965
rect 8878 864 9545 919
rect 8878 818 9451 864
rect 9497 818 9545 864
rect 8878 817 9545 818
rect 8878 802 9454 817
rect 8878 756 8926 802
rect 8972 756 9084 802
rect 9130 765 9454 802
rect 9506 765 9545 817
rect 9130 756 9545 765
rect 8878 694 9545 756
rect 8878 648 9451 694
rect 9497 648 9545 694
rect 8878 639 9545 648
rect 8878 593 8926 639
rect 8972 593 9084 639
rect 9130 599 9545 639
rect 9130 593 9454 599
rect 8878 547 9454 593
rect 9506 547 9545 599
rect 8878 524 9545 547
rect 8878 478 9451 524
rect 9497 478 9545 524
rect 8878 476 9545 478
rect 8878 430 8926 476
rect 8972 430 9084 476
rect 9130 430 9545 476
rect 8878 382 9545 430
rect 8878 354 9454 382
rect 8878 312 9451 354
rect 9506 330 9545 382
rect 8878 266 8926 312
rect 8972 266 9084 312
rect 9130 308 9451 312
rect 9497 308 9545 330
rect 9130 289 9545 308
rect 10088 4584 10300 4696
rect 10696 4869 10738 4909
rect 10650 4659 10696 4672
rect 10920 6335 10961 6376
rect 11056 8392 11095 8444
rect 11147 8392 11186 8444
rect 11056 8226 11098 8392
rect 11144 8226 11186 8392
rect 11056 8174 11095 8226
rect 11147 8174 11186 8226
rect 11056 8008 11098 8174
rect 11144 8008 11186 8174
rect 11056 7956 11095 8008
rect 11147 7956 11186 8008
rect 11056 7791 11098 7956
rect 11144 7791 11186 7956
rect 11056 7739 11095 7791
rect 11147 7739 11186 7791
rect 11056 7573 11098 7739
rect 11144 7573 11186 7739
rect 11056 7521 11095 7573
rect 11147 7521 11186 7573
rect 11056 7356 11098 7521
rect 11144 7356 11186 7521
rect 11056 7304 11095 7356
rect 11147 7304 11186 7356
rect 11056 7138 11098 7304
rect 11144 7138 11186 7304
rect 11056 7086 11095 7138
rect 11147 7086 11186 7138
rect 11056 6920 11098 7086
rect 11144 6920 11186 7086
rect 11056 6868 11095 6920
rect 11147 6868 11186 6920
rect 11056 6702 11098 6868
rect 11144 6702 11186 6868
rect 11056 6650 11095 6702
rect 11147 6650 11186 6702
rect 11056 6485 11098 6650
rect 11144 6485 11186 6650
rect 11056 6433 11095 6485
rect 11147 6433 11186 6485
rect 11056 6267 11098 6433
rect 11144 6267 11186 6433
rect 11281 8386 11322 8427
rect 11368 9126 11403 9182
rect 11546 9182 11592 9195
rect 11504 9097 11546 9137
rect 11935 9182 11981 9195
rect 11592 9097 11634 9137
rect 11504 9045 11543 9097
rect 11595 9045 11634 9097
rect 11504 8879 11546 9045
rect 11592 8879 11634 9045
rect 11504 8827 11543 8879
rect 11595 8827 11634 8879
rect 11504 8661 11546 8827
rect 11592 8661 11634 8827
rect 11504 8609 11543 8661
rect 11595 8609 11634 8661
rect 11504 8444 11546 8609
rect 11592 8444 11634 8609
rect 11368 8426 11400 8427
rect 11368 8386 11409 8426
rect 11281 8334 11319 8386
rect 11371 8334 11409 8386
rect 11281 8169 11322 8334
rect 11368 8169 11409 8334
rect 11281 8117 11319 8169
rect 11371 8117 11409 8169
rect 11281 7951 11322 8117
rect 11368 7951 11409 8117
rect 11281 7899 11319 7951
rect 11371 7899 11409 7951
rect 11281 7734 11322 7899
rect 11368 7734 11409 7899
rect 11281 7682 11319 7734
rect 11371 7682 11409 7734
rect 11281 7516 11322 7682
rect 11368 7516 11409 7682
rect 11281 7464 11319 7516
rect 11371 7464 11409 7516
rect 11281 7298 11322 7464
rect 11368 7298 11409 7464
rect 11281 7246 11319 7298
rect 11371 7246 11409 7298
rect 11281 7080 11322 7246
rect 11368 7080 11409 7246
rect 11281 7028 11319 7080
rect 11371 7028 11409 7080
rect 11281 6863 11322 7028
rect 11368 6863 11409 7028
rect 11281 6811 11319 6863
rect 11371 6811 11409 6863
rect 11281 6645 11322 6811
rect 11368 6645 11409 6811
rect 11281 6593 11319 6645
rect 11371 6593 11409 6645
rect 11281 6428 11322 6593
rect 11368 6428 11409 6593
rect 11281 6376 11319 6428
rect 11371 6376 11409 6428
rect 11281 6335 11322 6376
rect 11056 6215 11095 6267
rect 11147 6215 11186 6267
rect 11056 6050 11098 6215
rect 11144 6050 11186 6215
rect 11056 5998 11095 6050
rect 11147 5998 11186 6050
rect 11056 5832 11098 5998
rect 11144 5832 11186 5998
rect 11056 5780 11095 5832
rect 11147 5780 11186 5832
rect 11056 5614 11098 5780
rect 11144 5614 11186 5780
rect 11056 5562 11095 5614
rect 11147 5562 11186 5614
rect 11056 5397 11098 5562
rect 11144 5397 11186 5562
rect 11056 5345 11095 5397
rect 11147 5345 11186 5397
rect 11056 5179 11098 5345
rect 11144 5179 11186 5345
rect 11056 5127 11095 5179
rect 11147 5127 11186 5179
rect 11056 4961 11098 5127
rect 11144 4961 11186 5127
rect 11056 4909 11095 4961
rect 11147 4909 11186 4961
rect 11056 4869 11098 4909
rect 10874 4659 10920 4672
rect 11144 4869 11186 4909
rect 11098 4659 11144 4672
rect 11368 6335 11409 6376
rect 11504 8392 11543 8444
rect 11595 8392 11634 8444
rect 11504 8226 11546 8392
rect 11592 8226 11634 8392
rect 11504 8174 11543 8226
rect 11595 8174 11634 8226
rect 11504 8008 11546 8174
rect 11592 8008 11634 8174
rect 11504 7956 11543 8008
rect 11595 7956 11634 8008
rect 11504 7791 11546 7956
rect 11592 7791 11634 7956
rect 11504 7739 11543 7791
rect 11595 7739 11634 7791
rect 11504 7573 11546 7739
rect 11592 7573 11634 7739
rect 11504 7521 11543 7573
rect 11595 7521 11634 7573
rect 11504 7356 11546 7521
rect 11592 7356 11634 7521
rect 11504 7304 11543 7356
rect 11595 7304 11634 7356
rect 11504 7138 11546 7304
rect 11592 7138 11634 7304
rect 11504 7086 11543 7138
rect 11595 7086 11634 7138
rect 11504 6920 11546 7086
rect 11592 6920 11634 7086
rect 11504 6868 11543 6920
rect 11595 6868 11634 6920
rect 11504 6702 11546 6868
rect 11592 6702 11634 6868
rect 11504 6650 11543 6702
rect 11595 6650 11634 6702
rect 11504 6485 11546 6650
rect 11592 6485 11634 6650
rect 11504 6433 11543 6485
rect 11595 6433 11634 6485
rect 11504 6267 11546 6433
rect 11592 6267 11634 6433
rect 11504 6215 11543 6267
rect 11595 6215 11634 6267
rect 11504 6050 11546 6215
rect 11592 6050 11634 6215
rect 11504 5998 11543 6050
rect 11595 5998 11634 6050
rect 11504 5832 11546 5998
rect 11592 5832 11634 5998
rect 11504 5780 11543 5832
rect 11595 5780 11634 5832
rect 11504 5614 11546 5780
rect 11592 5614 11634 5780
rect 11504 5562 11543 5614
rect 11595 5562 11634 5614
rect 11504 5397 11546 5562
rect 11592 5397 11634 5562
rect 11504 5345 11543 5397
rect 11595 5345 11634 5397
rect 11504 5179 11546 5345
rect 11592 5179 11634 5345
rect 11504 5127 11543 5179
rect 11595 5127 11634 5179
rect 11504 4961 11546 5127
rect 11592 4961 11634 5127
rect 11504 4909 11543 4961
rect 11595 4909 11634 4961
rect 11504 4869 11546 4909
rect 11322 4659 11368 4672
rect 11592 4869 11634 4909
rect 11893 5413 11935 5453
rect 12124 9182 12239 9412
rect 12124 9126 12159 9182
rect 12115 8400 12159 8441
rect 12205 9126 12239 9182
rect 12383 9182 12429 9195
rect 12205 8440 12234 8441
rect 12115 8348 12153 8400
rect 12115 8183 12159 8348
rect 12115 8131 12153 8183
rect 12115 7965 12159 8131
rect 12115 7913 12153 7965
rect 12115 7748 12159 7913
rect 12115 7696 12153 7748
rect 12115 7530 12159 7696
rect 12115 7478 12153 7530
rect 12115 7312 12159 7478
rect 12115 7260 12153 7312
rect 12115 7094 12159 7260
rect 12115 7042 12153 7094
rect 12115 6877 12159 7042
rect 12115 6825 12153 6877
rect 12115 6659 12159 6825
rect 12115 6607 12153 6659
rect 12115 6442 12159 6607
rect 12115 6390 12153 6442
rect 12115 6349 12159 6390
rect 11981 5413 12021 5453
rect 11893 5361 11931 5413
rect 11983 5361 12021 5413
rect 11893 5195 11935 5361
rect 11981 5195 12021 5361
rect 11893 5143 11931 5195
rect 11983 5143 12021 5195
rect 11893 4977 11935 5143
rect 11981 4977 12021 5143
rect 11893 4925 11931 4977
rect 11983 4925 12021 4977
rect 11546 4659 11592 4672
rect 11893 4759 11935 4925
rect 11981 4759 12021 4925
rect 11893 4707 11931 4759
rect 11983 4712 12021 4759
rect 11983 4707 12022 4712
rect 11893 4672 11935 4707
rect 11981 4672 12022 4707
rect 10088 4538 10123 4584
rect 10169 4538 10300 4584
rect 11893 4574 12022 4672
rect 12205 6349 12243 8440
rect 12159 4659 12205 4672
rect 12341 5413 12383 5453
rect 12571 9182 12687 9412
rect 13217 9332 13491 9412
rect 13217 9286 13252 9332
rect 13298 9286 13410 9332
rect 13456 9286 13491 9332
rect 12571 9126 12607 9182
rect 12563 8400 12607 8441
rect 12653 9126 12687 9182
rect 12831 9182 12877 9195
rect 12653 8440 12682 8441
rect 12563 8348 12601 8400
rect 12563 8183 12607 8348
rect 12563 8131 12601 8183
rect 12563 7965 12607 8131
rect 12563 7913 12601 7965
rect 12563 7748 12607 7913
rect 12563 7696 12601 7748
rect 12563 7530 12607 7696
rect 12563 7478 12601 7530
rect 12563 7312 12607 7478
rect 12563 7260 12601 7312
rect 12563 7094 12607 7260
rect 12563 7042 12601 7094
rect 12563 6877 12607 7042
rect 12563 6825 12601 6877
rect 12563 6659 12607 6825
rect 12563 6607 12601 6659
rect 12563 6442 12607 6607
rect 12563 6390 12601 6442
rect 12563 6349 12607 6390
rect 12429 5413 12469 5453
rect 12341 5361 12379 5413
rect 12431 5361 12469 5413
rect 12341 5195 12383 5361
rect 12429 5195 12469 5361
rect 12341 5143 12379 5195
rect 12431 5143 12469 5195
rect 12341 4977 12383 5143
rect 12429 4977 12469 5143
rect 12341 4925 12379 4977
rect 12431 4925 12469 4977
rect 12341 4759 12383 4925
rect 12429 4759 12469 4925
rect 12341 4707 12379 4759
rect 12431 4707 12469 4759
rect 12341 4672 12383 4707
rect 12429 4672 12469 4707
rect 12341 4667 12469 4672
rect 12653 6349 12691 8440
rect 12383 4659 12429 4667
rect 12607 4659 12653 4672
rect 12789 5413 12831 5453
rect 13217 9169 13491 9286
rect 13217 9123 13252 9169
rect 13298 9123 13410 9169
rect 13456 9123 13491 9169
rect 13217 9006 13491 9123
rect 13217 8960 13252 9006
rect 13298 8960 13410 9006
rect 13456 8960 13491 9006
rect 13217 8843 13491 8960
rect 13217 8797 13252 8843
rect 13298 8797 13410 8843
rect 13456 8797 13491 8843
rect 13217 8679 13491 8797
rect 13217 8633 13252 8679
rect 13298 8633 13410 8679
rect 13456 8633 13491 8679
rect 13217 8516 13491 8633
rect 13217 8470 13252 8516
rect 13298 8470 13410 8516
rect 13456 8470 13491 8516
rect 13217 8400 13491 8470
rect 13217 8353 13400 8400
rect 13452 8353 13491 8400
rect 13217 8307 13252 8353
rect 13298 8348 13400 8353
rect 13298 8307 13410 8348
rect 13456 8307 13491 8353
rect 13217 8190 13491 8307
rect 13217 8144 13252 8190
rect 13298 8183 13410 8190
rect 13298 8144 13400 8183
rect 13456 8144 13491 8190
rect 13217 8131 13400 8144
rect 13452 8131 13491 8144
rect 13217 8026 13491 8131
rect 13217 7980 13252 8026
rect 13298 7980 13410 8026
rect 13456 7980 13491 8026
rect 13217 7965 13491 7980
rect 13217 7913 13400 7965
rect 13452 7913 13491 7965
rect 13217 7863 13491 7913
rect 13217 7817 13252 7863
rect 13298 7817 13410 7863
rect 13456 7817 13491 7863
rect 13217 7748 13491 7817
rect 13217 7700 13400 7748
rect 13452 7700 13491 7748
rect 13217 7654 13252 7700
rect 13298 7696 13400 7700
rect 13298 7654 13410 7696
rect 13456 7654 13491 7700
rect 13217 7537 13491 7654
rect 13217 7491 13252 7537
rect 13298 7530 13410 7537
rect 13298 7491 13400 7530
rect 13456 7491 13491 7537
rect 13217 7478 13400 7491
rect 13452 7478 13491 7491
rect 13217 7373 13491 7478
rect 13217 7327 13252 7373
rect 13298 7327 13410 7373
rect 13456 7327 13491 7373
rect 13217 7312 13491 7327
rect 13217 7260 13400 7312
rect 13452 7260 13491 7312
rect 13217 7210 13491 7260
rect 13217 7164 13252 7210
rect 13298 7164 13410 7210
rect 13456 7164 13491 7210
rect 13217 7094 13491 7164
rect 13217 7047 13400 7094
rect 13452 7047 13491 7094
rect 13217 7001 13252 7047
rect 13298 7042 13400 7047
rect 13298 7001 13410 7042
rect 13456 7001 13491 7047
rect 13217 6883 13491 7001
rect 13217 6837 13252 6883
rect 13298 6877 13410 6883
rect 13298 6837 13400 6877
rect 13456 6837 13491 6883
rect 13217 6825 13400 6837
rect 13452 6825 13491 6837
rect 13217 6720 13491 6825
rect 13217 6674 13252 6720
rect 13298 6674 13410 6720
rect 13456 6674 13491 6720
rect 13217 6659 13491 6674
rect 13217 6607 13400 6659
rect 13452 6607 13491 6659
rect 13217 6557 13491 6607
rect 13217 6511 13252 6557
rect 13298 6511 13410 6557
rect 13456 6511 13491 6557
rect 13217 6442 13491 6511
rect 13217 6394 13400 6442
rect 13452 6394 13491 6442
rect 13217 6348 13252 6394
rect 13298 6390 13400 6394
rect 13298 6348 13410 6390
rect 13456 6348 13491 6394
rect 13217 6230 13491 6348
rect 13217 6184 13252 6230
rect 13298 6184 13410 6230
rect 13456 6184 13491 6230
rect 13217 6067 13491 6184
rect 13217 6021 13252 6067
rect 13298 6021 13410 6067
rect 13456 6021 13491 6067
rect 13217 5904 13491 6021
rect 13217 5858 13252 5904
rect 13298 5858 13410 5904
rect 13456 5858 13491 5904
rect 13217 5741 13491 5858
rect 13217 5695 13252 5741
rect 13298 5695 13410 5741
rect 13456 5695 13491 5741
rect 13217 5577 13491 5695
rect 13217 5531 13252 5577
rect 13298 5531 13410 5577
rect 13456 5531 13491 5577
rect 12877 5413 12917 5453
rect 12789 5361 12827 5413
rect 12879 5361 12917 5413
rect 12789 5195 12831 5361
rect 12877 5195 12917 5361
rect 12789 5143 12827 5195
rect 12879 5143 12917 5195
rect 12789 4977 12831 5143
rect 12877 4977 12917 5143
rect 12789 4925 12827 4977
rect 12879 4925 12917 4977
rect 12789 4759 12831 4925
rect 12877 4759 12917 4925
rect 13217 5414 13491 5531
rect 13217 5368 13252 5414
rect 13298 5368 13410 5414
rect 13456 5368 13491 5414
rect 13217 5251 13491 5368
rect 13217 5205 13252 5251
rect 13298 5205 13410 5251
rect 13456 5205 13491 5251
rect 13217 5088 13491 5205
rect 13217 5042 13252 5088
rect 13298 5042 13410 5088
rect 13456 5042 13491 5088
rect 13217 4925 13491 5042
rect 13217 4879 13252 4925
rect 13298 4879 13410 4925
rect 13456 4879 13491 4925
rect 13217 4842 13491 4879
rect 12789 4707 12827 4759
rect 12879 4707 12917 4759
rect 12789 4672 12831 4707
rect 12877 4672 12917 4707
rect 12789 4667 12917 4672
rect 12831 4659 12877 4667
rect 10088 4417 10300 4538
rect 10727 4537 12022 4574
rect 12595 4540 12935 4553
rect 10727 4491 10763 4537
rect 10809 4491 11434 4537
rect 11480 4491 12022 4537
rect 10727 4454 12022 4491
rect 12268 4512 12935 4540
rect 12268 4506 12633 4512
rect 12268 4460 12294 4506
rect 12528 4460 12633 4506
rect 12685 4460 12845 4512
rect 12897 4460 12935 4512
rect 12268 4420 12935 4460
rect 10088 4371 10123 4417
rect 10169 4371 10300 4417
rect 10088 4356 10300 4371
rect 10088 4319 11258 4356
rect 10088 4273 11049 4319
rect 11189 4273 11258 4319
rect 10088 4249 11258 4273
rect 10088 4203 10123 4249
rect 10169 4236 11258 4249
rect 11557 4324 11897 4331
rect 11557 4290 12799 4324
rect 11557 4238 11595 4290
rect 11647 4238 11807 4290
rect 11859 4288 12799 4290
rect 11859 4242 12046 4288
rect 12092 4242 12718 4288
rect 12764 4242 12799 4288
rect 11859 4238 12799 4242
rect 10169 4203 10300 4236
rect 10088 4081 10300 4203
rect 11557 4204 12799 4238
rect 13305 4237 13605 4281
rect 11557 4198 11897 4204
rect 13305 4191 13353 4237
rect 13399 4191 13511 4237
rect 13557 4191 13605 4237
rect 13305 4104 13605 4191
rect 10088 4035 10123 4081
rect 10169 4035 10300 4081
rect 10088 3913 10300 4035
rect 10615 4068 10731 4104
rect 10615 4032 10650 4068
rect 10088 3867 10123 3913
rect 10169 3867 10300 3913
rect 10088 3746 10300 3867
rect 10088 3700 10123 3746
rect 10169 3700 10300 3746
rect 10088 3578 10300 3700
rect 10088 3532 10123 3578
rect 10169 3532 10300 3578
rect 10088 3410 10300 3532
rect 10088 3364 10123 3410
rect 10169 3364 10300 3410
rect 10088 3242 10300 3364
rect 10088 3196 10123 3242
rect 10169 3196 10300 3242
rect 10088 3075 10300 3196
rect 10088 3029 10123 3075
rect 10169 3029 10300 3075
rect 10088 2905 10300 3029
rect 10088 2859 10123 2905
rect 10169 2859 10300 2905
rect 10088 2735 10300 2859
rect 10088 2689 10123 2735
rect 10169 2689 10300 2735
rect 10088 2565 10300 2689
rect 10088 2519 10123 2565
rect 10169 2519 10300 2565
rect 10088 2395 10300 2519
rect 10088 2349 10123 2395
rect 10169 2349 10300 2395
rect 10088 2225 10300 2349
rect 10088 2179 10123 2225
rect 10169 2179 10300 2225
rect 10088 2055 10300 2179
rect 10088 2009 10123 2055
rect 10169 2009 10300 2055
rect 10088 1884 10300 2009
rect 10088 1838 10123 1884
rect 10169 1838 10300 1884
rect 10088 1714 10300 1838
rect 10088 1668 10123 1714
rect 10169 1668 10300 1714
rect 10088 1544 10300 1668
rect 10088 1498 10123 1544
rect 10169 1498 10300 1544
rect 10088 1374 10300 1498
rect 10088 1328 10123 1374
rect 10169 1328 10300 1374
rect 10088 1204 10300 1328
rect 10088 1158 10123 1204
rect 10169 1158 10300 1204
rect 10088 1034 10300 1158
rect 10088 988 10123 1034
rect 10169 988 10300 1034
rect 10088 864 10300 988
rect 10088 818 10123 864
rect 10169 818 10300 864
rect 10088 694 10300 818
rect 10088 648 10123 694
rect 10169 648 10300 694
rect 10088 524 10300 648
rect 10088 478 10123 524
rect 10169 478 10300 524
rect 10088 354 10300 478
rect 10088 308 10123 354
rect 10169 308 10300 354
rect 9130 266 9532 289
rect 10088 271 10300 308
rect 10609 4022 10650 4032
rect 10696 4032 10731 4068
rect 11057 4068 11186 4104
rect 11057 4064 11098 4068
rect 11144 4064 11186 4068
rect 10696 4022 10738 4032
rect 10609 3991 10738 4022
rect 10609 3939 10647 3991
rect 10699 3939 10738 3991
rect 10609 3900 10738 3939
rect 10609 3854 10650 3900
rect 10696 3854 10738 3900
rect 10609 3773 10738 3854
rect 10609 3721 10647 3773
rect 10699 3721 10738 3773
rect 10609 3686 10650 3721
rect 10696 3686 10738 3721
rect 10609 3564 10738 3686
rect 10609 3556 10650 3564
rect 10696 3556 10738 3564
rect 10609 3504 10647 3556
rect 10699 3504 10738 3556
rect 10609 3397 10738 3504
rect 10609 3351 10650 3397
rect 10696 3351 10738 3397
rect 10609 3338 10738 3351
rect 10609 3286 10647 3338
rect 10699 3286 10738 3338
rect 10609 3229 10738 3286
rect 10609 3183 10650 3229
rect 10696 3183 10738 3229
rect 10609 3120 10738 3183
rect 10609 3068 10647 3120
rect 10699 3068 10738 3120
rect 10609 3061 10738 3068
rect 10609 3015 10650 3061
rect 10696 3015 10738 3061
rect 10609 2903 10738 3015
rect 10609 2851 10647 2903
rect 10699 2851 10738 2903
rect 10609 2847 10650 2851
rect 10696 2847 10738 2851
rect 10609 2726 10738 2847
rect 10609 2685 10650 2726
rect 10696 2685 10738 2726
rect 10609 2633 10647 2685
rect 10699 2633 10738 2685
rect 10609 2558 10738 2633
rect 10609 2512 10650 2558
rect 10696 2512 10738 2558
rect 10609 2468 10738 2512
rect 10609 2416 10647 2468
rect 10699 2416 10738 2468
rect 10609 2390 10738 2416
rect 10609 2344 10650 2390
rect 10696 2344 10738 2390
rect 10609 2250 10738 2344
rect 10609 2198 10647 2250
rect 10699 2198 10738 2250
rect 11057 4012 11095 4064
rect 11147 4012 11186 4064
rect 11511 4068 11627 4104
rect 11511 4032 11546 4068
rect 11057 3900 11186 4012
rect 11057 3854 11098 3900
rect 11144 3854 11186 3900
rect 11057 3846 11186 3854
rect 11057 3794 11095 3846
rect 11147 3794 11186 3846
rect 11057 3732 11186 3794
rect 11057 3686 11098 3732
rect 11144 3686 11186 3732
rect 11057 3628 11186 3686
rect 11057 3576 11095 3628
rect 11147 3576 11186 3628
rect 11057 3564 11186 3576
rect 11057 3518 11098 3564
rect 11144 3518 11186 3564
rect 11057 3411 11186 3518
rect 11057 3359 11095 3411
rect 11147 3359 11186 3411
rect 11057 3351 11098 3359
rect 11144 3351 11186 3359
rect 11057 3229 11186 3351
rect 11057 3193 11098 3229
rect 11144 3193 11186 3229
rect 11057 3141 11095 3193
rect 11147 3141 11186 3193
rect 11057 3061 11186 3141
rect 11057 3015 11098 3061
rect 11144 3015 11186 3061
rect 11057 2975 11186 3015
rect 11057 2923 11095 2975
rect 11147 2923 11186 2975
rect 11057 2893 11186 2923
rect 11057 2847 11098 2893
rect 11144 2847 11186 2893
rect 11057 2758 11186 2847
rect 11057 2706 11095 2758
rect 11147 2706 11186 2758
rect 11057 2680 11098 2706
rect 11144 2680 11186 2706
rect 11057 2558 11186 2680
rect 11057 2540 11098 2558
rect 11144 2540 11186 2558
rect 11057 2488 11095 2540
rect 11147 2488 11186 2540
rect 11057 2390 11186 2488
rect 11057 2344 11098 2390
rect 11144 2344 11186 2390
rect 11057 2322 11186 2344
rect 11057 2270 11095 2322
rect 11147 2270 11186 2322
rect 11057 2230 11186 2270
rect 11505 4022 11546 4032
rect 11592 4032 11627 4068
rect 11900 4068 12015 4104
rect 11900 4032 11934 4068
rect 11592 4022 11634 4032
rect 11505 3991 11634 4022
rect 11505 3939 11543 3991
rect 11595 3939 11634 3991
rect 11505 3900 11634 3939
rect 11505 3854 11546 3900
rect 11592 3854 11634 3900
rect 11505 3773 11634 3854
rect 11505 3721 11543 3773
rect 11595 3721 11634 3773
rect 11505 3686 11546 3721
rect 11592 3686 11634 3721
rect 11505 3564 11634 3686
rect 11505 3556 11546 3564
rect 11592 3556 11634 3564
rect 11505 3504 11543 3556
rect 11595 3504 11634 3556
rect 11505 3397 11634 3504
rect 11505 3351 11546 3397
rect 11592 3351 11634 3397
rect 11505 3338 11634 3351
rect 11505 3286 11543 3338
rect 11595 3286 11634 3338
rect 11505 3229 11634 3286
rect 11505 3183 11546 3229
rect 11592 3183 11634 3229
rect 11505 3120 11634 3183
rect 11505 3068 11543 3120
rect 11595 3068 11634 3120
rect 11505 3061 11634 3068
rect 11505 3015 11546 3061
rect 11592 3015 11634 3061
rect 11505 2903 11634 3015
rect 11505 2851 11543 2903
rect 11595 2851 11634 2903
rect 11505 2847 11546 2851
rect 11592 2847 11634 2851
rect 11505 2726 11634 2847
rect 11505 2685 11546 2726
rect 11592 2685 11634 2726
rect 11505 2633 11543 2685
rect 11595 2633 11634 2685
rect 11505 2558 11634 2633
rect 11505 2512 11546 2558
rect 11592 2512 11634 2558
rect 11505 2468 11634 2512
rect 11505 2416 11543 2468
rect 11595 2416 11634 2468
rect 11505 2390 11634 2416
rect 11505 2344 11546 2390
rect 11592 2344 11634 2390
rect 11505 2250 11634 2344
rect 10609 2174 10650 2198
rect 10696 2174 10738 2198
rect 10609 2050 10738 2174
rect 10609 2032 10650 2050
rect 10696 2032 10738 2050
rect 10609 1980 10647 2032
rect 10699 1980 10738 2032
rect 10609 1880 10738 1980
rect 10609 1834 10650 1880
rect 10696 1834 10738 1880
rect 10609 1814 10738 1834
rect 10609 1762 10647 1814
rect 10699 1762 10738 1814
rect 10609 1710 10738 1762
rect 10609 1664 10650 1710
rect 10696 1664 10738 1710
rect 10609 1597 10738 1664
rect 10609 1545 10647 1597
rect 10699 1545 10738 1597
rect 10609 1540 10738 1545
rect 10609 1494 10650 1540
rect 10696 1494 10738 1540
rect 10609 1379 10738 1494
rect 10609 1327 10647 1379
rect 10699 1327 10738 1379
rect 10609 1324 10650 1327
rect 10696 1324 10738 1327
rect 10609 1200 10738 1324
rect 10609 1162 10650 1200
rect 10696 1162 10738 1200
rect 10609 1110 10647 1162
rect 10699 1110 10738 1162
rect 10609 1030 10738 1110
rect 10609 984 10650 1030
rect 10696 984 10738 1030
rect 10609 944 10738 984
rect 10609 892 10647 944
rect 10699 892 10738 944
rect 10609 860 10738 892
rect 10609 814 10650 860
rect 10696 814 10738 860
rect 10609 726 10738 814
rect 10609 674 10647 726
rect 10699 674 10738 726
rect 10609 644 10650 674
rect 10696 644 10738 674
rect 10609 509 10738 644
rect 10609 457 10647 509
rect 10699 457 10738 509
rect 11063 2220 11179 2230
rect 11063 2174 11098 2220
rect 11144 2174 11179 2220
rect 11063 2050 11179 2174
rect 11063 2004 11098 2050
rect 11144 2004 11179 2050
rect 11063 1880 11179 2004
rect 11063 1834 11098 1880
rect 11144 1834 11179 1880
rect 11063 1710 11179 1834
rect 11063 1664 11098 1710
rect 11144 1664 11179 1710
rect 11063 1540 11179 1664
rect 11063 1494 11098 1540
rect 11144 1494 11179 1540
rect 11063 1370 11179 1494
rect 11063 1324 11098 1370
rect 11144 1324 11179 1370
rect 11063 1200 11179 1324
rect 11063 1154 11098 1200
rect 11144 1154 11179 1200
rect 11063 1030 11179 1154
rect 11063 984 11098 1030
rect 11144 984 11179 1030
rect 11063 860 11179 984
rect 11063 814 11098 860
rect 11144 814 11179 860
rect 11063 690 11179 814
rect 11063 644 11098 690
rect 11144 644 11179 690
rect 11063 493 11179 644
rect 11505 2198 11543 2250
rect 11595 2198 11634 2250
rect 11505 2174 11546 2198
rect 11592 2174 11634 2198
rect 11505 2050 11634 2174
rect 11505 2032 11546 2050
rect 11592 2032 11634 2050
rect 11505 1980 11543 2032
rect 11595 1980 11634 2032
rect 11505 1880 11634 1980
rect 11505 1834 11546 1880
rect 11592 1834 11634 1880
rect 11505 1814 11634 1834
rect 11505 1762 11543 1814
rect 11595 1762 11634 1814
rect 11505 1710 11634 1762
rect 11505 1664 11546 1710
rect 11592 1664 11634 1710
rect 11505 1597 11634 1664
rect 11505 1545 11543 1597
rect 11595 1545 11634 1597
rect 11505 1540 11634 1545
rect 11505 1494 11546 1540
rect 11592 1494 11634 1540
rect 11505 1379 11634 1494
rect 11505 1327 11543 1379
rect 11595 1327 11634 1379
rect 11505 1324 11546 1327
rect 11592 1324 11634 1327
rect 11505 1200 11634 1324
rect 11505 1162 11546 1200
rect 11592 1162 11634 1200
rect 11505 1110 11543 1162
rect 11595 1110 11634 1162
rect 11505 1030 11634 1110
rect 11505 984 11546 1030
rect 11592 984 11634 1030
rect 11505 944 11634 984
rect 11505 892 11543 944
rect 11595 892 11634 944
rect 11505 860 11634 892
rect 11505 814 11546 860
rect 11592 814 11634 860
rect 11505 726 11634 814
rect 11505 674 11543 726
rect 11595 674 11634 726
rect 11505 644 11546 674
rect 11592 644 11634 674
rect 11505 509 11634 644
rect 10609 291 10738 457
rect 8878 149 9532 266
rect 10609 239 10647 291
rect 10699 239 10738 291
rect 10609 199 10738 239
rect 11505 457 11543 509
rect 11595 457 11634 509
rect 11505 291 11634 457
rect 11505 239 11543 291
rect 11595 239 11634 291
rect 11505 199 11634 239
rect 11893 4022 11934 4032
rect 11980 4032 12015 4068
rect 12341 4068 12470 4104
rect 12341 4064 12382 4068
rect 12428 4064 12470 4068
rect 11980 4022 12022 4032
rect 11893 3991 12022 4022
rect 11893 3939 11931 3991
rect 11983 3939 12022 3991
rect 11893 3900 12022 3939
rect 11893 3854 11934 3900
rect 11980 3854 12022 3900
rect 11893 3773 12022 3854
rect 11893 3721 11931 3773
rect 11983 3721 12022 3773
rect 11893 3686 11934 3721
rect 11980 3686 12022 3721
rect 11893 3564 12022 3686
rect 11893 3556 11934 3564
rect 11980 3556 12022 3564
rect 11893 3504 11931 3556
rect 11983 3504 12022 3556
rect 11893 3397 12022 3504
rect 11893 3351 11934 3397
rect 11980 3351 12022 3397
rect 11893 3338 12022 3351
rect 11893 3286 11931 3338
rect 11983 3286 12022 3338
rect 11893 3120 12022 3286
rect 11893 3068 11931 3120
rect 11983 3068 12022 3120
rect 11893 2903 12022 3068
rect 11893 2851 11931 2903
rect 11983 2851 12022 2903
rect 11893 2685 12022 2851
rect 11893 2633 11931 2685
rect 11983 2633 12022 2685
rect 11893 2468 12022 2633
rect 11893 2416 11931 2468
rect 11983 2416 12022 2468
rect 11893 2250 12022 2416
rect 11893 2198 11931 2250
rect 11983 2198 12022 2250
rect 12341 4012 12379 4064
rect 12431 4012 12470 4064
rect 12795 4074 13605 4104
rect 12795 4068 13353 4074
rect 12795 4032 12830 4068
rect 12341 3900 12470 4012
rect 12341 3854 12382 3900
rect 12428 3854 12470 3900
rect 12341 3846 12470 3854
rect 12341 3794 12379 3846
rect 12431 3794 12470 3846
rect 12341 3732 12470 3794
rect 12341 3686 12382 3732
rect 12428 3686 12470 3732
rect 12341 3628 12470 3686
rect 12341 3576 12379 3628
rect 12431 3576 12470 3628
rect 12341 3564 12470 3576
rect 12341 3518 12382 3564
rect 12428 3518 12470 3564
rect 12341 3411 12470 3518
rect 12341 3359 12379 3411
rect 12431 3359 12470 3411
rect 12341 3351 12382 3359
rect 12428 3351 12470 3359
rect 12341 3193 12470 3351
rect 12341 3141 12379 3193
rect 12431 3141 12470 3193
rect 12341 2975 12470 3141
rect 12341 2923 12379 2975
rect 12431 2923 12470 2975
rect 12341 2758 12470 2923
rect 12341 2706 12379 2758
rect 12431 2706 12470 2758
rect 12341 2540 12470 2706
rect 12341 2488 12379 2540
rect 12431 2488 12470 2540
rect 12341 2322 12470 2488
rect 12341 2270 12379 2322
rect 12431 2270 12470 2322
rect 12341 2230 12470 2270
rect 12789 4022 12830 4032
rect 12876 4028 13353 4068
rect 13399 4028 13511 4074
rect 13557 4032 13605 4074
rect 13557 4028 13606 4032
rect 12876 4022 13606 4028
rect 12789 3991 13606 4022
rect 12789 3939 12827 3991
rect 12879 3939 13515 3991
rect 13567 3939 13606 3991
rect 12789 3905 13606 3939
rect 12789 3859 13353 3905
rect 13399 3859 13511 3905
rect 13557 3859 13606 3905
rect 12789 3773 13606 3859
rect 12789 3721 12827 3773
rect 12879 3742 13515 3773
rect 12879 3721 13353 3742
rect 12789 3686 12830 3721
rect 12876 3696 13353 3721
rect 13399 3696 13511 3742
rect 13567 3721 13606 3773
rect 13557 3696 13606 3721
rect 12876 3686 13606 3696
rect 12789 3578 13606 3686
rect 12789 3564 13353 3578
rect 12789 3556 12830 3564
rect 12876 3556 13353 3564
rect 12789 3504 12827 3556
rect 12879 3532 13353 3556
rect 13399 3532 13511 3578
rect 13557 3556 13606 3578
rect 12879 3504 13515 3532
rect 13567 3504 13606 3556
rect 12789 3415 13606 3504
rect 12789 3397 13353 3415
rect 12789 3351 12830 3397
rect 12876 3369 13353 3397
rect 13399 3369 13511 3415
rect 13557 3369 13606 3415
rect 12876 3351 13606 3369
rect 12789 3338 13606 3351
rect 12789 3286 12827 3338
rect 12879 3286 13515 3338
rect 13567 3286 13606 3338
rect 12789 3252 13606 3286
rect 12789 3206 13353 3252
rect 13399 3206 13511 3252
rect 13557 3206 13606 3252
rect 12789 3120 13606 3206
rect 12789 3068 12827 3120
rect 12879 3089 13515 3120
rect 12879 3068 13353 3089
rect 12789 3043 13353 3068
rect 13399 3043 13511 3089
rect 13567 3068 13606 3120
rect 13557 3043 13606 3068
rect 12789 2925 13606 3043
rect 12789 2903 13353 2925
rect 12789 2851 12827 2903
rect 12879 2879 13353 2903
rect 13399 2879 13511 2925
rect 13557 2903 13606 2925
rect 12879 2851 13515 2879
rect 13567 2851 13606 2903
rect 12789 2762 13606 2851
rect 12789 2716 13353 2762
rect 13399 2716 13511 2762
rect 13557 2716 13606 2762
rect 12789 2685 13606 2716
rect 12789 2633 12827 2685
rect 12879 2633 13515 2685
rect 13567 2633 13606 2685
rect 12789 2599 13606 2633
rect 12789 2553 13353 2599
rect 13399 2553 13511 2599
rect 13557 2553 13606 2599
rect 12789 2468 13606 2553
rect 12789 2416 12827 2468
rect 12879 2436 13515 2468
rect 12879 2416 13353 2436
rect 12789 2390 13353 2416
rect 13399 2390 13511 2436
rect 13567 2416 13606 2468
rect 13557 2390 13606 2416
rect 12789 2272 13606 2390
rect 12789 2250 13353 2272
rect 11893 2032 12022 2198
rect 11893 1980 11931 2032
rect 11983 1980 12022 2032
rect 11893 1814 12022 1980
rect 11893 1762 11931 1814
rect 11983 1762 12022 1814
rect 11893 1597 12022 1762
rect 11893 1545 11931 1597
rect 11983 1545 12022 1597
rect 11893 1379 12022 1545
rect 11893 1327 11931 1379
rect 11983 1327 12022 1379
rect 11893 1162 12022 1327
rect 11893 1110 11931 1162
rect 11983 1110 12022 1162
rect 11893 944 12022 1110
rect 11893 892 11931 944
rect 11983 892 12022 944
rect 11893 726 12022 892
rect 11893 674 11931 726
rect 11983 674 12022 726
rect 11893 509 12022 674
rect 11893 457 11931 509
rect 11983 457 12022 509
rect 11893 291 12022 457
rect 11893 239 11931 291
rect 11983 239 12022 291
rect 11893 199 12022 239
rect 12789 2198 12827 2250
rect 12879 2226 13353 2250
rect 13399 2226 13511 2272
rect 13557 2250 13606 2272
rect 12879 2198 13515 2226
rect 13567 2198 13606 2250
rect 12789 2109 13606 2198
rect 12789 2063 13353 2109
rect 13399 2063 13511 2109
rect 13557 2063 13606 2109
rect 12789 2032 13606 2063
rect 12789 1980 12827 2032
rect 12879 1980 13515 2032
rect 13567 1980 13606 2032
rect 12789 1946 13606 1980
rect 12789 1900 13353 1946
rect 13399 1900 13511 1946
rect 13557 1900 13606 1946
rect 12789 1814 13606 1900
rect 12789 1762 12827 1814
rect 12879 1782 13515 1814
rect 12879 1762 13353 1782
rect 12789 1736 13353 1762
rect 13399 1736 13511 1782
rect 13567 1762 13606 1814
rect 13557 1736 13606 1762
rect 12789 1619 13606 1736
rect 12789 1597 13353 1619
rect 12789 1545 12827 1597
rect 12879 1573 13353 1597
rect 13399 1573 13511 1619
rect 13557 1597 13606 1619
rect 12879 1545 13515 1573
rect 13567 1545 13606 1597
rect 12789 1456 13606 1545
rect 12789 1410 13353 1456
rect 13399 1410 13511 1456
rect 13557 1410 13606 1456
rect 12789 1379 13606 1410
rect 12789 1327 12827 1379
rect 12879 1327 13515 1379
rect 13567 1327 13606 1379
rect 12789 1293 13606 1327
rect 12789 1247 13353 1293
rect 13399 1247 13511 1293
rect 13557 1247 13606 1293
rect 12789 1162 13606 1247
rect 12789 1110 12827 1162
rect 12879 1129 13515 1162
rect 12879 1110 13353 1129
rect 12789 1083 13353 1110
rect 13399 1083 13511 1129
rect 13567 1110 13606 1162
rect 13557 1083 13606 1110
rect 12789 966 13606 1083
rect 12789 944 13353 966
rect 12789 892 12827 944
rect 12879 920 13353 944
rect 13399 920 13511 966
rect 13557 944 13606 966
rect 12879 892 13515 920
rect 13567 892 13606 944
rect 12789 803 13606 892
rect 12789 757 13353 803
rect 13399 757 13511 803
rect 13557 757 13606 803
rect 12789 726 13606 757
rect 12789 674 12827 726
rect 12879 674 13515 726
rect 13567 674 13606 726
rect 12789 640 13606 674
rect 12789 594 13353 640
rect 13399 594 13511 640
rect 13557 594 13606 640
rect 12789 509 13606 594
rect 12789 457 12827 509
rect 12879 476 13515 509
rect 12879 457 13353 476
rect 12789 430 13353 457
rect 13399 430 13511 476
rect 13567 457 13606 509
rect 13557 430 13606 457
rect 12789 313 13606 430
rect 12789 291 13353 313
rect 12789 239 12827 291
rect 12879 267 13353 291
rect 13399 267 13511 313
rect 13557 291 13606 313
rect 12879 239 13515 267
rect 13567 239 13606 291
rect 12789 199 13606 239
rect 8878 103 8926 149
rect 8972 103 9084 149
rect 9130 103 9532 149
rect 8878 37 9532 103
rect 10615 37 10731 199
rect 11511 37 11627 199
rect 11900 37 12015 199
rect 12795 150 13605 199
rect 12795 104 13353 150
rect 13399 104 13511 150
rect 13557 104 13605 150
rect 12795 37 13605 104
rect 8878 36 9533 37
rect 10614 36 10732 37
rect 11510 36 11628 37
rect 11899 36 12017 37
rect 12795 36 13606 37
rect 8878 -13 13606 36
rect 8878 -14 13353 -13
rect 8878 -60 8926 -14
rect 8972 -60 9084 -14
rect 9130 -60 9401 -14
rect 9447 -60 9559 -14
rect 9605 -60 9717 -14
rect 9763 -60 9875 -14
rect 9921 -60 10033 -14
rect 10079 -60 10191 -14
rect 10237 -60 10349 -14
rect 10395 -60 10507 -14
rect 10553 -60 10665 -14
rect 10711 -60 10824 -14
rect 10870 -60 10982 -14
rect 11028 -60 11140 -14
rect 11186 -60 11298 -14
rect 11344 -60 11456 -14
rect 11502 -60 11614 -14
rect 11660 -60 11772 -14
rect 11818 -60 11931 -14
rect 11977 -60 12089 -14
rect 12135 -60 12247 -14
rect 12293 -60 12405 -14
rect 12451 -60 12563 -14
rect 12609 -60 12721 -14
rect 12767 -60 12879 -14
rect 12925 -60 13037 -14
rect 13083 -60 13195 -14
rect 13241 -59 13353 -14
rect 13399 -59 13511 -13
rect 13557 -59 13606 -13
rect 13241 -60 13606 -59
rect 8878 -110 13606 -60
rect 9036 -111 13606 -110
rect 8999 -477 13686 -384
rect 8999 -529 10253 -477
rect 10305 -529 10465 -477
rect 10517 -529 12976 -477
rect 13028 -529 13188 -477
rect 13240 -529 13686 -477
rect 8999 -695 13686 -529
rect 8999 -747 10253 -695
rect 10305 -747 10465 -695
rect 10517 -747 12976 -695
rect 13028 -747 13188 -695
rect 13240 -747 13686 -695
rect 8999 -840 13686 -747
<< via1 >>
rect 6329 16227 6350 16238
rect 6350 16227 6381 16238
rect 6777 16227 6824 16238
rect 6824 16227 6829 16238
rect 6329 16186 6381 16227
rect 6329 15968 6381 16020
rect 6777 16186 6829 16227
rect 6777 15968 6829 16020
rect 6329 15751 6333 15803
rect 6333 15751 6379 15803
rect 6379 15751 6381 15803
rect 6329 15533 6333 15585
rect 6333 15533 6379 15585
rect 6379 15533 6381 15585
rect 6329 15315 6333 15367
rect 6333 15315 6379 15367
rect 6379 15315 6381 15367
rect 6329 15097 6333 15149
rect 6333 15097 6379 15149
rect 6379 15097 6381 15149
rect 6329 14880 6333 14932
rect 6333 14880 6379 14932
rect 6379 14880 6381 14932
rect 6329 14662 6333 14714
rect 6333 14662 6379 14714
rect 6379 14662 6381 14714
rect 7225 16186 7277 16238
rect 7225 15968 7277 16020
rect 6777 15751 6781 15803
rect 6781 15751 6827 15803
rect 6827 15751 6829 15803
rect 6777 15533 6781 15585
rect 6781 15533 6827 15585
rect 6827 15533 6829 15585
rect 6777 15315 6781 15367
rect 6781 15315 6827 15367
rect 6827 15315 6829 15367
rect 6777 15097 6781 15149
rect 6781 15097 6827 15149
rect 6827 15097 6829 15149
rect 6777 14880 6781 14932
rect 6781 14880 6827 14932
rect 6827 14880 6829 14932
rect 6777 14662 6781 14714
rect 6781 14662 6827 14714
rect 6827 14662 6829 14714
rect 6551 14381 6557 14433
rect 6557 14381 6603 14433
rect 6551 14164 6557 14216
rect 6557 14164 6603 14216
rect 6551 13946 6557 13998
rect 6557 13946 6603 13998
rect 6551 13728 6557 13780
rect 6557 13728 6603 13780
rect 6551 13511 6557 13563
rect 6557 13511 6603 13563
rect 7673 16186 7725 16238
rect 8121 16227 8135 16238
rect 8135 16227 8173 16238
rect 8569 16227 8609 16238
rect 8609 16227 8621 16238
rect 8859 16227 8880 16238
rect 8880 16227 8911 16238
rect 9307 16227 9354 16238
rect 9354 16227 9359 16238
rect 7673 15968 7725 16020
rect 7225 15751 7229 15803
rect 7229 15751 7275 15803
rect 7275 15751 7277 15803
rect 7225 15533 7229 15585
rect 7229 15533 7275 15585
rect 7275 15533 7277 15585
rect 7225 15315 7229 15367
rect 7229 15315 7275 15367
rect 7275 15315 7277 15367
rect 7225 15097 7229 15149
rect 7229 15097 7275 15149
rect 7275 15097 7277 15149
rect 7225 14880 7229 14932
rect 7229 14880 7275 14932
rect 7275 14880 7277 14932
rect 7225 14662 7229 14714
rect 7229 14662 7275 14714
rect 7275 14662 7277 14714
rect 6999 14381 7005 14433
rect 7005 14381 7051 14433
rect 6999 14164 7005 14216
rect 7005 14164 7051 14216
rect 6999 13946 7005 13998
rect 7005 13946 7051 13998
rect 6999 13728 7005 13780
rect 7005 13728 7051 13780
rect 6999 13511 7005 13563
rect 7005 13511 7051 13563
rect 8121 16186 8173 16227
rect 8121 15968 8173 16020
rect 7673 15751 7677 15803
rect 7677 15751 7723 15803
rect 7723 15751 7725 15803
rect 7673 15533 7677 15585
rect 7677 15533 7723 15585
rect 7723 15533 7725 15585
rect 7673 15315 7677 15367
rect 7677 15315 7723 15367
rect 7723 15315 7725 15367
rect 7673 15097 7677 15149
rect 7677 15097 7723 15149
rect 7723 15097 7725 15149
rect 7673 14880 7677 14932
rect 7677 14880 7723 14932
rect 7723 14880 7725 14932
rect 7673 14662 7677 14714
rect 7677 14662 7723 14714
rect 7723 14662 7725 14714
rect 7447 14381 7453 14433
rect 7453 14381 7499 14433
rect 7447 14164 7453 14216
rect 7453 14164 7499 14216
rect 7447 13946 7453 13998
rect 7453 13946 7499 13998
rect 7447 13728 7453 13780
rect 7453 13728 7499 13780
rect 7447 13511 7453 13563
rect 7453 13511 7499 13563
rect 8569 16186 8621 16227
rect 8569 15968 8621 16020
rect 8121 15751 8125 15803
rect 8125 15751 8171 15803
rect 8171 15751 8173 15803
rect 8121 15533 8125 15585
rect 8125 15533 8171 15585
rect 8171 15533 8173 15585
rect 8121 15315 8125 15367
rect 8125 15315 8171 15367
rect 8171 15315 8173 15367
rect 8121 15097 8125 15149
rect 8125 15097 8171 15149
rect 8171 15097 8173 15149
rect 8121 14880 8125 14932
rect 8125 14880 8171 14932
rect 8171 14880 8173 14932
rect 8121 14662 8125 14714
rect 8125 14662 8171 14714
rect 8171 14662 8173 14714
rect 7895 14381 7901 14433
rect 7901 14381 7947 14433
rect 7895 14164 7901 14216
rect 7901 14164 7947 14216
rect 7895 13946 7901 13998
rect 7901 13946 7947 13998
rect 7895 13728 7901 13780
rect 7901 13728 7947 13780
rect 7895 13511 7901 13563
rect 7901 13511 7947 13563
rect 8569 15751 8573 15803
rect 8573 15751 8619 15803
rect 8619 15751 8621 15803
rect 8569 15533 8573 15585
rect 8573 15533 8619 15585
rect 8619 15533 8621 15585
rect 8569 15315 8573 15367
rect 8573 15315 8619 15367
rect 8619 15315 8621 15367
rect 8569 15097 8573 15149
rect 8573 15097 8619 15149
rect 8619 15097 8621 15149
rect 8569 14880 8573 14932
rect 8573 14880 8619 14932
rect 8619 14880 8621 14932
rect 8569 14662 8573 14714
rect 8573 14662 8619 14714
rect 8619 14662 8621 14714
rect 8343 14381 8349 14433
rect 8349 14381 8395 14433
rect 8343 14164 8349 14216
rect 8349 14164 8395 14216
rect 8343 13946 8349 13998
rect 8349 13946 8395 13998
rect 8343 13728 8349 13780
rect 8349 13728 8395 13780
rect 8343 13511 8349 13563
rect 8349 13511 8395 13563
rect 8859 16186 8911 16227
rect 8859 15968 8911 16020
rect 9307 16186 9359 16227
rect 9307 15968 9359 16020
rect 8859 15751 8862 15803
rect 8862 15751 8908 15803
rect 8908 15751 8911 15803
rect 8859 15533 8862 15585
rect 8862 15533 8908 15585
rect 8908 15533 8911 15585
rect 8859 15315 8862 15367
rect 8862 15315 8908 15367
rect 8908 15315 8911 15367
rect 8859 15097 8862 15149
rect 8862 15097 8908 15149
rect 8908 15097 8911 15149
rect 8859 14880 8862 14932
rect 8862 14880 8908 14932
rect 8908 14880 8911 14932
rect 8859 14662 8862 14714
rect 8862 14662 8908 14714
rect 8908 14662 8911 14714
rect 6577 13284 6629 13336
rect 6788 13284 6840 13336
rect 7000 13284 7052 13336
rect 7211 13284 7263 13336
rect 9755 16186 9807 16238
rect 9755 15968 9807 16020
rect 9307 15751 9310 15803
rect 9310 15751 9356 15803
rect 9356 15751 9359 15803
rect 9307 15533 9310 15585
rect 9310 15533 9356 15585
rect 9356 15533 9359 15585
rect 9307 15315 9310 15367
rect 9310 15315 9356 15367
rect 9356 15315 9359 15367
rect 9307 15097 9310 15149
rect 9310 15097 9356 15149
rect 9356 15097 9359 15149
rect 9307 14880 9310 14932
rect 9310 14880 9356 14932
rect 9356 14880 9359 14932
rect 9307 14662 9310 14714
rect 9310 14662 9356 14714
rect 9356 14662 9359 14714
rect 9083 14284 9086 14336
rect 9086 14284 9132 14336
rect 9132 14284 9135 14336
rect 9083 14066 9086 14118
rect 9086 14066 9132 14118
rect 9132 14066 9135 14118
rect 9083 13848 9086 13900
rect 9086 13848 9132 13900
rect 9132 13848 9135 13900
rect 9083 13631 9086 13683
rect 9086 13631 9132 13683
rect 9132 13631 9135 13683
rect 9083 13413 9086 13465
rect 9086 13413 9132 13465
rect 9132 13413 9135 13465
rect 9083 13195 9086 13247
rect 9086 13195 9132 13247
rect 9132 13195 9135 13247
rect 9083 12978 9086 13030
rect 9086 12978 9132 13030
rect 9132 12978 9135 13030
rect 9083 12760 9086 12812
rect 9086 12760 9132 12812
rect 9132 12760 9135 12812
rect 9083 12542 9086 12594
rect 9086 12542 9132 12594
rect 9132 12542 9135 12594
rect 10203 16186 10255 16238
rect 10651 16227 10665 16238
rect 10665 16227 10703 16238
rect 11099 16227 11139 16238
rect 11139 16227 11151 16238
rect 11547 16227 11567 16238
rect 11567 16227 11599 16238
rect 11995 16227 12042 16238
rect 12042 16227 12047 16238
rect 10203 15968 10255 16020
rect 9755 15751 9758 15803
rect 9758 15751 9804 15803
rect 9804 15751 9807 15803
rect 9755 15533 9758 15585
rect 9758 15533 9804 15585
rect 9804 15533 9807 15585
rect 9755 15315 9758 15367
rect 9758 15315 9804 15367
rect 9804 15315 9807 15367
rect 9755 15097 9758 15149
rect 9758 15097 9804 15149
rect 9804 15097 9807 15149
rect 9755 14880 9758 14932
rect 9758 14880 9804 14932
rect 9804 14880 9807 14932
rect 9755 14662 9758 14714
rect 9758 14662 9804 14714
rect 9804 14662 9807 14714
rect 9531 14284 9534 14336
rect 9534 14284 9580 14336
rect 9580 14284 9583 14336
rect 9531 14066 9534 14118
rect 9534 14066 9580 14118
rect 9580 14066 9583 14118
rect 9531 13848 9534 13900
rect 9534 13848 9580 13900
rect 9580 13848 9583 13900
rect 9531 13631 9534 13683
rect 9534 13631 9580 13683
rect 9580 13631 9583 13683
rect 9531 13413 9534 13465
rect 9534 13413 9580 13465
rect 9580 13413 9583 13465
rect 9531 13195 9534 13247
rect 9534 13195 9580 13247
rect 9580 13195 9583 13247
rect 9531 12978 9534 13030
rect 9534 12978 9580 13030
rect 9580 12978 9583 13030
rect 9531 12760 9534 12812
rect 9534 12760 9580 12812
rect 9580 12760 9583 12812
rect 9531 12542 9534 12594
rect 9534 12542 9580 12594
rect 9580 12542 9583 12594
rect 10651 16186 10703 16227
rect 10651 15968 10703 16020
rect 10203 15751 10206 15803
rect 10206 15751 10252 15803
rect 10252 15751 10255 15803
rect 10203 15533 10206 15585
rect 10206 15533 10252 15585
rect 10252 15533 10255 15585
rect 10203 15315 10206 15367
rect 10206 15315 10252 15367
rect 10252 15315 10255 15367
rect 10203 15097 10206 15149
rect 10206 15097 10252 15149
rect 10252 15097 10255 15149
rect 10203 14880 10206 14932
rect 10206 14880 10252 14932
rect 10252 14880 10255 14932
rect 10203 14662 10206 14714
rect 10206 14662 10252 14714
rect 10252 14662 10255 14714
rect 9979 14284 9982 14336
rect 9982 14284 10028 14336
rect 10028 14284 10031 14336
rect 9979 14066 9982 14118
rect 9982 14066 10028 14118
rect 10028 14066 10031 14118
rect 9979 13848 9982 13900
rect 9982 13848 10028 13900
rect 10028 13848 10031 13900
rect 9979 13631 9982 13683
rect 9982 13631 10028 13683
rect 10028 13631 10031 13683
rect 9979 13413 9982 13465
rect 9982 13413 10028 13465
rect 10028 13413 10031 13465
rect 9979 13195 9982 13247
rect 9982 13195 10028 13247
rect 10028 13195 10031 13247
rect 9979 12978 9982 13030
rect 9982 12978 10028 13030
rect 10028 12978 10031 13030
rect 9979 12760 9982 12812
rect 9982 12760 10028 12812
rect 10028 12760 10031 12812
rect 9979 12542 9982 12594
rect 9982 12542 10028 12594
rect 10028 12542 10031 12594
rect 11099 16186 11151 16227
rect 11099 15968 11151 16020
rect 10651 15751 10654 15803
rect 10654 15751 10700 15803
rect 10700 15751 10703 15803
rect 10651 15533 10654 15585
rect 10654 15533 10700 15585
rect 10700 15533 10703 15585
rect 10651 15315 10654 15367
rect 10654 15315 10700 15367
rect 10700 15315 10703 15367
rect 10651 15097 10654 15149
rect 10654 15097 10700 15149
rect 10700 15097 10703 15149
rect 10651 14880 10654 14932
rect 10654 14880 10700 14932
rect 10700 14880 10703 14932
rect 10651 14662 10654 14714
rect 10654 14662 10700 14714
rect 10700 14662 10703 14714
rect 10427 14284 10430 14336
rect 10430 14284 10476 14336
rect 10476 14284 10479 14336
rect 10427 14066 10430 14118
rect 10430 14066 10476 14118
rect 10476 14066 10479 14118
rect 10427 13848 10430 13900
rect 10430 13848 10476 13900
rect 10476 13848 10479 13900
rect 10427 13631 10430 13683
rect 10430 13631 10476 13683
rect 10476 13631 10479 13683
rect 10427 13413 10430 13465
rect 10430 13413 10476 13465
rect 10476 13413 10479 13465
rect 10427 13195 10430 13247
rect 10430 13195 10476 13247
rect 10476 13195 10479 13247
rect 10427 12978 10430 13030
rect 10430 12978 10476 13030
rect 10476 12978 10479 13030
rect 10427 12760 10430 12812
rect 10430 12760 10476 12812
rect 10476 12760 10479 12812
rect 10427 12542 10430 12594
rect 10430 12542 10476 12594
rect 10476 12542 10479 12594
rect 11547 16186 11599 16227
rect 11547 15968 11599 16020
rect 11099 15751 11102 15803
rect 11102 15751 11148 15803
rect 11148 15751 11151 15803
rect 11099 15533 11102 15585
rect 11102 15533 11148 15585
rect 11148 15533 11151 15585
rect 11099 15315 11102 15367
rect 11102 15315 11148 15367
rect 11148 15315 11151 15367
rect 11099 15097 11102 15149
rect 11102 15097 11148 15149
rect 11148 15097 11151 15149
rect 11099 14880 11102 14932
rect 11102 14880 11148 14932
rect 11148 14880 11151 14932
rect 11099 14662 11102 14714
rect 11102 14662 11148 14714
rect 11148 14662 11151 14714
rect 10875 14284 10878 14336
rect 10878 14284 10924 14336
rect 10924 14284 10927 14336
rect 10875 14066 10878 14118
rect 10878 14066 10924 14118
rect 10924 14066 10927 14118
rect 10875 13848 10878 13900
rect 10878 13848 10924 13900
rect 10924 13848 10927 13900
rect 10875 13631 10878 13683
rect 10878 13631 10924 13683
rect 10924 13631 10927 13683
rect 10875 13413 10878 13465
rect 10878 13413 10924 13465
rect 10924 13413 10927 13465
rect 10875 13195 10878 13247
rect 10878 13195 10924 13247
rect 10924 13195 10927 13247
rect 10875 12978 10878 13030
rect 10878 12978 10924 13030
rect 10924 12978 10927 13030
rect 10875 12760 10878 12812
rect 10878 12760 10924 12812
rect 10924 12760 10927 12812
rect 10875 12542 10878 12594
rect 10878 12542 10924 12594
rect 10924 12542 10927 12594
rect 11995 16186 12047 16227
rect 11995 15968 12047 16020
rect 11547 15751 11550 15803
rect 11550 15751 11596 15803
rect 11596 15751 11599 15803
rect 11547 15533 11550 15585
rect 11550 15533 11596 15585
rect 11596 15533 11599 15585
rect 11547 15315 11550 15367
rect 11550 15315 11596 15367
rect 11596 15315 11599 15367
rect 11547 15097 11550 15149
rect 11550 15097 11596 15149
rect 11596 15097 11599 15149
rect 11547 14880 11550 14932
rect 11550 14880 11596 14932
rect 11596 14880 11599 14932
rect 11547 14662 11550 14714
rect 11550 14662 11596 14714
rect 11596 14662 11599 14714
rect 11323 14284 11326 14336
rect 11326 14284 11372 14336
rect 11372 14284 11375 14336
rect 11323 14066 11326 14118
rect 11326 14066 11372 14118
rect 11372 14066 11375 14118
rect 11323 13848 11326 13900
rect 11326 13848 11372 13900
rect 11372 13848 11375 13900
rect 11323 13631 11326 13683
rect 11326 13631 11372 13683
rect 11372 13631 11375 13683
rect 11323 13413 11326 13465
rect 11326 13413 11372 13465
rect 11372 13413 11375 13465
rect 11323 13195 11326 13247
rect 11326 13195 11372 13247
rect 11372 13195 11375 13247
rect 11323 12978 11326 13030
rect 11326 12978 11372 13030
rect 11372 12978 11375 13030
rect 11323 12760 11326 12812
rect 11326 12760 11372 12812
rect 11372 12760 11375 12812
rect 11323 12542 11326 12594
rect 11326 12542 11372 12594
rect 11372 12542 11375 12594
rect 12443 16186 12495 16238
rect 12443 15968 12495 16020
rect 11995 15751 11998 15803
rect 11998 15751 12044 15803
rect 12044 15751 12047 15803
rect 11995 15533 11998 15585
rect 11998 15533 12044 15585
rect 12044 15533 12047 15585
rect 11995 15315 11998 15367
rect 11998 15315 12044 15367
rect 12044 15315 12047 15367
rect 11995 15097 11998 15149
rect 11998 15097 12044 15149
rect 12044 15097 12047 15149
rect 11995 14880 11998 14932
rect 11998 14880 12044 14932
rect 12044 14880 12047 14932
rect 11995 14662 11998 14714
rect 11998 14662 12044 14714
rect 12044 14662 12047 14714
rect 11771 14284 11774 14336
rect 11774 14284 11820 14336
rect 11820 14284 11823 14336
rect 11771 14066 11774 14118
rect 11774 14066 11820 14118
rect 11820 14066 11823 14118
rect 11771 13848 11774 13900
rect 11774 13848 11820 13900
rect 11820 13848 11823 13900
rect 11771 13631 11774 13683
rect 11774 13631 11820 13683
rect 11820 13631 11823 13683
rect 11771 13413 11774 13465
rect 11774 13413 11820 13465
rect 11820 13413 11823 13465
rect 11771 13195 11774 13247
rect 11774 13195 11820 13247
rect 11820 13195 11823 13247
rect 11771 12978 11774 13030
rect 11774 12978 11820 13030
rect 11820 12978 11823 13030
rect 11771 12760 11774 12812
rect 11774 12760 11820 12812
rect 11820 12760 11823 12812
rect 11771 12542 11774 12594
rect 11774 12542 11820 12594
rect 11820 12542 11823 12594
rect 12891 16186 12943 16238
rect 13339 16227 13353 16238
rect 13353 16227 13391 16238
rect 12891 15968 12943 16020
rect 12443 15751 12446 15803
rect 12446 15751 12492 15803
rect 12492 15751 12495 15803
rect 12443 15533 12446 15585
rect 12446 15533 12492 15585
rect 12492 15533 12495 15585
rect 12443 15315 12446 15367
rect 12446 15315 12492 15367
rect 12492 15315 12495 15367
rect 12443 15097 12446 15149
rect 12446 15097 12492 15149
rect 12492 15097 12495 15149
rect 12443 14880 12446 14932
rect 12446 14880 12492 14932
rect 12492 14880 12495 14932
rect 12443 14662 12446 14714
rect 12446 14662 12492 14714
rect 12492 14662 12495 14714
rect 12219 14284 12222 14336
rect 12222 14284 12268 14336
rect 12268 14284 12271 14336
rect 12219 14066 12222 14118
rect 12222 14066 12268 14118
rect 12268 14066 12271 14118
rect 12219 13848 12222 13900
rect 12222 13848 12268 13900
rect 12268 13848 12271 13900
rect 12219 13631 12222 13683
rect 12222 13631 12268 13683
rect 12268 13631 12271 13683
rect 12219 13413 12222 13465
rect 12222 13413 12268 13465
rect 12268 13413 12271 13465
rect 12219 13195 12222 13247
rect 12222 13195 12268 13247
rect 12268 13195 12271 13247
rect 12219 12978 12222 13030
rect 12222 12978 12268 13030
rect 12268 12978 12271 13030
rect 12219 12760 12222 12812
rect 12222 12760 12268 12812
rect 12268 12760 12271 12812
rect 12219 12542 12222 12594
rect 12222 12542 12268 12594
rect 12268 12542 12271 12594
rect 13339 16186 13391 16227
rect 13339 15968 13391 16020
rect 12891 15751 12894 15803
rect 12894 15751 12940 15803
rect 12940 15751 12943 15803
rect 12891 15533 12894 15585
rect 12894 15533 12940 15585
rect 12940 15533 12943 15585
rect 12891 15315 12894 15367
rect 12894 15315 12940 15367
rect 12940 15315 12943 15367
rect 12891 15097 12894 15149
rect 12894 15097 12940 15149
rect 12940 15097 12943 15149
rect 12891 14880 12894 14932
rect 12894 14880 12940 14932
rect 12940 14880 12943 14932
rect 12891 14662 12894 14714
rect 12894 14662 12940 14714
rect 12940 14662 12943 14714
rect 12667 14284 12670 14336
rect 12670 14284 12716 14336
rect 12716 14284 12719 14336
rect 12667 14066 12670 14118
rect 12670 14066 12716 14118
rect 12716 14066 12719 14118
rect 12667 13848 12670 13900
rect 12670 13848 12716 13900
rect 12716 13848 12719 13900
rect 12667 13631 12670 13683
rect 12670 13631 12716 13683
rect 12716 13631 12719 13683
rect 12667 13413 12670 13465
rect 12670 13413 12716 13465
rect 12716 13413 12719 13465
rect 12667 13195 12670 13247
rect 12670 13195 12716 13247
rect 12716 13195 12719 13247
rect 12667 12978 12670 13030
rect 12670 12978 12716 13030
rect 12716 12978 12719 13030
rect 12667 12760 12670 12812
rect 12670 12760 12716 12812
rect 12716 12760 12719 12812
rect 12667 12542 12670 12594
rect 12670 12542 12716 12594
rect 12716 12542 12719 12594
rect 13339 15751 13342 15803
rect 13342 15751 13388 15803
rect 13388 15751 13391 15803
rect 13339 15533 13342 15585
rect 13342 15533 13388 15585
rect 13388 15533 13391 15585
rect 13339 15315 13342 15367
rect 13342 15315 13388 15367
rect 13388 15315 13391 15367
rect 13339 15097 13342 15149
rect 13342 15097 13388 15149
rect 13388 15097 13391 15149
rect 13339 14880 13342 14932
rect 13342 14880 13388 14932
rect 13388 14880 13391 14932
rect 13339 14662 13342 14714
rect 13342 14662 13388 14714
rect 13388 14662 13391 14714
rect 13115 14284 13118 14336
rect 13118 14284 13164 14336
rect 13164 14284 13167 14336
rect 13115 14066 13118 14118
rect 13118 14066 13164 14118
rect 13164 14066 13167 14118
rect 13115 13848 13118 13900
rect 13118 13848 13164 13900
rect 13164 13848 13167 13900
rect 13115 13631 13118 13683
rect 13118 13631 13164 13683
rect 13164 13631 13167 13683
rect 13115 13413 13118 13465
rect 13118 13413 13164 13465
rect 13164 13413 13167 13465
rect 13115 13195 13118 13247
rect 13118 13195 13164 13247
rect 13164 13195 13167 13247
rect 13115 12978 13118 13030
rect 13118 12978 13164 13030
rect 13164 12978 13167 13030
rect 13115 12760 13118 12812
rect 13118 12760 13164 12812
rect 13164 12760 13167 12812
rect 13115 12542 13118 12594
rect 13118 12542 13164 12594
rect 13164 12542 13167 12594
rect 9142 12158 9194 12170
rect 9353 12158 9405 12170
rect 9564 12158 9616 12170
rect 9774 12158 9826 12170
rect 9985 12158 10037 12170
rect 10197 12158 10249 12170
rect 10408 12158 10460 12170
rect 10618 12158 10670 12170
rect 10829 12158 10881 12170
rect 11040 12158 11092 12170
rect 9142 12118 9194 12158
rect 9353 12118 9405 12158
rect 9564 12118 9616 12158
rect 9774 12118 9826 12158
rect 9985 12118 10037 12158
rect 10197 12118 10249 12158
rect 10408 12118 10460 12158
rect 10618 12118 10670 12158
rect 10829 12118 10881 12158
rect 11040 12118 11092 12158
rect 6314 11269 6323 11293
rect 6323 11269 6366 11293
rect 6314 11241 6366 11269
rect 9142 11438 9194 11477
rect 9353 11438 9405 11477
rect 9564 11438 9616 11477
rect 9774 11438 9826 11477
rect 9985 11438 10037 11477
rect 10197 11438 10249 11477
rect 10408 11438 10460 11477
rect 10618 11438 10670 11477
rect 10829 11438 10881 11477
rect 11040 11438 11092 11477
rect 9142 11425 9194 11438
rect 9353 11425 9405 11438
rect 9564 11425 9616 11438
rect 9774 11425 9826 11438
rect 9985 11425 10037 11438
rect 10197 11425 10249 11438
rect 10408 11425 10460 11438
rect 10618 11425 10670 11438
rect 10829 11425 10881 11438
rect 11040 11425 11092 11438
rect 6607 11148 6659 11200
rect 6818 11160 6870 11200
rect 7030 11160 7082 11200
rect 7241 11160 7293 11200
rect 6818 11148 6870 11160
rect 7030 11148 7082 11160
rect 7241 11148 7293 11160
rect 6314 11023 6366 11075
rect 6314 10825 6366 10858
rect 6314 10806 6323 10825
rect 6323 10806 6366 10825
rect 6314 10616 6323 10640
rect 6323 10616 6366 10640
rect 6314 10588 6366 10616
rect 6314 10370 6366 10422
rect 6314 10172 6366 10205
rect 6314 10153 6323 10172
rect 6323 10153 6366 10172
rect 6314 9963 6323 9987
rect 6323 9963 6366 9987
rect 6314 9935 6366 9963
rect 6846 10863 6849 10915
rect 6849 10863 6895 10915
rect 6895 10863 6898 10915
rect 6846 10645 6849 10697
rect 6849 10645 6895 10697
rect 6895 10645 6898 10697
rect 6846 10428 6849 10480
rect 6849 10428 6895 10480
rect 6895 10428 6898 10480
rect 6846 10210 6849 10262
rect 6849 10210 6895 10262
rect 6895 10210 6898 10262
rect 6846 9992 6849 10044
rect 6849 9992 6895 10044
rect 6895 9992 6898 10044
rect 6846 9775 6849 9827
rect 6849 9775 6895 9827
rect 6895 9775 6898 9827
rect 6846 9557 6849 9609
rect 6849 9557 6895 9609
rect 6895 9557 6898 9609
rect 7293 10863 7297 10915
rect 7297 10863 7343 10915
rect 7343 10863 7345 10915
rect 7293 10645 7297 10697
rect 7297 10645 7343 10697
rect 7343 10645 7345 10697
rect 7293 10428 7297 10480
rect 7297 10428 7343 10480
rect 7343 10428 7345 10480
rect 7070 10210 7073 10262
rect 7073 10210 7119 10262
rect 7119 10210 7122 10262
rect 7070 9992 7073 10044
rect 7073 9992 7119 10044
rect 7119 9992 7122 10044
rect 7070 9774 7073 9826
rect 7073 9774 7119 9826
rect 7119 9774 7122 9826
rect 7070 9556 7073 9608
rect 7073 9556 7119 9608
rect 7119 9556 7122 9608
rect 7293 10210 7297 10262
rect 7297 10210 7343 10262
rect 7343 10210 7345 10262
rect 7293 9992 7297 10044
rect 7297 9992 7343 10044
rect 7343 9992 7345 10044
rect 7293 9775 7297 9827
rect 7297 9775 7343 9827
rect 7343 9775 7345 9827
rect 7293 9557 7297 9609
rect 7297 9557 7343 9609
rect 7343 9557 7345 9609
rect 7741 10863 7745 10915
rect 7745 10863 7791 10915
rect 7791 10863 7793 10915
rect 7741 10645 7745 10697
rect 7745 10645 7791 10697
rect 7791 10645 7793 10697
rect 9083 11143 9086 11195
rect 9086 11143 9132 11195
rect 9132 11143 9135 11195
rect 9083 10926 9086 10978
rect 9086 10926 9132 10978
rect 9132 10926 9135 10978
rect 9083 10708 9086 10760
rect 9086 10708 9132 10760
rect 9132 10708 9135 10760
rect 8861 10541 8862 10593
rect 8862 10541 8908 10593
rect 8908 10541 8913 10593
rect 7741 10428 7745 10480
rect 7745 10428 7791 10480
rect 7791 10428 7793 10480
rect 7517 10210 7521 10262
rect 7521 10210 7567 10262
rect 7567 10210 7569 10262
rect 7517 9992 7521 10044
rect 7521 9992 7567 10044
rect 7567 9992 7569 10044
rect 7517 9774 7521 9826
rect 7521 9774 7567 9826
rect 7567 9774 7569 9826
rect 7517 9556 7521 9608
rect 7521 9556 7567 9608
rect 7567 9556 7569 9608
rect 7741 10210 7745 10262
rect 7745 10210 7791 10262
rect 7791 10210 7793 10262
rect 7741 9992 7745 10044
rect 7745 9992 7791 10044
rect 7791 9992 7793 10044
rect 7741 9775 7745 9827
rect 7745 9775 7791 9827
rect 7791 9775 7793 9827
rect 7741 9557 7745 9609
rect 7745 9557 7791 9609
rect 7791 9557 7793 9609
rect 8017 10427 8069 10474
rect 8229 10427 8281 10474
rect 8017 10422 8045 10427
rect 8045 10422 8069 10427
rect 8229 10422 8249 10427
rect 8249 10422 8281 10427
rect 8017 10218 8045 10257
rect 8045 10218 8069 10257
rect 8229 10218 8249 10257
rect 8249 10218 8281 10257
rect 8017 10205 8069 10218
rect 8229 10205 8281 10218
rect 8017 9987 8069 10039
rect 8229 9987 8281 10039
rect 8861 10323 8862 10375
rect 8862 10323 8908 10375
rect 8908 10323 8913 10375
rect 8861 10105 8862 10157
rect 8862 10105 8908 10157
rect 8908 10105 8913 10157
rect 9083 10490 9086 10542
rect 9086 10490 9132 10542
rect 9132 10490 9135 10542
rect 9083 10272 9086 10324
rect 9086 10272 9132 10324
rect 9132 10272 9135 10324
rect 9083 10055 9086 10107
rect 9086 10055 9132 10107
rect 9132 10055 9135 10107
rect 8861 9887 8862 9939
rect 8862 9887 8908 9939
rect 8908 9887 8913 9939
rect 9531 11143 9534 11195
rect 9534 11143 9580 11195
rect 9580 11143 9583 11195
rect 9531 10926 9534 10978
rect 9534 10926 9580 10978
rect 9580 10926 9583 10978
rect 9531 10708 9534 10760
rect 9534 10708 9580 10760
rect 9580 10708 9583 10760
rect 9309 10541 9310 10593
rect 9310 10541 9356 10593
rect 9356 10541 9361 10593
rect 9309 10323 9310 10375
rect 9310 10323 9356 10375
rect 9356 10323 9361 10375
rect 9309 10105 9310 10157
rect 9310 10105 9356 10157
rect 9356 10105 9361 10157
rect 9531 10490 9534 10542
rect 9534 10490 9580 10542
rect 9580 10490 9583 10542
rect 9531 10272 9534 10324
rect 9534 10272 9580 10324
rect 9580 10272 9583 10324
rect 9531 10055 9534 10107
rect 9534 10055 9580 10107
rect 9580 10055 9583 10107
rect 9309 9887 9310 9939
rect 9310 9887 9356 9939
rect 9356 9887 9361 9939
rect 9979 11143 9982 11195
rect 9982 11143 10028 11195
rect 10028 11143 10031 11195
rect 9979 10926 9982 10978
rect 9982 10926 10028 10978
rect 10028 10926 10031 10978
rect 9979 10708 9982 10760
rect 9982 10708 10028 10760
rect 10028 10708 10031 10760
rect 9757 10541 9758 10593
rect 9758 10541 9804 10593
rect 9804 10541 9809 10593
rect 9757 10323 9758 10375
rect 9758 10323 9804 10375
rect 9804 10323 9809 10375
rect 9757 10105 9758 10157
rect 9758 10105 9804 10157
rect 9804 10105 9809 10157
rect 9979 10490 9982 10542
rect 9982 10490 10028 10542
rect 10028 10490 10031 10542
rect 9979 10272 9982 10324
rect 9982 10272 10028 10324
rect 10028 10272 10031 10324
rect 9979 10055 9982 10107
rect 9982 10055 10028 10107
rect 10028 10055 10031 10107
rect 9757 9887 9758 9939
rect 9758 9887 9804 9939
rect 9804 9887 9809 9939
rect 10427 11143 10430 11195
rect 10430 11143 10476 11195
rect 10476 11143 10479 11195
rect 10427 10926 10430 10978
rect 10430 10926 10476 10978
rect 10476 10926 10479 10978
rect 10427 10708 10430 10760
rect 10430 10708 10476 10760
rect 10476 10708 10479 10760
rect 10205 10541 10206 10593
rect 10206 10541 10252 10593
rect 10252 10541 10257 10593
rect 10205 10323 10206 10375
rect 10206 10323 10252 10375
rect 10252 10323 10257 10375
rect 10205 10105 10206 10157
rect 10206 10105 10252 10157
rect 10252 10105 10257 10157
rect 10427 10490 10430 10542
rect 10430 10490 10476 10542
rect 10476 10490 10479 10542
rect 10427 10272 10430 10324
rect 10430 10272 10476 10324
rect 10476 10272 10479 10324
rect 10427 10055 10430 10107
rect 10430 10055 10476 10107
rect 10476 10055 10479 10107
rect 10205 9887 10206 9939
rect 10206 9887 10252 9939
rect 10252 9887 10257 9939
rect 10875 11143 10878 11195
rect 10878 11143 10924 11195
rect 10924 11143 10927 11195
rect 10875 10926 10878 10978
rect 10878 10926 10924 10978
rect 10924 10926 10927 10978
rect 10875 10708 10878 10760
rect 10878 10708 10924 10760
rect 10924 10708 10927 10760
rect 10653 10541 10654 10593
rect 10654 10541 10700 10593
rect 10700 10541 10705 10593
rect 10653 10323 10654 10375
rect 10654 10323 10700 10375
rect 10700 10323 10705 10375
rect 10653 10105 10654 10157
rect 10654 10105 10700 10157
rect 10700 10105 10705 10157
rect 10875 10490 10878 10542
rect 10878 10490 10924 10542
rect 10924 10490 10927 10542
rect 10875 10272 10878 10324
rect 10878 10272 10924 10324
rect 10924 10272 10927 10324
rect 10875 10055 10878 10107
rect 10878 10055 10924 10107
rect 10924 10055 10927 10107
rect 10653 9887 10654 9939
rect 10654 9887 10700 9939
rect 10700 9887 10705 9939
rect 11323 11143 11326 11195
rect 11326 11143 11372 11195
rect 11372 11143 11375 11195
rect 11323 10926 11326 10978
rect 11326 10926 11372 10978
rect 11372 10926 11375 10978
rect 11323 10708 11326 10760
rect 11326 10708 11372 10760
rect 11372 10708 11375 10760
rect 11101 10541 11102 10593
rect 11102 10541 11148 10593
rect 11148 10541 11153 10593
rect 11101 10323 11102 10375
rect 11102 10323 11148 10375
rect 11148 10323 11153 10375
rect 11101 10105 11102 10157
rect 11102 10105 11148 10157
rect 11148 10105 11153 10157
rect 11323 10490 11326 10542
rect 11326 10490 11372 10542
rect 11372 10490 11375 10542
rect 11323 10272 11326 10324
rect 11326 10272 11372 10324
rect 11372 10272 11375 10324
rect 11323 10055 11326 10107
rect 11326 10055 11372 10107
rect 11372 10055 11375 10107
rect 11101 9887 11102 9939
rect 11102 9887 11148 9939
rect 11148 9887 11153 9939
rect 11771 11143 11774 11195
rect 11774 11143 11820 11195
rect 11820 11143 11823 11195
rect 11771 10926 11774 10978
rect 11774 10926 11820 10978
rect 11820 10926 11823 10978
rect 11771 10708 11774 10760
rect 11774 10708 11820 10760
rect 11820 10708 11823 10760
rect 11549 10541 11550 10593
rect 11550 10541 11596 10593
rect 11596 10541 11601 10593
rect 11549 10323 11550 10375
rect 11550 10323 11596 10375
rect 11596 10323 11601 10375
rect 11549 10105 11550 10157
rect 11550 10105 11596 10157
rect 11596 10105 11601 10157
rect 11771 10490 11774 10542
rect 11774 10490 11820 10542
rect 11820 10490 11823 10542
rect 11771 10272 11774 10324
rect 11774 10272 11820 10324
rect 11820 10272 11823 10324
rect 11771 10055 11774 10107
rect 11774 10055 11820 10107
rect 11820 10055 11823 10107
rect 11549 9887 11550 9939
rect 11550 9887 11596 9939
rect 11596 9887 11601 9939
rect 12219 11143 12222 11195
rect 12222 11143 12268 11195
rect 12268 11143 12271 11195
rect 12219 10926 12222 10978
rect 12222 10926 12268 10978
rect 12268 10926 12271 10978
rect 12219 10708 12222 10760
rect 12222 10708 12268 10760
rect 12268 10708 12271 10760
rect 11997 10541 11998 10593
rect 11998 10541 12044 10593
rect 12044 10541 12049 10593
rect 11997 10323 11998 10375
rect 11998 10323 12044 10375
rect 12044 10323 12049 10375
rect 11997 10105 11998 10157
rect 11998 10105 12044 10157
rect 12044 10105 12049 10157
rect 12219 10490 12222 10542
rect 12222 10490 12268 10542
rect 12268 10490 12271 10542
rect 12219 10272 12222 10324
rect 12222 10272 12268 10324
rect 12268 10272 12271 10324
rect 12219 10055 12222 10107
rect 12222 10055 12268 10107
rect 12268 10055 12271 10107
rect 11997 9887 11998 9939
rect 11998 9887 12044 9939
rect 12044 9887 12049 9939
rect 12667 11143 12670 11195
rect 12670 11143 12716 11195
rect 12716 11143 12719 11195
rect 12667 10926 12670 10978
rect 12670 10926 12716 10978
rect 12716 10926 12719 10978
rect 12667 10708 12670 10760
rect 12670 10708 12716 10760
rect 12716 10708 12719 10760
rect 12445 10541 12446 10593
rect 12446 10541 12492 10593
rect 12492 10541 12497 10593
rect 12445 10323 12446 10375
rect 12446 10323 12492 10375
rect 12492 10323 12497 10375
rect 12445 10105 12446 10157
rect 12446 10105 12492 10157
rect 12492 10105 12497 10157
rect 12667 10490 12670 10542
rect 12670 10490 12716 10542
rect 12716 10490 12719 10542
rect 12667 10272 12670 10324
rect 12670 10272 12716 10324
rect 12716 10272 12719 10324
rect 12667 10055 12670 10107
rect 12670 10055 12716 10107
rect 12716 10055 12719 10107
rect 12445 9887 12446 9939
rect 12446 9887 12492 9939
rect 12492 9887 12497 9939
rect 13115 11143 13118 11195
rect 13118 11143 13164 11195
rect 13164 11143 13167 11195
rect 13115 10926 13118 10978
rect 13118 10926 13164 10978
rect 13164 10926 13167 10978
rect 13115 10708 13118 10760
rect 13118 10708 13164 10760
rect 13164 10708 13167 10760
rect 12893 10541 12894 10593
rect 12894 10541 12940 10593
rect 12940 10541 12945 10593
rect 12893 10323 12894 10375
rect 12894 10323 12940 10375
rect 12940 10323 12945 10375
rect 12893 10105 12894 10157
rect 12894 10105 12940 10157
rect 12940 10105 12945 10157
rect 13115 10490 13118 10542
rect 13118 10490 13164 10542
rect 13164 10490 13167 10542
rect 13115 10272 13118 10324
rect 13118 10272 13164 10324
rect 13164 10272 13167 10324
rect 13115 10055 13118 10107
rect 13118 10055 13164 10107
rect 13164 10055 13167 10107
rect 12893 9887 12894 9939
rect 12894 9887 12940 9939
rect 12940 9887 12945 9939
rect 13640 10617 13692 10627
rect 13339 10541 13342 10593
rect 13342 10541 13388 10593
rect 13388 10541 13391 10593
rect 13640 10575 13643 10617
rect 13643 10575 13689 10617
rect 13689 10575 13692 10617
rect 13640 10407 13643 10409
rect 13643 10407 13689 10409
rect 13689 10407 13692 10409
rect 13339 10323 13342 10375
rect 13342 10323 13388 10375
rect 13388 10323 13391 10375
rect 13640 10357 13692 10407
rect 13339 10105 13342 10157
rect 13342 10105 13388 10157
rect 13388 10105 13391 10157
rect 13640 10139 13692 10191
rect 13640 9964 13692 9973
rect 13339 9887 13342 9939
rect 13342 9887 13388 9939
rect 13388 9887 13391 9939
rect 13640 9921 13643 9964
rect 13643 9921 13689 9964
rect 13689 9921 13692 9964
rect 8017 9774 8069 9821
rect 8229 9774 8281 9821
rect 8017 9769 8045 9774
rect 8045 9769 8069 9774
rect 8229 9769 8249 9774
rect 8249 9769 8281 9774
rect 8017 9564 8045 9604
rect 8045 9564 8069 9604
rect 8229 9564 8249 9604
rect 8249 9564 8281 9604
rect 8017 9552 8069 9564
rect 8229 9552 8281 9564
rect 457 8206 509 8258
rect 668 8206 720 8258
rect 878 8206 930 8258
rect 1089 8206 1141 8258
rect 1300 8206 1352 8258
rect 1511 8206 1563 8258
rect 1722 8206 1774 8258
rect 1932 8206 1984 8258
rect 2143 8206 2195 8258
rect 2355 8206 2407 8258
rect 2566 8206 2618 8258
rect 2776 8206 2828 8258
rect 2987 8206 3039 8258
rect 3198 8206 3250 8258
rect 3409 8206 3461 8258
rect 3620 8206 3672 8258
rect 3830 8206 3882 8258
rect 4041 8206 4093 8258
rect 457 7988 509 8040
rect 668 7988 720 8040
rect 878 7988 930 8040
rect 1089 7988 1141 8040
rect 1300 7988 1352 8040
rect 1511 7988 1563 8040
rect 1722 7988 1774 8040
rect 1932 7988 1984 8040
rect 2143 7988 2195 8040
rect 2355 7988 2407 8040
rect 2566 7988 2618 8040
rect 2776 7988 2828 8040
rect 2987 7988 3039 8040
rect 3198 7988 3250 8040
rect 3409 7988 3461 8040
rect 3620 7988 3672 8040
rect 3830 7988 3882 8040
rect 4041 7988 4093 8040
rect 9672 8938 9675 8990
rect 9675 8938 9721 8990
rect 9721 8938 9724 8990
rect 9672 8720 9675 8772
rect 9675 8720 9721 8772
rect 9721 8720 9724 8772
rect 457 7770 509 7822
rect 668 7770 720 7822
rect 878 7770 930 7822
rect 1089 7770 1141 7822
rect 1300 7770 1352 7822
rect 1511 7770 1563 7822
rect 1722 7770 1774 7822
rect 1932 7770 1984 7822
rect 2143 7770 2195 7822
rect 2355 7770 2407 7822
rect 2566 7770 2618 7822
rect 2776 7770 2828 7822
rect 2987 7770 3039 7822
rect 3198 7770 3250 7822
rect 3409 7770 3461 7822
rect 3620 7770 3672 7822
rect 3830 7770 3882 7822
rect 4041 7770 4093 7822
rect 5411 7861 5463 7913
rect 5623 7861 5675 7913
rect 7118 8101 7170 8153
rect 7118 7883 7170 7935
rect 8977 8353 9029 8395
rect 8977 8343 8982 8353
rect 8982 8343 9028 8353
rect 9028 8343 9029 8353
rect 9189 8343 9241 8395
rect 9448 8343 9451 8395
rect 9451 8343 9497 8395
rect 9497 8343 9500 8395
rect 8977 8144 8982 8178
rect 8982 8144 9028 8178
rect 9028 8144 9029 8178
rect 8977 8126 9029 8144
rect 9189 8126 9241 8178
rect 9448 8126 9451 8178
rect 9451 8126 9497 8178
rect 9497 8126 9500 8178
rect 6192 7345 6240 7391
rect 6240 7345 6244 7391
rect 6404 7345 6444 7391
rect 6444 7345 6456 7391
rect 6192 7339 6244 7345
rect 6404 7339 6456 7345
rect 4976 7013 5028 7065
rect 743 6809 795 6861
rect 954 6809 1006 6861
rect 1164 6809 1216 6861
rect 1375 6809 1427 6861
rect 1586 6809 1638 6861
rect 1797 6809 1849 6861
rect 2008 6809 2060 6861
rect 2218 6809 2270 6861
rect 2429 6809 2481 6861
rect 2641 6809 2693 6861
rect 2852 6809 2904 6861
rect 3062 6809 3114 6861
rect 3273 6809 3325 6861
rect 3484 6809 3536 6861
rect 3695 6809 3747 6861
rect 3906 6809 3958 6861
rect 4116 6809 4168 6861
rect 4327 6809 4379 6861
rect 743 6591 795 6643
rect 954 6591 1006 6643
rect 1164 6591 1216 6643
rect 1375 6591 1427 6643
rect 1586 6591 1638 6643
rect 1797 6591 1849 6643
rect 2008 6591 2060 6643
rect 2218 6591 2270 6643
rect 2429 6591 2481 6643
rect 2641 6591 2693 6643
rect 2852 6591 2904 6643
rect 3062 6591 3114 6643
rect 3273 6591 3325 6643
rect 3484 6591 3536 6643
rect 3695 6591 3747 6643
rect 3906 6591 3958 6643
rect 4116 6591 4168 6643
rect 4327 6591 4379 6643
rect 4976 6795 5028 6847
rect 4976 6577 5028 6629
rect 6894 7212 6897 7222
rect 6897 7212 6943 7222
rect 6943 7212 6946 7222
rect 6894 7170 6946 7212
rect 6894 7000 6897 7004
rect 6897 7000 6943 7004
rect 6943 7000 6946 7004
rect 6894 6952 6946 7000
rect 6386 6805 6438 6857
rect 5431 6678 5483 6730
rect 5431 6460 5483 6512
rect 6386 6587 6438 6639
rect 4840 5968 4892 6020
rect 5052 5978 5054 6020
rect 5054 5978 5100 6020
rect 5100 5978 5104 6020
rect 5052 5968 5104 5978
rect 743 5825 795 5877
rect 954 5825 1006 5877
rect 1164 5825 1216 5877
rect 1375 5825 1427 5877
rect 1586 5825 1638 5877
rect 1797 5825 1849 5877
rect 2008 5825 2060 5877
rect 2218 5825 2270 5877
rect 2429 5825 2481 5877
rect 2641 5825 2693 5877
rect 2852 5825 2904 5877
rect 3062 5825 3114 5877
rect 3273 5825 3325 5877
rect 3484 5825 3536 5877
rect 3695 5825 3747 5877
rect 3906 5825 3958 5877
rect 4116 5825 4168 5877
rect 4327 5825 4379 5877
rect 6386 6375 6429 6421
rect 6429 6375 6438 6421
rect 6386 6369 6438 6375
rect 7831 8031 7883 8083
rect 7831 7821 7883 7865
rect 7831 7813 7874 7821
rect 7874 7813 7883 7821
rect 8977 7908 9029 7960
rect 9189 7908 9241 7960
rect 9448 7908 9451 7960
rect 9451 7908 9497 7960
rect 9497 7908 9500 7960
rect 8977 7700 9029 7743
rect 8977 7691 8982 7700
rect 8982 7691 9028 7700
rect 9028 7691 9029 7700
rect 9189 7691 9241 7743
rect 9448 7691 9451 7743
rect 9451 7691 9497 7743
rect 9497 7691 9500 7743
rect 7118 7046 7170 7075
rect 7118 7023 7121 7046
rect 7121 7023 7167 7046
rect 7167 7023 7170 7046
rect 7118 6834 7170 6857
rect 7118 6805 7121 6834
rect 7121 6805 7167 6834
rect 7167 6805 7170 6834
rect 7118 6622 7170 6639
rect 7118 6587 7121 6622
rect 7121 6587 7167 6622
rect 7167 6587 7170 6622
rect 7118 6410 7170 6421
rect 7118 6369 7121 6410
rect 7121 6369 7167 6410
rect 7167 6369 7170 6410
rect 8977 7490 8982 7525
rect 8982 7490 9028 7525
rect 9028 7490 9029 7525
rect 8977 7473 9029 7490
rect 9189 7473 9241 7525
rect 9448 7473 9451 7525
rect 9451 7473 9497 7525
rect 9497 7473 9500 7525
rect 7831 7376 7883 7428
rect 7831 7158 7883 7210
rect 8977 7255 9029 7307
rect 9189 7255 9241 7307
rect 9448 7255 9451 7307
rect 9451 7255 9497 7307
rect 9497 7255 9500 7307
rect 6894 6066 6946 6118
rect 6386 5918 6438 5970
rect 6894 5848 6946 5900
rect 743 5607 795 5659
rect 954 5607 1006 5659
rect 1164 5607 1216 5659
rect 1375 5607 1427 5659
rect 1586 5607 1638 5659
rect 1797 5607 1849 5659
rect 2008 5607 2060 5659
rect 2218 5607 2270 5659
rect 2429 5607 2481 5659
rect 2641 5607 2693 5659
rect 2852 5607 2904 5659
rect 3062 5607 3114 5659
rect 3273 5607 3325 5659
rect 3484 5607 3536 5659
rect 3695 5607 3747 5659
rect 3906 5607 3958 5659
rect 4116 5607 4168 5659
rect 4327 5607 4379 5659
rect 5200 5574 5204 5626
rect 5204 5574 5250 5626
rect 5250 5574 5252 5626
rect 5200 5356 5252 5408
rect 5789 5765 5834 5807
rect 5834 5765 5841 5807
rect 5789 5755 5841 5765
rect 5789 5537 5841 5589
rect 6386 5707 6438 5752
rect 8977 7046 9029 7089
rect 8977 7037 8982 7046
rect 8982 7037 9028 7046
rect 9028 7037 9029 7046
rect 9189 7037 9241 7089
rect 9448 7037 9451 7089
rect 9451 7037 9497 7089
rect 9497 7037 9500 7089
rect 8977 6837 8982 6872
rect 8982 6837 9028 6872
rect 9028 6837 9029 6872
rect 8977 6820 9029 6837
rect 9189 6820 9241 6872
rect 9448 6820 9451 6872
rect 9451 6820 9497 6872
rect 9497 6820 9500 6872
rect 8977 6602 9029 6654
rect 9189 6602 9241 6654
rect 9448 6602 9451 6654
rect 9451 6602 9497 6654
rect 9497 6602 9500 6654
rect 8977 6394 9029 6437
rect 8977 6385 8982 6394
rect 8982 6385 9028 6394
rect 9028 6385 9029 6394
rect 9189 6385 9241 6437
rect 9448 6385 9451 6437
rect 9451 6385 9497 6437
rect 9497 6385 9500 6437
rect 6386 5700 6429 5707
rect 6429 5700 6438 5707
rect 10122 8938 10123 8990
rect 10123 8938 10169 8990
rect 10169 8938 10174 8990
rect 10122 8720 10123 8772
rect 10123 8720 10169 8772
rect 10169 8720 10174 8772
rect 9896 8343 9899 8395
rect 9899 8343 9945 8395
rect 9945 8343 9948 8395
rect 9896 8126 9899 8178
rect 9899 8126 9945 8178
rect 9945 8126 9948 8178
rect 9896 7908 9899 7960
rect 9899 7908 9945 7960
rect 9945 7908 9948 7960
rect 9896 7691 9899 7743
rect 9899 7691 9945 7743
rect 9945 7691 9948 7743
rect 9896 7473 9899 7525
rect 9899 7473 9945 7525
rect 9945 7473 9948 7525
rect 9896 7255 9899 7307
rect 9899 7255 9945 7307
rect 9945 7255 9948 7307
rect 9896 7037 9899 7089
rect 9899 7037 9945 7089
rect 9945 7037 9948 7089
rect 9896 6820 9899 6872
rect 9899 6820 9945 6872
rect 9945 6820 9948 6872
rect 9896 6602 9899 6654
rect 9899 6602 9945 6654
rect 9945 6602 9948 6654
rect 9896 6385 9899 6437
rect 9899 6385 9945 6437
rect 9945 6385 9948 6437
rect 8623 5156 8675 5208
rect 8835 5156 8887 5208
rect 9784 5109 9836 5161
rect 255 4885 307 4937
rect 466 4885 518 4937
rect 677 4885 729 4937
rect 887 4885 939 4937
rect 1098 4885 1150 4937
rect 1309 4885 1361 4937
rect 1520 4885 1572 4937
rect 1731 4885 1783 4937
rect 1941 4885 1993 4937
rect 2152 4885 2204 4937
rect 2363 4885 2415 4937
rect 2574 4885 2626 4937
rect 2785 4885 2837 4937
rect 2996 4885 3048 4937
rect 3207 4885 3259 4937
rect 3418 4885 3470 4937
rect 3629 4885 3681 4937
rect 3839 4885 3891 4937
rect 4050 4885 4102 4937
rect 4261 4885 4313 4937
rect 4472 4885 4524 4937
rect 4683 4885 4735 4937
rect 4893 4885 4945 4937
rect 5104 4885 5156 4937
rect 5315 4885 5367 4937
rect 255 4667 307 4719
rect 466 4667 518 4719
rect 677 4667 729 4719
rect 887 4667 939 4719
rect 1098 4667 1150 4719
rect 1309 4667 1361 4719
rect 1520 4667 1572 4719
rect 1731 4667 1783 4719
rect 1941 4667 1993 4719
rect 2152 4667 2204 4719
rect 2363 4667 2415 4719
rect 2574 4667 2626 4719
rect 2785 4667 2837 4719
rect 2996 4667 3048 4719
rect 3207 4667 3259 4719
rect 3418 4667 3470 4719
rect 3629 4667 3681 4719
rect 3839 4667 3891 4719
rect 4050 4667 4102 4719
rect 4261 4667 4313 4719
rect 4472 4667 4524 4719
rect 4683 4667 4735 4719
rect 4893 4667 4945 4719
rect 5104 4667 5156 4719
rect 5315 4667 5367 4719
rect 255 4449 307 4501
rect 466 4449 518 4501
rect 677 4449 729 4501
rect 887 4449 939 4501
rect 1098 4449 1150 4501
rect 1309 4449 1361 4501
rect 1520 4449 1572 4501
rect 1731 4449 1783 4501
rect 1941 4449 1993 4501
rect 2152 4449 2204 4501
rect 2363 4449 2415 4501
rect 2574 4449 2626 4501
rect 2785 4449 2837 4501
rect 2996 4449 3048 4501
rect 3207 4449 3259 4501
rect 3418 4449 3470 4501
rect 3629 4449 3681 4501
rect 3839 4449 3891 4501
rect 4050 4449 4102 4501
rect 4261 4449 4313 4501
rect 4472 4449 4524 4501
rect 4683 4449 4735 4501
rect 4893 4449 4945 4501
rect 5104 4449 5156 4501
rect 5315 4449 5367 4501
rect 255 4231 307 4283
rect 466 4231 518 4283
rect 677 4231 729 4283
rect 887 4231 939 4283
rect 1098 4231 1150 4283
rect 1309 4231 1361 4283
rect 1520 4231 1572 4283
rect 1731 4231 1783 4283
rect 1941 4231 1993 4283
rect 2152 4231 2204 4283
rect 2363 4231 2415 4283
rect 2574 4231 2626 4283
rect 2785 4231 2837 4283
rect 2996 4231 3048 4283
rect 3207 4231 3259 4283
rect 3418 4231 3470 4283
rect 3629 4231 3681 4283
rect 3839 4231 3891 4283
rect 4050 4231 4102 4283
rect 4261 4231 4313 4283
rect 4472 4231 4524 4283
rect 4683 4231 4735 4283
rect 4893 4231 4945 4283
rect 5104 4231 5156 4283
rect 5315 4231 5367 4283
rect 9784 4891 9836 4943
rect 10010 5109 10062 5161
rect 10010 4891 10062 4943
rect 8981 4649 9033 4701
rect 9454 4706 9497 4734
rect 9497 4706 9506 4734
rect 9193 4649 9245 4701
rect 9454 4682 9506 4706
rect 10647 9045 10650 9097
rect 10650 9045 10696 9097
rect 10696 9045 10699 9097
rect 10647 8827 10650 8879
rect 10650 8827 10696 8879
rect 10696 8827 10699 8879
rect 10647 8609 10650 8661
rect 10650 8609 10696 8661
rect 10696 8609 10699 8661
rect 10647 8392 10650 8444
rect 10650 8392 10696 8444
rect 10696 8392 10699 8444
rect 10647 8174 10650 8226
rect 10650 8174 10696 8226
rect 10696 8174 10699 8226
rect 10647 7956 10650 8008
rect 10650 7956 10696 8008
rect 10696 7956 10699 8008
rect 10647 7739 10650 7791
rect 10650 7739 10696 7791
rect 10696 7739 10699 7791
rect 10647 7521 10650 7573
rect 10650 7521 10696 7573
rect 10696 7521 10699 7573
rect 10647 7304 10650 7356
rect 10650 7304 10696 7356
rect 10696 7304 10699 7356
rect 10647 7086 10650 7138
rect 10650 7086 10696 7138
rect 10696 7086 10699 7138
rect 10647 6868 10650 6920
rect 10650 6868 10696 6920
rect 10696 6868 10699 6920
rect 10647 6650 10650 6702
rect 10650 6650 10696 6702
rect 10696 6650 10699 6702
rect 10647 6433 10650 6485
rect 10650 6433 10696 6485
rect 10696 6433 10699 6485
rect 11095 9045 11098 9097
rect 11098 9045 11144 9097
rect 11144 9045 11147 9097
rect 11095 8827 11098 8879
rect 11098 8827 11144 8879
rect 11144 8827 11147 8879
rect 11095 8609 11098 8661
rect 11098 8609 11144 8661
rect 11144 8609 11147 8661
rect 10871 8334 10874 8386
rect 10874 8334 10920 8386
rect 10920 8334 10923 8386
rect 10871 8117 10874 8169
rect 10874 8117 10920 8169
rect 10920 8117 10923 8169
rect 10871 7899 10874 7951
rect 10874 7899 10920 7951
rect 10920 7899 10923 7951
rect 10871 7682 10874 7734
rect 10874 7682 10920 7734
rect 10920 7682 10923 7734
rect 10871 7464 10874 7516
rect 10874 7464 10920 7516
rect 10920 7464 10923 7516
rect 10871 7246 10874 7298
rect 10874 7246 10920 7298
rect 10920 7246 10923 7298
rect 10871 7028 10874 7080
rect 10874 7028 10920 7080
rect 10920 7028 10923 7080
rect 10871 6811 10874 6863
rect 10874 6811 10920 6863
rect 10920 6811 10923 6863
rect 10871 6593 10874 6645
rect 10874 6593 10920 6645
rect 10920 6593 10923 6645
rect 10871 6376 10874 6428
rect 10874 6376 10920 6428
rect 10920 6376 10923 6428
rect 10647 6215 10650 6267
rect 10650 6215 10696 6267
rect 10696 6215 10699 6267
rect 10647 5998 10650 6050
rect 10650 5998 10696 6050
rect 10696 5998 10699 6050
rect 10647 5780 10650 5832
rect 10650 5780 10696 5832
rect 10696 5780 10699 5832
rect 10647 5562 10650 5614
rect 10650 5562 10696 5614
rect 10696 5562 10699 5614
rect 10647 5345 10650 5397
rect 10650 5345 10696 5397
rect 10696 5345 10699 5397
rect 10647 5127 10650 5179
rect 10650 5127 10696 5179
rect 10696 5127 10699 5179
rect 10647 4909 10650 4961
rect 10650 4909 10696 4961
rect 10696 4909 10699 4961
rect 8981 4431 9033 4483
rect 9193 4431 9245 4483
rect 9454 4465 9506 4517
rect 5362 3557 5414 3558
rect 5362 3511 5391 3557
rect 5391 3511 5414 3557
rect 5362 3506 5414 3511
rect 5574 3506 5626 3558
rect 2526 2678 2578 2730
rect 2658 2678 2710 2730
rect 2790 2678 2842 2730
rect 2922 2678 2974 2730
rect 3054 2678 3106 2730
rect 3186 2678 3238 2730
rect 3318 2678 3370 2730
rect 3450 2678 3502 2730
rect 3582 2678 3634 2730
rect 3714 2678 3766 2730
rect 3846 2719 3898 2730
rect 3978 2719 4030 2730
rect 4110 2719 4162 2730
rect 4242 2719 4294 2730
rect 4374 2719 4426 2730
rect 4506 2719 4558 2730
rect 4638 2719 4690 2730
rect 4770 2719 4822 2730
rect 4902 2719 4954 2730
rect 5034 2719 5086 2730
rect 5166 2719 5218 2730
rect 5298 2719 5350 2730
rect 3846 2678 3896 2719
rect 3896 2678 3898 2719
rect 3978 2678 4020 2719
rect 4020 2678 4030 2719
rect 4110 2678 4144 2719
rect 4144 2678 4162 2719
rect 4242 2678 4268 2719
rect 4268 2678 4294 2719
rect 4374 2678 4392 2719
rect 4392 2678 4426 2719
rect 4506 2678 4516 2719
rect 4516 2678 4558 2719
rect 4638 2678 4640 2719
rect 4640 2678 4686 2719
rect 4686 2678 4690 2719
rect 4770 2678 4810 2719
rect 4810 2678 4822 2719
rect 4902 2678 4934 2719
rect 4934 2678 4954 2719
rect 5034 2678 5058 2719
rect 5058 2678 5086 2719
rect 5166 2678 5182 2719
rect 5182 2678 5218 2719
rect 5298 2678 5306 2719
rect 5306 2678 5350 2719
rect 5430 2678 5482 2730
rect 5562 2678 5614 2730
rect 5694 2678 5746 2730
rect 5826 2678 5878 2730
rect 5958 2719 6010 2730
rect 6090 2719 6142 2730
rect 6222 2719 6274 2730
rect 6354 2719 6406 2730
rect 6486 2719 6538 2730
rect 6618 2719 6670 2730
rect 6750 2719 6802 2730
rect 6882 2719 6934 2730
rect 7014 2719 7066 2730
rect 7146 2719 7198 2730
rect 7278 2719 7330 2730
rect 7410 2719 7462 2730
rect 5958 2678 6004 2719
rect 6004 2678 6010 2719
rect 6090 2678 6128 2719
rect 6128 2678 6142 2719
rect 6222 2678 6252 2719
rect 6252 2678 6274 2719
rect 6354 2678 6376 2719
rect 6376 2678 6406 2719
rect 6486 2678 6500 2719
rect 6500 2678 6538 2719
rect 6618 2678 6624 2719
rect 6624 2678 6670 2719
rect 6750 2678 6794 2719
rect 6794 2678 6802 2719
rect 6882 2678 6918 2719
rect 6918 2678 6934 2719
rect 7014 2678 7042 2719
rect 7042 2678 7066 2719
rect 7146 2678 7166 2719
rect 7166 2678 7198 2719
rect 7278 2678 7290 2719
rect 7290 2678 7330 2719
rect 7410 2678 7414 2719
rect 7414 2678 7462 2719
rect 7542 2678 7594 2730
rect 2526 2546 2578 2598
rect 2658 2546 2710 2598
rect 2790 2546 2842 2598
rect 2922 2546 2974 2598
rect 3054 2546 3106 2598
rect 3186 2546 3238 2598
rect 3318 2546 3370 2598
rect 3450 2546 3502 2598
rect 3582 2546 3634 2598
rect 3714 2546 3766 2598
rect 3846 2595 3898 2598
rect 3978 2595 4030 2598
rect 4110 2595 4162 2598
rect 4242 2595 4294 2598
rect 4374 2595 4426 2598
rect 4506 2595 4558 2598
rect 4638 2595 4690 2598
rect 4770 2595 4822 2598
rect 4902 2595 4954 2598
rect 5034 2595 5086 2598
rect 5166 2595 5218 2598
rect 5298 2595 5350 2598
rect 3846 2549 3896 2595
rect 3896 2549 3898 2595
rect 3978 2549 4020 2595
rect 4020 2549 4030 2595
rect 4110 2549 4144 2595
rect 4144 2549 4162 2595
rect 4242 2549 4268 2595
rect 4268 2549 4294 2595
rect 4374 2549 4392 2595
rect 4392 2549 4426 2595
rect 4506 2549 4516 2595
rect 4516 2549 4558 2595
rect 4638 2549 4640 2595
rect 4640 2549 4686 2595
rect 4686 2549 4690 2595
rect 4770 2549 4810 2595
rect 4810 2549 4822 2595
rect 4902 2549 4934 2595
rect 4934 2549 4954 2595
rect 5034 2549 5058 2595
rect 5058 2549 5086 2595
rect 5166 2549 5182 2595
rect 5182 2549 5218 2595
rect 5298 2549 5306 2595
rect 5306 2549 5350 2595
rect 3846 2546 3898 2549
rect 3978 2546 4030 2549
rect 4110 2546 4162 2549
rect 4242 2546 4294 2549
rect 4374 2546 4426 2549
rect 4506 2546 4558 2549
rect 4638 2546 4690 2549
rect 4770 2546 4822 2549
rect 4902 2546 4954 2549
rect 5034 2546 5086 2549
rect 5166 2546 5218 2549
rect 5298 2546 5350 2549
rect 5430 2546 5482 2598
rect 5562 2546 5614 2598
rect 5694 2546 5746 2598
rect 5826 2546 5878 2598
rect 5958 2595 6010 2598
rect 6090 2595 6142 2598
rect 6222 2595 6274 2598
rect 6354 2595 6406 2598
rect 6486 2595 6538 2598
rect 6618 2595 6670 2598
rect 6750 2595 6802 2598
rect 6882 2595 6934 2598
rect 7014 2595 7066 2598
rect 7146 2595 7198 2598
rect 7278 2595 7330 2598
rect 7410 2595 7462 2598
rect 5958 2549 6004 2595
rect 6004 2549 6010 2595
rect 6090 2549 6128 2595
rect 6128 2549 6142 2595
rect 6222 2549 6252 2595
rect 6252 2549 6274 2595
rect 6354 2549 6376 2595
rect 6376 2549 6406 2595
rect 6486 2549 6500 2595
rect 6500 2549 6538 2595
rect 6618 2549 6624 2595
rect 6624 2549 6670 2595
rect 6750 2549 6794 2595
rect 6794 2549 6802 2595
rect 6882 2549 6918 2595
rect 6918 2549 6934 2595
rect 7014 2549 7042 2595
rect 7042 2549 7066 2595
rect 7146 2549 7166 2595
rect 7166 2549 7198 2595
rect 7278 2549 7290 2595
rect 7290 2549 7330 2595
rect 7410 2549 7414 2595
rect 7414 2549 7462 2595
rect 5958 2546 6010 2549
rect 6090 2546 6142 2549
rect 6222 2546 6274 2549
rect 6354 2546 6406 2549
rect 6486 2546 6538 2549
rect 6618 2546 6670 2549
rect 6750 2546 6802 2549
rect 6882 2546 6934 2549
rect 7014 2546 7066 2549
rect 7146 2546 7198 2549
rect 7278 2546 7330 2549
rect 7410 2546 7462 2549
rect 7542 2546 7594 2598
rect 8036 3019 8088 3063
rect 8036 2973 8039 3019
rect 8039 2973 8085 3019
rect 8085 2973 8088 3019
rect 8036 2905 8088 2973
rect 8036 2859 8039 2905
rect 8039 2859 8085 2905
rect 8085 2859 8088 2905
rect 8036 2791 8088 2859
rect 8036 2745 8039 2791
rect 8039 2745 8085 2791
rect 8085 2745 8088 2791
rect 8036 2699 8088 2745
rect 8981 4213 9033 4265
rect 9193 4213 9245 4265
rect 9454 4249 9506 4299
rect 9454 4247 9497 4249
rect 9497 4247 9506 4249
rect 8981 3995 9033 4047
rect 9193 3995 9245 4047
rect 9454 4035 9497 4081
rect 9497 4035 9506 4081
rect 9454 4029 9506 4035
rect 9454 3812 9506 3864
rect 9454 3594 9506 3646
rect 9454 3410 9506 3429
rect 9454 3377 9497 3410
rect 9497 3377 9506 3410
rect 8484 3019 8536 3063
rect 8484 2973 8487 3019
rect 8487 2973 8533 3019
rect 8533 2973 8536 3019
rect 8484 2905 8536 2973
rect 8484 2859 8487 2905
rect 8487 2859 8533 2905
rect 8533 2859 8536 2905
rect 8484 2791 8536 2859
rect 8484 2745 8487 2791
rect 8487 2745 8533 2791
rect 8533 2745 8536 2791
rect 8484 2699 8536 2745
rect 9454 3196 9497 3211
rect 9497 3196 9506 3211
rect 9454 3159 9506 3196
rect 9454 2941 9506 2993
rect 9454 2735 9506 2776
rect 9454 2724 9497 2735
rect 9497 2724 9506 2735
rect 9454 2519 9497 2558
rect 9497 2519 9506 2558
rect 9454 2506 9506 2519
rect 2526 2414 2578 2466
rect 2658 2414 2710 2466
rect 2790 2414 2842 2466
rect 2922 2414 2974 2466
rect 3054 2414 3106 2466
rect 3186 2414 3238 2466
rect 3318 2414 3370 2466
rect 3450 2414 3502 2466
rect 3582 2414 3634 2466
rect 3714 2414 3766 2466
rect 3846 2425 3896 2466
rect 3896 2425 3898 2466
rect 3978 2425 4020 2466
rect 4020 2425 4030 2466
rect 4110 2425 4144 2466
rect 4144 2425 4162 2466
rect 4242 2425 4268 2466
rect 4268 2425 4294 2466
rect 4374 2425 4392 2466
rect 4392 2425 4426 2466
rect 4506 2425 4516 2466
rect 4516 2425 4558 2466
rect 4638 2425 4640 2466
rect 4640 2425 4686 2466
rect 4686 2425 4690 2466
rect 4770 2425 4810 2466
rect 4810 2425 4822 2466
rect 4902 2425 4934 2466
rect 4934 2425 4954 2466
rect 5034 2425 5058 2466
rect 5058 2425 5086 2466
rect 5166 2425 5182 2466
rect 5182 2425 5218 2466
rect 5298 2425 5306 2466
rect 5306 2425 5350 2466
rect 3846 2414 3898 2425
rect 3978 2414 4030 2425
rect 4110 2414 4162 2425
rect 4242 2414 4294 2425
rect 4374 2414 4426 2425
rect 4506 2414 4558 2425
rect 4638 2414 4690 2425
rect 4770 2414 4822 2425
rect 4902 2414 4954 2425
rect 5034 2414 5086 2425
rect 5166 2414 5218 2425
rect 5298 2414 5350 2425
rect 5430 2414 5482 2466
rect 5562 2414 5614 2466
rect 5694 2414 5746 2466
rect 5826 2414 5878 2466
rect 5958 2425 6004 2466
rect 6004 2425 6010 2466
rect 6090 2425 6128 2466
rect 6128 2425 6142 2466
rect 6222 2425 6252 2466
rect 6252 2425 6274 2466
rect 6354 2425 6376 2466
rect 6376 2425 6406 2466
rect 6486 2425 6500 2466
rect 6500 2425 6538 2466
rect 6618 2425 6624 2466
rect 6624 2425 6670 2466
rect 6750 2425 6794 2466
rect 6794 2425 6802 2466
rect 6882 2425 6918 2466
rect 6918 2425 6934 2466
rect 7014 2425 7042 2466
rect 7042 2425 7066 2466
rect 7146 2425 7166 2466
rect 7166 2425 7198 2466
rect 7278 2425 7290 2466
rect 7290 2425 7330 2466
rect 7410 2425 7414 2466
rect 7414 2425 7462 2466
rect 5958 2414 6010 2425
rect 6090 2414 6142 2425
rect 6222 2414 6274 2425
rect 6354 2414 6406 2425
rect 6486 2414 6538 2425
rect 6618 2414 6670 2425
rect 6750 2414 6802 2425
rect 6882 2414 6934 2425
rect 7014 2414 7066 2425
rect 7146 2414 7198 2425
rect 7278 2414 7330 2425
rect 7410 2414 7462 2425
rect 7542 2414 7594 2466
rect 2526 2282 2578 2334
rect 2658 2282 2710 2334
rect 2790 2282 2842 2334
rect 2922 2282 2974 2334
rect 3054 2282 3106 2334
rect 3186 2282 3238 2334
rect 3318 2282 3370 2334
rect 3450 2282 3502 2334
rect 3582 2282 3634 2334
rect 3714 2282 3766 2334
rect 3846 2301 3896 2334
rect 3896 2301 3898 2334
rect 3978 2301 4020 2334
rect 4020 2301 4030 2334
rect 4110 2301 4144 2334
rect 4144 2301 4162 2334
rect 4242 2301 4268 2334
rect 4268 2301 4294 2334
rect 4374 2301 4392 2334
rect 4392 2301 4426 2334
rect 4506 2301 4516 2334
rect 4516 2301 4558 2334
rect 4638 2301 4640 2334
rect 4640 2301 4686 2334
rect 4686 2301 4690 2334
rect 4770 2301 4810 2334
rect 4810 2301 4822 2334
rect 4902 2301 4934 2334
rect 4934 2301 4954 2334
rect 5034 2301 5058 2334
rect 5058 2301 5086 2334
rect 5166 2301 5182 2334
rect 5182 2301 5218 2334
rect 5298 2301 5306 2334
rect 5306 2301 5350 2334
rect 3846 2282 3898 2301
rect 3978 2282 4030 2301
rect 4110 2282 4162 2301
rect 4242 2282 4294 2301
rect 4374 2282 4426 2301
rect 4506 2282 4558 2301
rect 4638 2282 4690 2301
rect 4770 2282 4822 2301
rect 4902 2282 4954 2301
rect 5034 2282 5086 2301
rect 5166 2282 5218 2301
rect 5298 2282 5350 2301
rect 5430 2282 5482 2334
rect 5562 2282 5614 2334
rect 5694 2282 5746 2334
rect 5826 2282 5878 2334
rect 5958 2301 6004 2334
rect 6004 2301 6010 2334
rect 6090 2301 6128 2334
rect 6128 2301 6142 2334
rect 6222 2301 6252 2334
rect 6252 2301 6274 2334
rect 6354 2301 6376 2334
rect 6376 2301 6406 2334
rect 6486 2301 6500 2334
rect 6500 2301 6538 2334
rect 6618 2301 6624 2334
rect 6624 2301 6670 2334
rect 6750 2301 6794 2334
rect 6794 2301 6802 2334
rect 6882 2301 6918 2334
rect 6918 2301 6934 2334
rect 7014 2301 7042 2334
rect 7042 2301 7066 2334
rect 7146 2301 7166 2334
rect 7166 2301 7198 2334
rect 7278 2301 7290 2334
rect 7290 2301 7330 2334
rect 7410 2301 7414 2334
rect 7414 2301 7462 2334
rect 5958 2282 6010 2301
rect 6090 2282 6142 2301
rect 6222 2282 6274 2301
rect 6354 2282 6406 2301
rect 6486 2282 6538 2301
rect 6618 2282 6670 2301
rect 6750 2282 6802 2301
rect 6882 2282 6934 2301
rect 7014 2282 7066 2301
rect 7146 2282 7198 2301
rect 7278 2282 7330 2301
rect 7410 2282 7462 2301
rect 7542 2282 7594 2334
rect 9454 2288 9506 2340
rect 9454 2071 9506 2123
rect 9454 1884 9506 1905
rect 9454 1853 9497 1884
rect 9497 1853 9506 1884
rect 9454 1668 9497 1687
rect 9497 1668 9506 1687
rect 9454 1635 9506 1668
rect 9454 1418 9506 1470
rect 9454 1204 9506 1252
rect 9454 1200 9497 1204
rect 9497 1200 9506 1204
rect 9454 1034 9506 1035
rect 9454 988 9497 1034
rect 9497 988 9506 1034
rect 9454 983 9506 988
rect 9454 765 9506 817
rect 9454 547 9506 599
rect 9454 354 9506 382
rect 9454 330 9497 354
rect 9497 330 9506 354
rect 11095 8392 11098 8444
rect 11098 8392 11144 8444
rect 11144 8392 11147 8444
rect 11095 8174 11098 8226
rect 11098 8174 11144 8226
rect 11144 8174 11147 8226
rect 11095 7956 11098 8008
rect 11098 7956 11144 8008
rect 11144 7956 11147 8008
rect 11095 7739 11098 7791
rect 11098 7739 11144 7791
rect 11144 7739 11147 7791
rect 11095 7521 11098 7573
rect 11098 7521 11144 7573
rect 11144 7521 11147 7573
rect 11095 7304 11098 7356
rect 11098 7304 11144 7356
rect 11144 7304 11147 7356
rect 11095 7086 11098 7138
rect 11098 7086 11144 7138
rect 11144 7086 11147 7138
rect 11095 6868 11098 6920
rect 11098 6868 11144 6920
rect 11144 6868 11147 6920
rect 11095 6650 11098 6702
rect 11098 6650 11144 6702
rect 11144 6650 11147 6702
rect 11095 6433 11098 6485
rect 11098 6433 11144 6485
rect 11144 6433 11147 6485
rect 11543 9045 11546 9097
rect 11546 9045 11592 9097
rect 11592 9045 11595 9097
rect 11543 8827 11546 8879
rect 11546 8827 11592 8879
rect 11592 8827 11595 8879
rect 11543 8609 11546 8661
rect 11546 8609 11592 8661
rect 11592 8609 11595 8661
rect 11319 8334 11322 8386
rect 11322 8334 11368 8386
rect 11368 8334 11371 8386
rect 11319 8117 11322 8169
rect 11322 8117 11368 8169
rect 11368 8117 11371 8169
rect 11319 7899 11322 7951
rect 11322 7899 11368 7951
rect 11368 7899 11371 7951
rect 11319 7682 11322 7734
rect 11322 7682 11368 7734
rect 11368 7682 11371 7734
rect 11319 7464 11322 7516
rect 11322 7464 11368 7516
rect 11368 7464 11371 7516
rect 11319 7246 11322 7298
rect 11322 7246 11368 7298
rect 11368 7246 11371 7298
rect 11319 7028 11322 7080
rect 11322 7028 11368 7080
rect 11368 7028 11371 7080
rect 11319 6811 11322 6863
rect 11322 6811 11368 6863
rect 11368 6811 11371 6863
rect 11319 6593 11322 6645
rect 11322 6593 11368 6645
rect 11368 6593 11371 6645
rect 11319 6376 11322 6428
rect 11322 6376 11368 6428
rect 11368 6376 11371 6428
rect 11095 6215 11098 6267
rect 11098 6215 11144 6267
rect 11144 6215 11147 6267
rect 11095 5998 11098 6050
rect 11098 5998 11144 6050
rect 11144 5998 11147 6050
rect 11095 5780 11098 5832
rect 11098 5780 11144 5832
rect 11144 5780 11147 5832
rect 11095 5562 11098 5614
rect 11098 5562 11144 5614
rect 11144 5562 11147 5614
rect 11095 5345 11098 5397
rect 11098 5345 11144 5397
rect 11144 5345 11147 5397
rect 11095 5127 11098 5179
rect 11098 5127 11144 5179
rect 11144 5127 11147 5179
rect 11095 4909 11098 4961
rect 11098 4909 11144 4961
rect 11144 4909 11147 4961
rect 11543 8392 11546 8444
rect 11546 8392 11592 8444
rect 11592 8392 11595 8444
rect 11543 8174 11546 8226
rect 11546 8174 11592 8226
rect 11592 8174 11595 8226
rect 11543 7956 11546 8008
rect 11546 7956 11592 8008
rect 11592 7956 11595 8008
rect 11543 7739 11546 7791
rect 11546 7739 11592 7791
rect 11592 7739 11595 7791
rect 11543 7521 11546 7573
rect 11546 7521 11592 7573
rect 11592 7521 11595 7573
rect 11543 7304 11546 7356
rect 11546 7304 11592 7356
rect 11592 7304 11595 7356
rect 11543 7086 11546 7138
rect 11546 7086 11592 7138
rect 11592 7086 11595 7138
rect 11543 6868 11546 6920
rect 11546 6868 11592 6920
rect 11592 6868 11595 6920
rect 11543 6650 11546 6702
rect 11546 6650 11592 6702
rect 11592 6650 11595 6702
rect 11543 6433 11546 6485
rect 11546 6433 11592 6485
rect 11592 6433 11595 6485
rect 11543 6215 11546 6267
rect 11546 6215 11592 6267
rect 11592 6215 11595 6267
rect 11543 5998 11546 6050
rect 11546 5998 11592 6050
rect 11592 5998 11595 6050
rect 11543 5780 11546 5832
rect 11546 5780 11592 5832
rect 11592 5780 11595 5832
rect 11543 5562 11546 5614
rect 11546 5562 11592 5614
rect 11592 5562 11595 5614
rect 11543 5345 11546 5397
rect 11546 5345 11592 5397
rect 11592 5345 11595 5397
rect 11543 5127 11546 5179
rect 11546 5127 11592 5179
rect 11592 5127 11595 5179
rect 11543 4909 11546 4961
rect 11546 4909 11592 4961
rect 11592 4909 11595 4961
rect 12153 8348 12159 8400
rect 12159 8348 12205 8400
rect 12153 8131 12159 8183
rect 12159 8131 12205 8183
rect 12153 7913 12159 7965
rect 12159 7913 12205 7965
rect 12153 7696 12159 7748
rect 12159 7696 12205 7748
rect 12153 7478 12159 7530
rect 12159 7478 12205 7530
rect 12153 7260 12159 7312
rect 12159 7260 12205 7312
rect 12153 7042 12159 7094
rect 12159 7042 12205 7094
rect 12153 6825 12159 6877
rect 12159 6825 12205 6877
rect 12153 6607 12159 6659
rect 12159 6607 12205 6659
rect 12153 6390 12159 6442
rect 12159 6390 12205 6442
rect 11931 5361 11935 5413
rect 11935 5361 11981 5413
rect 11981 5361 11983 5413
rect 11931 5143 11935 5195
rect 11935 5143 11981 5195
rect 11981 5143 11983 5195
rect 11931 4925 11935 4977
rect 11935 4925 11981 4977
rect 11981 4925 11983 4977
rect 11931 4707 11935 4759
rect 11935 4707 11981 4759
rect 11981 4707 11983 4759
rect 12601 8348 12607 8400
rect 12607 8348 12653 8400
rect 12601 8131 12607 8183
rect 12607 8131 12653 8183
rect 12601 7913 12607 7965
rect 12607 7913 12653 7965
rect 12601 7696 12607 7748
rect 12607 7696 12653 7748
rect 12601 7478 12607 7530
rect 12607 7478 12653 7530
rect 12601 7260 12607 7312
rect 12607 7260 12653 7312
rect 12601 7042 12607 7094
rect 12607 7042 12653 7094
rect 12601 6825 12607 6877
rect 12607 6825 12653 6877
rect 12601 6607 12607 6659
rect 12607 6607 12653 6659
rect 12601 6390 12607 6442
rect 12607 6390 12653 6442
rect 12379 5361 12383 5413
rect 12383 5361 12429 5413
rect 12429 5361 12431 5413
rect 12379 5143 12383 5195
rect 12383 5143 12429 5195
rect 12429 5143 12431 5195
rect 12379 4925 12383 4977
rect 12383 4925 12429 4977
rect 12429 4925 12431 4977
rect 12379 4707 12383 4759
rect 12383 4707 12429 4759
rect 12429 4707 12431 4759
rect 13400 8353 13452 8400
rect 13400 8348 13410 8353
rect 13410 8348 13452 8353
rect 13400 8144 13410 8183
rect 13410 8144 13452 8183
rect 13400 8131 13452 8144
rect 13400 7913 13452 7965
rect 13400 7700 13452 7748
rect 13400 7696 13410 7700
rect 13410 7696 13452 7700
rect 13400 7491 13410 7530
rect 13410 7491 13452 7530
rect 13400 7478 13452 7491
rect 13400 7260 13452 7312
rect 13400 7047 13452 7094
rect 13400 7042 13410 7047
rect 13410 7042 13452 7047
rect 13400 6837 13410 6877
rect 13410 6837 13452 6877
rect 13400 6825 13452 6837
rect 13400 6607 13452 6659
rect 13400 6394 13452 6442
rect 13400 6390 13410 6394
rect 13410 6390 13452 6394
rect 12827 5361 12831 5413
rect 12831 5361 12877 5413
rect 12877 5361 12879 5413
rect 12827 5143 12831 5195
rect 12831 5143 12877 5195
rect 12877 5143 12879 5195
rect 12827 4925 12831 4977
rect 12831 4925 12877 4977
rect 12877 4925 12879 4977
rect 12827 4707 12831 4759
rect 12831 4707 12877 4759
rect 12877 4707 12879 4759
rect 12633 4460 12685 4512
rect 12845 4460 12897 4512
rect 11595 4238 11647 4290
rect 11807 4238 11859 4290
rect 10647 3939 10699 3991
rect 10647 3732 10699 3773
rect 10647 3721 10650 3732
rect 10650 3721 10696 3732
rect 10696 3721 10699 3732
rect 10647 3518 10650 3556
rect 10650 3518 10696 3556
rect 10696 3518 10699 3556
rect 10647 3504 10699 3518
rect 10647 3286 10699 3338
rect 10647 3068 10699 3120
rect 10647 2893 10699 2903
rect 10647 2851 10650 2893
rect 10650 2851 10696 2893
rect 10696 2851 10699 2893
rect 10647 2680 10650 2685
rect 10650 2680 10696 2685
rect 10696 2680 10699 2685
rect 10647 2633 10699 2680
rect 10647 2416 10699 2468
rect 10647 2220 10699 2250
rect 10647 2198 10650 2220
rect 10650 2198 10696 2220
rect 10696 2198 10699 2220
rect 11095 4022 11098 4064
rect 11098 4022 11144 4064
rect 11144 4022 11147 4064
rect 11095 4012 11147 4022
rect 11095 3794 11147 3846
rect 11095 3576 11147 3628
rect 11095 3397 11147 3411
rect 11095 3359 11098 3397
rect 11098 3359 11144 3397
rect 11144 3359 11147 3397
rect 11095 3183 11098 3193
rect 11098 3183 11144 3193
rect 11144 3183 11147 3193
rect 11095 3141 11147 3183
rect 11095 2923 11147 2975
rect 11095 2726 11147 2758
rect 11095 2706 11098 2726
rect 11098 2706 11144 2726
rect 11144 2706 11147 2726
rect 11095 2512 11098 2540
rect 11098 2512 11144 2540
rect 11144 2512 11147 2540
rect 11095 2488 11147 2512
rect 11095 2270 11147 2322
rect 11543 3939 11595 3991
rect 11543 3732 11595 3773
rect 11543 3721 11546 3732
rect 11546 3721 11592 3732
rect 11592 3721 11595 3732
rect 11543 3518 11546 3556
rect 11546 3518 11592 3556
rect 11592 3518 11595 3556
rect 11543 3504 11595 3518
rect 11543 3286 11595 3338
rect 11543 3068 11595 3120
rect 11543 2893 11595 2903
rect 11543 2851 11546 2893
rect 11546 2851 11592 2893
rect 11592 2851 11595 2893
rect 11543 2680 11546 2685
rect 11546 2680 11592 2685
rect 11592 2680 11595 2685
rect 11543 2633 11595 2680
rect 11543 2416 11595 2468
rect 10647 2004 10650 2032
rect 10650 2004 10696 2032
rect 10696 2004 10699 2032
rect 10647 1980 10699 2004
rect 10647 1762 10699 1814
rect 10647 1545 10699 1597
rect 10647 1370 10699 1379
rect 10647 1327 10650 1370
rect 10650 1327 10696 1370
rect 10696 1327 10699 1370
rect 10647 1154 10650 1162
rect 10650 1154 10696 1162
rect 10696 1154 10699 1162
rect 10647 1110 10699 1154
rect 10647 892 10699 944
rect 10647 690 10699 726
rect 10647 674 10650 690
rect 10650 674 10696 690
rect 10696 674 10699 690
rect 10647 457 10699 509
rect 11543 2220 11595 2250
rect 11543 2198 11546 2220
rect 11546 2198 11592 2220
rect 11592 2198 11595 2220
rect 11543 2004 11546 2032
rect 11546 2004 11592 2032
rect 11592 2004 11595 2032
rect 11543 1980 11595 2004
rect 11543 1762 11595 1814
rect 11543 1545 11595 1597
rect 11543 1370 11595 1379
rect 11543 1327 11546 1370
rect 11546 1327 11592 1370
rect 11592 1327 11595 1370
rect 11543 1154 11546 1162
rect 11546 1154 11592 1162
rect 11592 1154 11595 1162
rect 11543 1110 11595 1154
rect 11543 892 11595 944
rect 11543 690 11595 726
rect 11543 674 11546 690
rect 11546 674 11592 690
rect 11592 674 11595 690
rect 10647 239 10699 291
rect 11543 457 11595 509
rect 11543 239 11595 291
rect 11931 3939 11983 3991
rect 11931 3732 11983 3773
rect 11931 3721 11934 3732
rect 11934 3721 11980 3732
rect 11980 3721 11983 3732
rect 11931 3518 11934 3556
rect 11934 3518 11980 3556
rect 11980 3518 11983 3556
rect 11931 3504 11983 3518
rect 11931 3286 11983 3338
rect 11931 3068 11983 3120
rect 11931 2851 11983 2903
rect 11931 2633 11983 2685
rect 11931 2416 11983 2468
rect 11931 2198 11983 2250
rect 12379 4022 12382 4064
rect 12382 4022 12428 4064
rect 12428 4022 12431 4064
rect 12379 4012 12431 4022
rect 12379 3794 12431 3846
rect 12379 3576 12431 3628
rect 12379 3397 12431 3411
rect 12379 3359 12382 3397
rect 12382 3359 12428 3397
rect 12428 3359 12431 3397
rect 12379 3141 12431 3193
rect 12379 2923 12431 2975
rect 12379 2706 12431 2758
rect 12379 2488 12431 2540
rect 12379 2270 12431 2322
rect 12827 3939 12879 3991
rect 13515 3939 13567 3991
rect 12827 3732 12879 3773
rect 13515 3742 13567 3773
rect 12827 3721 12830 3732
rect 12830 3721 12876 3732
rect 12876 3721 12879 3732
rect 13515 3721 13557 3742
rect 13557 3721 13567 3742
rect 12827 3518 12830 3556
rect 12830 3518 12876 3556
rect 12876 3518 12879 3556
rect 13515 3532 13557 3556
rect 13557 3532 13567 3556
rect 12827 3504 12879 3518
rect 13515 3504 13567 3532
rect 12827 3286 12879 3338
rect 13515 3286 13567 3338
rect 12827 3068 12879 3120
rect 13515 3089 13567 3120
rect 13515 3068 13557 3089
rect 13557 3068 13567 3089
rect 12827 2851 12879 2903
rect 13515 2879 13557 2903
rect 13557 2879 13567 2903
rect 13515 2851 13567 2879
rect 12827 2633 12879 2685
rect 13515 2633 13567 2685
rect 12827 2416 12879 2468
rect 13515 2436 13567 2468
rect 13515 2416 13557 2436
rect 13557 2416 13567 2436
rect 11931 1980 11983 2032
rect 11931 1762 11983 1814
rect 11931 1545 11983 1597
rect 11931 1327 11983 1379
rect 11931 1110 11983 1162
rect 11931 892 11983 944
rect 11931 674 11983 726
rect 11931 457 11983 509
rect 11931 239 11983 291
rect 12827 2198 12879 2250
rect 13515 2226 13557 2250
rect 13557 2226 13567 2250
rect 13515 2198 13567 2226
rect 12827 1980 12879 2032
rect 13515 1980 13567 2032
rect 12827 1762 12879 1814
rect 13515 1782 13567 1814
rect 13515 1762 13557 1782
rect 13557 1762 13567 1782
rect 12827 1545 12879 1597
rect 13515 1573 13557 1597
rect 13557 1573 13567 1597
rect 13515 1545 13567 1573
rect 12827 1327 12879 1379
rect 13515 1327 13567 1379
rect 12827 1110 12879 1162
rect 13515 1129 13567 1162
rect 13515 1110 13557 1129
rect 13557 1110 13567 1129
rect 12827 892 12879 944
rect 13515 920 13557 944
rect 13557 920 13567 944
rect 13515 892 13567 920
rect 12827 674 12879 726
rect 13515 674 13567 726
rect 12827 457 12879 509
rect 13515 476 13567 509
rect 13515 457 13557 476
rect 13557 457 13567 476
rect 12827 239 12879 291
rect 13515 267 13557 291
rect 13557 267 13567 291
rect 13515 239 13567 267
rect 10253 -529 10305 -477
rect 10465 -529 10517 -477
rect 12976 -529 13028 -477
rect 13188 -529 13240 -477
rect 10253 -747 10305 -695
rect 10465 -747 10517 -695
rect 12976 -747 13028 -695
rect 13188 -747 13240 -695
<< metal2 >>
rect 6225 16240 13430 16278
rect 6225 16184 6327 16240
rect 6383 16184 6775 16240
rect 6831 16184 7223 16240
rect 7279 16184 7671 16240
rect 7727 16184 8119 16240
rect 8175 16184 8567 16240
rect 8623 16184 8857 16240
rect 8913 16184 9305 16240
rect 9361 16184 9753 16240
rect 9809 16184 10201 16240
rect 10257 16184 10649 16240
rect 10705 16184 11097 16240
rect 11153 16184 11545 16240
rect 11601 16184 11993 16240
rect 12049 16184 12441 16240
rect 12497 16184 12889 16240
rect 12945 16184 13337 16240
rect 13393 16184 13430 16240
rect 6225 16022 13430 16184
rect 6225 15966 6327 16022
rect 6383 15966 6775 16022
rect 6831 15966 7223 16022
rect 7279 15966 7671 16022
rect 7727 15966 8119 16022
rect 8175 15966 8567 16022
rect 8623 15966 8857 16022
rect 8913 15966 9305 16022
rect 9361 15966 9753 16022
rect 9809 15966 10201 16022
rect 10257 15966 10649 16022
rect 10705 15966 11097 16022
rect 11153 15966 11545 16022
rect 11601 15966 11993 16022
rect 12049 15966 12441 16022
rect 12497 15966 12889 16022
rect 12945 15966 13337 16022
rect 13393 15966 13430 16022
rect 6225 15805 13430 15966
rect 6225 15749 6327 15805
rect 6383 15749 6775 15805
rect 6831 15749 7223 15805
rect 7279 15749 7671 15805
rect 7727 15749 8119 15805
rect 8175 15749 8567 15805
rect 8623 15749 8857 15805
rect 8913 15749 9305 15805
rect 9361 15749 9753 15805
rect 9809 15749 10201 15805
rect 10257 15749 10649 15805
rect 10705 15749 11097 15805
rect 11153 15749 11545 15805
rect 11601 15749 11993 15805
rect 12049 15749 12441 15805
rect 12497 15749 12889 15805
rect 12945 15749 13337 15805
rect 13393 15749 13430 15805
rect 6225 15587 13430 15749
rect 6225 15531 6327 15587
rect 6383 15531 6775 15587
rect 6831 15531 7223 15587
rect 7279 15531 7671 15587
rect 7727 15531 8119 15587
rect 8175 15531 8567 15587
rect 8623 15531 8857 15587
rect 8913 15531 9305 15587
rect 9361 15531 9753 15587
rect 9809 15531 10201 15587
rect 10257 15531 10649 15587
rect 10705 15531 11097 15587
rect 11153 15531 11545 15587
rect 11601 15531 11993 15587
rect 12049 15531 12441 15587
rect 12497 15531 12889 15587
rect 12945 15531 13337 15587
rect 13393 15531 13430 15587
rect 6225 15369 13430 15531
rect 6225 15313 6327 15369
rect 6383 15313 6775 15369
rect 6831 15313 7223 15369
rect 7279 15313 7671 15369
rect 7727 15313 8119 15369
rect 8175 15313 8567 15369
rect 8623 15313 8857 15369
rect 8913 15313 9305 15369
rect 9361 15313 9753 15369
rect 9809 15313 10201 15369
rect 10257 15313 10649 15369
rect 10705 15313 11097 15369
rect 11153 15313 11545 15369
rect 11601 15313 11993 15369
rect 12049 15313 12441 15369
rect 12497 15313 12889 15369
rect 12945 15313 13337 15369
rect 13393 15313 13430 15369
rect 6225 15151 13430 15313
rect 6225 15095 6327 15151
rect 6383 15095 6775 15151
rect 6831 15095 7223 15151
rect 7279 15095 7671 15151
rect 7727 15095 8119 15151
rect 8175 15095 8567 15151
rect 8623 15095 8857 15151
rect 8913 15095 9305 15151
rect 9361 15095 9753 15151
rect 9809 15095 10201 15151
rect 10257 15095 10649 15151
rect 10705 15095 11097 15151
rect 11153 15095 11545 15151
rect 11601 15095 11993 15151
rect 12049 15095 12441 15151
rect 12497 15095 12889 15151
rect 12945 15095 13337 15151
rect 13393 15095 13430 15151
rect 6225 14934 13430 15095
rect 6225 14878 6327 14934
rect 6383 14878 6775 14934
rect 6831 14878 7223 14934
rect 7279 14878 7671 14934
rect 7727 14878 8119 14934
rect 8175 14878 8567 14934
rect 8623 14878 8857 14934
rect 8913 14878 9305 14934
rect 9361 14878 9753 14934
rect 9809 14878 10201 14934
rect 10257 14878 10649 14934
rect 10705 14878 11097 14934
rect 11153 14878 11545 14934
rect 11601 14878 11993 14934
rect 12049 14878 12441 14934
rect 12497 14878 12889 14934
rect 12945 14878 13337 14934
rect 13393 14878 13430 14934
rect 6225 14716 13430 14878
rect 6225 14660 6327 14716
rect 6383 14660 6775 14716
rect 6831 14660 7223 14716
rect 7279 14660 7671 14716
rect 7727 14660 8119 14716
rect 8175 14660 8567 14716
rect 8623 14660 8857 14716
rect 8913 14660 9305 14716
rect 9361 14660 9753 14716
rect 9809 14660 10201 14716
rect 10257 14660 10649 14716
rect 10705 14660 11097 14716
rect 11153 14660 11545 14716
rect 11601 14660 11993 14716
rect 12049 14660 12441 14716
rect 12497 14660 12889 14716
rect 12945 14660 13337 14716
rect 13393 14660 13430 14716
rect 6225 14621 13430 14660
rect 6513 14433 8434 14474
rect 6513 14381 6551 14433
rect 6603 14381 6999 14433
rect 7051 14381 7447 14433
rect 7499 14381 7895 14433
rect 7947 14381 8343 14433
rect 8395 14381 8434 14433
rect 6513 14216 8434 14381
rect 6513 14164 6551 14216
rect 6603 14164 6999 14216
rect 7051 14164 7447 14216
rect 7499 14164 7895 14216
rect 7947 14164 8343 14216
rect 8395 14164 8434 14216
rect 6513 13998 8434 14164
rect 6513 13946 6551 13998
rect 6603 13946 6999 13998
rect 7051 13946 7447 13998
rect 7499 13946 7895 13998
rect 7947 13946 8343 13998
rect 8395 13946 8434 13998
rect 6513 13780 8434 13946
rect 6513 13728 6551 13780
rect 6603 13728 6999 13780
rect 7051 13728 7447 13780
rect 7499 13728 7895 13780
rect 7947 13728 8343 13780
rect 8395 13728 8434 13780
rect 6513 13563 8434 13728
rect 6513 13511 6551 13563
rect 6603 13511 6999 13563
rect 7051 13511 7447 13563
rect 7499 13511 7895 13563
rect 7947 13511 8343 13563
rect 8395 13511 8434 13563
rect 6513 13470 8434 13511
rect 9045 14336 13206 14376
rect 9045 14284 9083 14336
rect 9135 14284 9531 14336
rect 9583 14284 9979 14336
rect 10031 14284 10427 14336
rect 10479 14284 10875 14336
rect 10927 14284 11323 14336
rect 11375 14284 11771 14336
rect 11823 14284 12219 14336
rect 12271 14284 12667 14336
rect 12719 14284 13115 14336
rect 13167 14284 13206 14336
rect 9045 14118 13206 14284
rect 9045 14066 9083 14118
rect 9135 14066 9531 14118
rect 9583 14066 9979 14118
rect 10031 14066 10427 14118
rect 10479 14066 10875 14118
rect 10927 14066 11323 14118
rect 11375 14066 11771 14118
rect 11823 14066 12219 14118
rect 12271 14066 12667 14118
rect 12719 14066 13115 14118
rect 13167 14066 13206 14118
rect 9045 13900 13206 14066
rect 9045 13848 9083 13900
rect 9135 13848 9531 13900
rect 9583 13848 9979 13900
rect 10031 13848 10427 13900
rect 10479 13848 10875 13900
rect 10927 13848 11323 13900
rect 11375 13848 11771 13900
rect 11823 13848 12219 13900
rect 12271 13848 12667 13900
rect 12719 13848 13115 13900
rect 13167 13848 13206 13900
rect 9045 13683 13206 13848
rect 9045 13631 9083 13683
rect 9135 13631 9531 13683
rect 9583 13631 9979 13683
rect 10031 13631 10427 13683
rect 10479 13631 10875 13683
rect 10927 13631 11323 13683
rect 11375 13631 11771 13683
rect 11823 13631 12219 13683
rect 12271 13631 12667 13683
rect 12719 13631 13115 13683
rect 13167 13631 13206 13683
rect 6497 13336 7364 13376
rect 6497 13284 6577 13336
rect 6629 13284 6788 13336
rect 6840 13284 7000 13336
rect 7052 13284 7211 13336
rect 7263 13284 7364 13336
rect 6276 11295 6404 11332
rect 6276 11239 6312 11295
rect 6368 11239 6404 11295
rect 6276 11077 6404 11239
rect 6276 11021 6312 11077
rect 6368 11021 6404 11077
rect 6276 10860 6404 11021
rect 6276 10804 6312 10860
rect 6368 10804 6404 10860
rect 6276 10642 6404 10804
rect 6276 10586 6312 10642
rect 6368 10586 6404 10642
rect 6276 10424 6404 10586
rect 6276 10368 6312 10424
rect 6368 10368 6404 10424
rect 6276 10207 6404 10368
rect 6276 10151 6312 10207
rect 6368 10151 6404 10207
rect 6276 9989 6404 10151
rect 6276 9933 6312 9989
rect 6368 9933 6404 9989
rect 6276 9895 6404 9933
rect 6497 11200 7364 13284
rect 6497 11148 6607 11200
rect 6659 11148 6818 11200
rect 6870 11148 7030 11200
rect 7082 11148 7241 11200
rect 7293 11148 7364 11200
rect 6497 11107 7364 11148
rect 7591 12211 8192 13470
rect 9045 13465 13206 13631
rect 9045 13413 9083 13465
rect 9135 13413 9531 13465
rect 9583 13413 9979 13465
rect 10031 13413 10427 13465
rect 10479 13413 10875 13465
rect 10927 13413 11323 13465
rect 11375 13413 11771 13465
rect 11823 13413 12219 13465
rect 12271 13413 12667 13465
rect 12719 13413 13115 13465
rect 13167 13413 13206 13465
rect 9045 13247 13206 13413
rect 9045 13195 9083 13247
rect 9135 13195 9531 13247
rect 9583 13195 9979 13247
rect 10031 13195 10427 13247
rect 10479 13195 10875 13247
rect 10927 13195 11323 13247
rect 11375 13195 11771 13247
rect 11823 13195 12219 13247
rect 12271 13195 12667 13247
rect 12719 13195 13115 13247
rect 13167 13195 13206 13247
rect 9045 13030 13206 13195
rect 9045 12978 9083 13030
rect 9135 12978 9531 13030
rect 9583 12978 9979 13030
rect 10031 12978 10427 13030
rect 10479 12978 10875 13030
rect 10927 12978 11323 13030
rect 11375 12978 11771 13030
rect 11823 12978 12219 13030
rect 12271 12978 12667 13030
rect 12719 12978 13115 13030
rect 13167 12978 13206 13030
rect 9045 12812 13206 12978
rect 9045 12760 9083 12812
rect 9135 12760 9531 12812
rect 9583 12760 9979 12812
rect 10031 12760 10427 12812
rect 10479 12760 10875 12812
rect 10927 12760 11323 12812
rect 11375 12760 11771 12812
rect 11823 12760 12219 12812
rect 12271 12760 12667 12812
rect 12719 12760 13115 12812
rect 13167 12760 13206 12812
rect 9045 12594 13206 12760
rect 9045 12542 9083 12594
rect 9135 12542 9531 12594
rect 9583 12542 9979 12594
rect 10031 12542 10427 12594
rect 10479 12542 10875 12594
rect 10927 12542 11323 12594
rect 11375 12542 11771 12594
rect 11823 12542 12219 12594
rect 12271 12542 12667 12594
rect 12719 12542 13115 12594
rect 13167 12542 13206 12594
rect 9045 12502 13206 12542
rect 7591 12170 11159 12211
rect 7591 12118 9142 12170
rect 9194 12118 9353 12170
rect 9405 12118 9564 12170
rect 9616 12118 9774 12170
rect 9826 12118 9985 12170
rect 10037 12118 10197 12170
rect 10249 12118 10408 12170
rect 10460 12118 10618 12170
rect 10670 12118 10829 12170
rect 10881 12118 11040 12170
rect 11092 12118 11159 12170
rect 7591 11477 11159 12118
rect 7591 11425 9142 11477
rect 9194 11425 9353 11477
rect 9405 11425 9564 11477
rect 9616 11425 9774 11477
rect 9826 11425 9985 11477
rect 10037 11425 10197 11477
rect 10249 11425 10408 11477
rect 10460 11425 10618 11477
rect 10670 11425 10829 11477
rect 10881 11425 11040 11477
rect 11092 11425 11159 11477
rect 7591 11384 11159 11425
rect 6497 9258 6725 11107
rect 7591 10955 8192 11384
rect 11555 11282 13206 12502
rect 6838 10954 8192 10955
rect 6808 10915 8192 10954
rect 6808 10863 6846 10915
rect 6898 10863 7293 10915
rect 7345 10863 7741 10915
rect 7793 10863 8192 10915
rect 6808 10697 8192 10863
rect 6808 10645 6846 10697
rect 6898 10656 7293 10697
rect 6898 10645 6936 10656
rect 6808 10480 6936 10645
rect 6808 10428 6846 10480
rect 6898 10428 6936 10480
rect 6808 10262 6936 10428
rect 7255 10645 7293 10656
rect 7345 10656 7741 10697
rect 7345 10645 7383 10656
rect 7255 10480 7383 10645
rect 7255 10428 7293 10480
rect 7345 10428 7383 10480
rect 6808 10210 6846 10262
rect 6898 10210 6936 10262
rect 6808 10044 6936 10210
rect 6808 9992 6846 10044
rect 6898 9992 6936 10044
rect 6808 9827 6936 9992
rect 6808 9775 6846 9827
rect 6898 9775 6936 9827
rect 6808 9609 6936 9775
rect 6808 9557 6846 9609
rect 6898 9557 6936 9609
rect 6808 9517 6936 9557
rect 7032 10264 7160 10301
rect 7032 10208 7068 10264
rect 7124 10208 7160 10264
rect 7032 10046 7160 10208
rect 7032 9990 7068 10046
rect 7124 9990 7160 10046
rect 7032 9828 7160 9990
rect 7032 9772 7068 9828
rect 7124 9772 7160 9828
rect 7032 9610 7160 9772
rect 7032 9554 7068 9610
rect 7124 9554 7160 9610
rect 7032 9516 7160 9554
rect 7255 10262 7383 10428
rect 7703 10645 7741 10656
rect 7793 10656 8192 10697
rect 8428 11195 13206 11282
rect 8428 11143 9083 11195
rect 9135 11143 9531 11195
rect 9583 11143 9979 11195
rect 10031 11143 10427 11195
rect 10479 11143 10875 11195
rect 10927 11143 11323 11195
rect 11375 11143 11771 11195
rect 11823 11143 12219 11195
rect 12271 11143 12667 11195
rect 12719 11143 13115 11195
rect 13167 11143 13206 11195
rect 8428 10978 13206 11143
rect 8428 10926 9083 10978
rect 9135 10926 9531 10978
rect 9583 10926 9979 10978
rect 10031 10926 10427 10978
rect 10479 10926 10875 10978
rect 10927 10926 11323 10978
rect 11375 10926 11771 10978
rect 11823 10926 12219 10978
rect 12271 10926 12667 10978
rect 12719 10926 13115 10978
rect 13167 10926 13206 10978
rect 8428 10760 13206 10926
rect 8428 10731 9083 10760
rect 7793 10645 7831 10656
rect 7703 10480 7831 10645
rect 7703 10428 7741 10480
rect 7793 10428 7831 10480
rect 7255 10210 7293 10262
rect 7345 10210 7383 10262
rect 7255 10044 7383 10210
rect 7255 9992 7293 10044
rect 7345 9992 7383 10044
rect 7255 9827 7383 9992
rect 7255 9775 7293 9827
rect 7345 9775 7383 9827
rect 7255 9609 7383 9775
rect 7255 9557 7293 9609
rect 7345 9557 7383 9609
rect 7255 9517 7383 9557
rect 7479 10264 7607 10301
rect 7479 10208 7515 10264
rect 7571 10208 7607 10264
rect 7479 10046 7607 10208
rect 7479 9990 7515 10046
rect 7571 9990 7607 10046
rect 7479 9828 7607 9990
rect 7479 9772 7515 9828
rect 7571 9772 7607 9828
rect 7479 9610 7607 9772
rect 7479 9554 7515 9610
rect 7571 9554 7607 9610
rect 7479 9516 7607 9554
rect 7703 10262 7831 10428
rect 7703 10210 7741 10262
rect 7793 10210 7831 10262
rect 7703 10044 7831 10210
rect 7703 9992 7741 10044
rect 7793 9992 7831 10044
rect 7703 9827 7831 9992
rect 7703 9775 7741 9827
rect 7793 9775 7831 9827
rect 7703 9609 7831 9775
rect 7703 9557 7741 9609
rect 7793 9557 7831 9609
rect 7703 9517 7831 9557
rect 7980 10476 8319 10515
rect 7980 10420 8015 10476
rect 8071 10420 8227 10476
rect 8283 10420 8319 10476
rect 7980 10259 8319 10420
rect 7980 10203 8015 10259
rect 8071 10203 8227 10259
rect 8283 10203 8319 10259
rect 7980 10041 8319 10203
rect 7980 9985 8015 10041
rect 8071 9985 8227 10041
rect 8283 9985 8319 10041
rect 7980 9823 8319 9985
rect 7980 9767 8015 9823
rect 8071 9767 8227 9823
rect 8283 9767 8319 9823
rect 7980 9606 8319 9767
rect 7980 9550 8015 9606
rect 8071 9550 8227 9606
rect 8283 9550 8319 9606
rect 7980 9511 8319 9550
rect 8428 9736 8719 10731
rect 9045 10708 9083 10731
rect 9135 10731 9531 10760
rect 9135 10708 9174 10731
rect 8823 10595 8951 10632
rect 8823 10539 8859 10595
rect 8915 10539 8951 10595
rect 8823 10377 8951 10539
rect 8823 10321 8859 10377
rect 8915 10321 8951 10377
rect 8823 10159 8951 10321
rect 8823 10103 8859 10159
rect 8915 10103 8951 10159
rect 8823 9941 8951 10103
rect 8823 9885 8859 9941
rect 8915 9885 8951 9941
rect 8823 9847 8951 9885
rect 9045 10542 9174 10708
rect 9493 10708 9531 10731
rect 9583 10731 9979 10760
rect 9583 10708 9622 10731
rect 9045 10490 9083 10542
rect 9135 10490 9174 10542
rect 9045 10324 9174 10490
rect 9045 10272 9083 10324
rect 9135 10272 9174 10324
rect 9045 10107 9174 10272
rect 9045 10055 9083 10107
rect 9135 10055 9174 10107
rect 9045 9736 9174 10055
rect 9271 10595 9399 10632
rect 9271 10539 9307 10595
rect 9363 10539 9399 10595
rect 9271 10377 9399 10539
rect 9271 10321 9307 10377
rect 9363 10321 9399 10377
rect 9271 10159 9399 10321
rect 9271 10103 9307 10159
rect 9363 10103 9399 10159
rect 9271 9941 9399 10103
rect 9271 9885 9307 9941
rect 9363 9885 9399 9941
rect 9271 9847 9399 9885
rect 9493 10542 9622 10708
rect 9941 10708 9979 10731
rect 10031 10731 10427 10760
rect 10031 10708 10070 10731
rect 9493 10490 9531 10542
rect 9583 10490 9622 10542
rect 9493 10324 9622 10490
rect 9493 10272 9531 10324
rect 9583 10272 9622 10324
rect 9493 10107 9622 10272
rect 9493 10055 9531 10107
rect 9583 10055 9622 10107
rect 9493 9736 9622 10055
rect 9719 10595 9847 10632
rect 9719 10539 9755 10595
rect 9811 10539 9847 10595
rect 9719 10377 9847 10539
rect 9719 10321 9755 10377
rect 9811 10321 9847 10377
rect 9719 10159 9847 10321
rect 9719 10103 9755 10159
rect 9811 10103 9847 10159
rect 9719 9941 9847 10103
rect 9719 9885 9755 9941
rect 9811 9885 9847 9941
rect 9719 9847 9847 9885
rect 9941 10542 10070 10708
rect 10389 10708 10427 10731
rect 10479 10731 10875 10760
rect 10479 10708 10518 10731
rect 9941 10490 9979 10542
rect 10031 10490 10070 10542
rect 9941 10324 10070 10490
rect 9941 10272 9979 10324
rect 10031 10272 10070 10324
rect 9941 10107 10070 10272
rect 9941 10055 9979 10107
rect 10031 10055 10070 10107
rect 9941 9736 10070 10055
rect 10167 10595 10295 10632
rect 10167 10539 10203 10595
rect 10259 10539 10295 10595
rect 10167 10377 10295 10539
rect 10167 10321 10203 10377
rect 10259 10321 10295 10377
rect 10167 10159 10295 10321
rect 10167 10103 10203 10159
rect 10259 10103 10295 10159
rect 10167 9941 10295 10103
rect 10167 9885 10203 9941
rect 10259 9885 10295 9941
rect 10167 9847 10295 9885
rect 10389 10542 10518 10708
rect 10837 10708 10875 10731
rect 10927 10731 11323 10760
rect 10927 10708 10966 10731
rect 10389 10490 10427 10542
rect 10479 10490 10518 10542
rect 10389 10324 10518 10490
rect 10389 10272 10427 10324
rect 10479 10272 10518 10324
rect 10389 10107 10518 10272
rect 10389 10055 10427 10107
rect 10479 10055 10518 10107
rect 10389 9736 10518 10055
rect 10615 10595 10743 10632
rect 10615 10539 10651 10595
rect 10707 10539 10743 10595
rect 10615 10377 10743 10539
rect 10615 10321 10651 10377
rect 10707 10321 10743 10377
rect 10615 10159 10743 10321
rect 10615 10103 10651 10159
rect 10707 10103 10743 10159
rect 10615 9941 10743 10103
rect 10615 9885 10651 9941
rect 10707 9885 10743 9941
rect 10615 9847 10743 9885
rect 10837 10542 10966 10708
rect 11285 10708 11323 10731
rect 11375 10731 11771 10760
rect 11375 10708 11414 10731
rect 10837 10490 10875 10542
rect 10927 10490 10966 10542
rect 10837 10324 10966 10490
rect 10837 10272 10875 10324
rect 10927 10272 10966 10324
rect 10837 10107 10966 10272
rect 10837 10055 10875 10107
rect 10927 10055 10966 10107
rect 10837 9736 10966 10055
rect 11063 10595 11191 10632
rect 11063 10539 11099 10595
rect 11155 10539 11191 10595
rect 11063 10377 11191 10539
rect 11063 10321 11099 10377
rect 11155 10321 11191 10377
rect 11063 10159 11191 10321
rect 11063 10103 11099 10159
rect 11155 10103 11191 10159
rect 11063 9941 11191 10103
rect 11063 9885 11099 9941
rect 11155 9885 11191 9941
rect 11063 9847 11191 9885
rect 11285 10542 11414 10708
rect 11733 10708 11771 10731
rect 11823 10731 12219 10760
rect 11823 10708 11862 10731
rect 11285 10490 11323 10542
rect 11375 10490 11414 10542
rect 11285 10324 11414 10490
rect 11285 10272 11323 10324
rect 11375 10272 11414 10324
rect 11285 10107 11414 10272
rect 11285 10055 11323 10107
rect 11375 10055 11414 10107
rect 11285 9736 11414 10055
rect 11511 10595 11639 10632
rect 11511 10539 11547 10595
rect 11603 10539 11639 10595
rect 11511 10377 11639 10539
rect 11511 10321 11547 10377
rect 11603 10321 11639 10377
rect 11511 10159 11639 10321
rect 11511 10103 11547 10159
rect 11603 10103 11639 10159
rect 11511 9941 11639 10103
rect 11511 9885 11547 9941
rect 11603 9885 11639 9941
rect 11511 9847 11639 9885
rect 11733 10542 11862 10708
rect 12181 10708 12219 10731
rect 12271 10731 12667 10760
rect 12271 10708 12310 10731
rect 11733 10490 11771 10542
rect 11823 10490 11862 10542
rect 11733 10324 11862 10490
rect 11733 10272 11771 10324
rect 11823 10272 11862 10324
rect 11733 10107 11862 10272
rect 11733 10055 11771 10107
rect 11823 10055 11862 10107
rect 11733 9736 11862 10055
rect 11959 10595 12087 10632
rect 11959 10539 11995 10595
rect 12051 10539 12087 10595
rect 11959 10377 12087 10539
rect 11959 10321 11995 10377
rect 12051 10321 12087 10377
rect 11959 10159 12087 10321
rect 11959 10103 11995 10159
rect 12051 10103 12087 10159
rect 11959 9941 12087 10103
rect 11959 9885 11995 9941
rect 12051 9885 12087 9941
rect 11959 9847 12087 9885
rect 12181 10542 12310 10708
rect 12629 10708 12667 10731
rect 12719 10731 13115 10760
rect 12719 10708 12758 10731
rect 12181 10490 12219 10542
rect 12271 10490 12310 10542
rect 12181 10324 12310 10490
rect 12181 10272 12219 10324
rect 12271 10272 12310 10324
rect 12181 10107 12310 10272
rect 12181 10055 12219 10107
rect 12271 10055 12310 10107
rect 12181 9736 12310 10055
rect 12407 10595 12535 10632
rect 12407 10539 12443 10595
rect 12499 10539 12535 10595
rect 12407 10377 12535 10539
rect 12407 10321 12443 10377
rect 12499 10321 12535 10377
rect 12407 10159 12535 10321
rect 12407 10103 12443 10159
rect 12499 10103 12535 10159
rect 12407 9941 12535 10103
rect 12407 9885 12443 9941
rect 12499 9885 12535 9941
rect 12407 9847 12535 9885
rect 12629 10542 12758 10708
rect 13077 10708 13115 10731
rect 13167 10708 13206 10760
rect 12629 10490 12667 10542
rect 12719 10490 12758 10542
rect 12629 10324 12758 10490
rect 12629 10272 12667 10324
rect 12719 10272 12758 10324
rect 12629 10107 12758 10272
rect 12629 10055 12667 10107
rect 12719 10055 12758 10107
rect 12629 9736 12758 10055
rect 12855 10595 12983 10632
rect 12855 10539 12891 10595
rect 12947 10539 12983 10595
rect 12855 10377 12983 10539
rect 12855 10321 12891 10377
rect 12947 10321 12983 10377
rect 12855 10159 12983 10321
rect 12855 10103 12891 10159
rect 12947 10103 12983 10159
rect 12855 9941 12983 10103
rect 12855 9885 12891 9941
rect 12947 9885 12983 9941
rect 12855 9847 12983 9885
rect 13077 10542 13206 10708
rect 13077 10490 13115 10542
rect 13167 10490 13206 10542
rect 13077 10324 13206 10490
rect 13077 10272 13115 10324
rect 13167 10272 13206 10324
rect 13077 10107 13206 10272
rect 13077 10055 13115 10107
rect 13167 10055 13206 10107
rect 13077 9736 13206 10055
rect 13301 10595 13429 10632
rect 13301 10539 13337 10595
rect 13393 10539 13429 10595
rect 13301 10377 13429 10539
rect 13301 10321 13337 10377
rect 13393 10321 13429 10377
rect 13301 10159 13429 10321
rect 13301 10103 13337 10159
rect 13393 10103 13429 10159
rect 13301 9941 13429 10103
rect 13301 9885 13337 9941
rect 13393 9885 13429 9941
rect 13301 9847 13429 9885
rect 13602 10629 13730 10666
rect 13602 10573 13638 10629
rect 13694 10573 13730 10629
rect 13602 10411 13730 10573
rect 13602 10355 13638 10411
rect 13694 10355 13730 10411
rect 13602 10193 13730 10355
rect 13602 10137 13638 10193
rect 13694 10137 13730 10193
rect 13602 9975 13730 10137
rect 13602 9919 13638 9975
rect 13694 9919 13730 9975
rect 13602 9881 13730 9919
rect 8428 9355 13206 9736
rect 6497 9257 6768 9258
rect 6497 9219 6888 9257
rect 6497 9163 6584 9219
rect 6640 9163 6796 9219
rect 6852 9163 6888 9219
rect 6497 9001 6888 9163
rect 6497 8945 6584 9001
rect 6640 8945 6796 9001
rect 6852 8945 6888 9001
rect 6497 8906 6888 8945
rect 8428 8808 8719 9355
rect 4611 8760 8719 8808
rect 4611 8704 4647 8760
rect 4703 8704 4859 8760
rect 4915 8704 8719 8760
rect 4611 8659 8719 8704
rect 9633 8990 10212 9030
rect 9633 8938 9672 8990
rect 9724 8938 10122 8990
rect 10174 8938 10212 8990
rect 9633 8772 10212 8938
rect 9633 8720 9672 8772
rect 9724 8720 10122 8772
rect 10174 8720 10212 8772
rect 9633 8679 10212 8720
rect 419 8260 4132 8298
rect 419 8204 455 8260
rect 511 8204 666 8260
rect 722 8204 876 8260
rect 932 8204 1087 8260
rect 1143 8204 1298 8260
rect 1354 8204 1509 8260
rect 1565 8204 1720 8260
rect 1776 8204 1930 8260
rect 1986 8204 2141 8260
rect 2197 8204 2353 8260
rect 2409 8204 2564 8260
rect 2620 8204 2774 8260
rect 2830 8204 2985 8260
rect 3041 8204 3196 8260
rect 3252 8204 3407 8260
rect 3463 8204 3618 8260
rect 3674 8204 3828 8260
rect 3884 8204 4039 8260
rect 4095 8204 4132 8260
rect 419 8042 4132 8204
rect 419 7986 455 8042
rect 511 7986 666 8042
rect 722 7986 876 8042
rect 932 7986 1087 8042
rect 1143 7986 1298 8042
rect 1354 7986 1509 8042
rect 1565 7986 1720 8042
rect 1776 7986 1930 8042
rect 1986 7986 2141 8042
rect 2197 7986 2353 8042
rect 2409 7986 2564 8042
rect 2620 7986 2774 8042
rect 2830 7986 2985 8042
rect 3041 7986 3196 8042
rect 3252 7986 3407 8042
rect 3463 7986 3618 8042
rect 3674 7986 3828 8042
rect 3884 7986 4039 8042
rect 4095 7986 4132 8042
rect 419 7824 4132 7986
rect 419 7768 455 7824
rect 511 7768 666 7824
rect 722 7768 876 7824
rect 932 7768 1087 7824
rect 1143 7768 1298 7824
rect 1354 7768 1509 7824
rect 1565 7768 1720 7824
rect 1776 7768 1930 7824
rect 1986 7768 2141 7824
rect 2197 7768 2353 7824
rect 2409 7768 2564 7824
rect 2620 7768 2774 7824
rect 2830 7768 2985 7824
rect 3041 7768 3196 7824
rect 3252 7768 3407 7824
rect 3463 7768 3618 7824
rect 3674 7768 3828 7824
rect 3884 7768 4039 7824
rect 4095 7768 4132 7824
rect 419 7730 4132 7768
rect -319 7396 21 7435
rect -319 7340 -283 7396
rect -227 7340 -71 7396
rect -15 7340 21 7396
rect -319 7301 21 7340
rect -279 -2007 -146 7301
rect 704 6863 4418 6902
rect 704 6807 741 6863
rect 797 6807 952 6863
rect 1008 6807 1162 6863
rect 1218 6807 1373 6863
rect 1429 6807 1584 6863
rect 1640 6807 1795 6863
rect 1851 6807 2006 6863
rect 2062 6807 2216 6863
rect 2272 6807 2427 6863
rect 2483 6807 2639 6863
rect 2695 6807 2850 6863
rect 2906 6807 3060 6863
rect 3116 6807 3271 6863
rect 3327 6807 3482 6863
rect 3538 6807 3693 6863
rect 3749 6807 3904 6863
rect 3960 6807 4114 6863
rect 4170 6807 4325 6863
rect 4381 6807 4418 6863
rect 704 6645 4418 6807
rect 704 6589 741 6645
rect 797 6589 952 6645
rect 1008 6589 1162 6645
rect 1218 6589 1373 6645
rect 1429 6589 1584 6645
rect 1640 6589 1795 6645
rect 1851 6589 2006 6645
rect 2062 6589 2216 6645
rect 2272 6589 2427 6645
rect 2483 6589 2639 6645
rect 2695 6589 2850 6645
rect 2906 6589 3060 6645
rect 3116 6589 3271 6645
rect 3327 6589 3482 6645
rect 3538 6589 3693 6645
rect 3749 6589 3904 6645
rect 3960 6589 4114 6645
rect 4170 6589 4325 6645
rect 4381 6589 4418 6645
rect 704 6551 4418 6589
rect 4714 6061 4848 8659
rect 5474 8565 5713 8566
rect 7897 8565 8027 8566
rect 5374 8527 5713 8565
rect 5374 8471 5409 8527
rect 5465 8471 5621 8527
rect 5677 8471 5713 8527
rect 5374 8432 5713 8471
rect 7688 8527 8027 8565
rect 7688 8471 7723 8527
rect 7779 8471 7935 8527
rect 7991 8471 8027 8527
rect 7688 8432 8027 8471
rect 5474 7954 5603 8432
rect 7081 8155 7206 8194
rect 7081 8099 7116 8155
rect 7172 8099 7206 8155
rect 5373 7913 5713 7954
rect 5373 7861 5411 7913
rect 5463 7861 5623 7913
rect 5675 7861 5713 7913
rect 5373 7820 5713 7861
rect 7081 7937 7206 8099
rect 7081 7881 7116 7937
rect 7172 7881 7206 7937
rect 7081 7843 7206 7881
rect 7793 8083 7922 8432
rect 7793 8031 7831 8083
rect 7883 8031 7922 8083
rect 7793 7865 7922 8031
rect 7793 7813 7831 7865
rect 7883 7813 7922 7865
rect 7793 7773 7922 7813
rect 8939 8397 9279 8436
rect 8939 8341 8975 8397
rect 9031 8341 9187 8397
rect 9243 8341 9279 8397
rect 8939 8180 9279 8341
rect 8939 8124 8975 8180
rect 9031 8124 9187 8180
rect 9243 8124 9279 8180
rect 8939 7962 9279 8124
rect 8939 7906 8975 7962
rect 9031 7906 9187 7962
rect 9243 7906 9279 7962
rect 8939 7745 9279 7906
rect 8939 7689 8975 7745
rect 9031 7689 9187 7745
rect 9243 7689 9279 7745
rect 5391 7528 7926 7666
rect 4938 7067 5066 7104
rect 4938 7011 4974 7067
rect 5030 7011 5066 7067
rect 4938 6849 5066 7011
rect 4938 6793 4974 6849
rect 5030 6793 5066 6849
rect 4938 6631 5066 6793
rect 4938 6575 4974 6631
rect 5030 6575 5066 6631
rect 4938 6537 5066 6575
rect 5391 6730 5524 7528
rect 5641 7396 5981 7435
rect 5641 7340 5677 7396
rect 5733 7340 5889 7396
rect 5945 7340 5981 7396
rect 5641 7301 5981 7340
rect 6154 7391 6494 7432
rect 6154 7339 6192 7391
rect 6244 7339 6404 7391
rect 6456 7339 6494 7391
rect 5391 6678 5431 6730
rect 5483 6678 5524 6730
rect 5391 6512 5524 6678
rect 5391 6460 5431 6512
rect 5483 6460 5524 6512
rect 5391 6451 5524 6460
rect 5395 6420 5519 6451
rect 4714 6020 5142 6061
rect 4714 5968 4840 6020
rect 4892 5968 5052 6020
rect 5104 5968 5142 6020
rect 4714 5928 5142 5968
rect 4714 5927 4848 5928
rect 704 5879 4418 5918
rect 704 5823 741 5879
rect 797 5823 952 5879
rect 1008 5823 1162 5879
rect 1218 5823 1373 5879
rect 1429 5823 1584 5879
rect 1640 5823 1795 5879
rect 1851 5823 2006 5879
rect 2062 5823 2216 5879
rect 2272 5823 2427 5879
rect 2483 5823 2639 5879
rect 2695 5823 2850 5879
rect 2906 5823 3060 5879
rect 3116 5823 3271 5879
rect 3327 5823 3482 5879
rect 3538 5823 3693 5879
rect 3749 5823 3904 5879
rect 3960 5823 4114 5879
rect 4170 5823 4325 5879
rect 4381 5823 4418 5879
rect 704 5661 4418 5823
rect 5738 5807 5886 7301
rect 6154 7298 6494 7339
rect 7793 7428 7926 7528
rect 7793 7376 7831 7428
rect 7883 7376 7926 7428
rect 6273 7149 6407 7298
rect 6858 7222 6982 7262
rect 6858 7170 6894 7222
rect 6946 7170 6982 7222
rect 6858 7149 6982 7170
rect 6273 7011 6982 7149
rect 7793 7210 7926 7376
rect 7793 7158 7831 7210
rect 7883 7158 7926 7210
rect 7793 7117 7926 7158
rect 8939 7527 9279 7689
rect 8939 7471 8975 7527
rect 9031 7471 9187 7527
rect 9243 7471 9279 7527
rect 8939 7309 9279 7471
rect 8939 7253 8975 7309
rect 9031 7253 9187 7309
rect 9243 7253 9279 7309
rect 6858 7004 6982 7011
rect 6858 6952 6894 7004
rect 6946 6952 6982 7004
rect 6858 6912 6982 6952
rect 7080 7077 7208 7114
rect 7080 7021 7116 7077
rect 7172 7021 7208 7077
rect 6348 6859 6476 6896
rect 6348 6803 6384 6859
rect 6440 6803 6476 6859
rect 6348 6641 6476 6803
rect 6348 6585 6384 6641
rect 6440 6585 6476 6641
rect 6348 6423 6476 6585
rect 6348 6367 6384 6423
rect 6440 6367 6476 6423
rect 6348 6329 6476 6367
rect 7080 6859 7208 7021
rect 7080 6803 7116 6859
rect 7172 6803 7208 6859
rect 7080 6641 7208 6803
rect 7080 6585 7116 6641
rect 7172 6585 7208 6641
rect 7080 6423 7208 6585
rect 7080 6367 7116 6423
rect 7172 6367 7208 6423
rect 7080 6329 7208 6367
rect 8939 7091 9279 7253
rect 8939 7035 8975 7091
rect 9031 7035 9187 7091
rect 9243 7035 9279 7091
rect 8939 6874 9279 7035
rect 8939 6818 8975 6874
rect 9031 6818 9187 6874
rect 9243 6818 9279 6874
rect 8939 6656 9279 6818
rect 8939 6600 8975 6656
rect 9031 6600 9187 6656
rect 9243 6600 9279 6656
rect 8939 6439 9279 6600
rect 8939 6383 8975 6439
rect 9031 6383 9187 6439
rect 9243 6383 9279 6439
rect 8939 6344 9279 6383
rect 9410 8397 9538 8435
rect 9410 8341 9446 8397
rect 9502 8341 9538 8397
rect 9410 8180 9538 8341
rect 9410 8124 9446 8180
rect 9502 8124 9538 8180
rect 9410 7962 9538 8124
rect 9410 7906 9446 7962
rect 9502 7906 9538 7962
rect 9410 7745 9538 7906
rect 9410 7689 9446 7745
rect 9502 7689 9538 7745
rect 9410 7527 9538 7689
rect 9410 7471 9446 7527
rect 9502 7471 9538 7527
rect 9410 7309 9538 7471
rect 9410 7253 9446 7309
rect 9502 7253 9538 7309
rect 9410 7091 9538 7253
rect 9410 7035 9446 7091
rect 9502 7035 9538 7091
rect 9410 6874 9538 7035
rect 9410 6818 9446 6874
rect 9502 6818 9538 6874
rect 9410 6656 9538 6818
rect 9410 6600 9446 6656
rect 9502 6600 9538 6656
rect 9410 6439 9538 6600
rect 9410 6383 9446 6439
rect 9502 6383 9538 6439
rect 9410 6344 9538 6383
rect 9858 8397 9986 8435
rect 9858 8341 9894 8397
rect 9950 8341 9986 8397
rect 9858 8180 9986 8341
rect 9858 8124 9894 8180
rect 9950 8124 9986 8180
rect 9858 7962 9986 8124
rect 9858 7906 9894 7962
rect 9950 7906 9986 7962
rect 9858 7745 9986 7906
rect 9858 7689 9894 7745
rect 9950 7689 9986 7745
rect 9858 7527 9986 7689
rect 9858 7471 9894 7527
rect 9950 7471 9986 7527
rect 9858 7309 9986 7471
rect 9858 7253 9894 7309
rect 9950 7253 9986 7309
rect 9858 7091 9986 7253
rect 9858 7035 9894 7091
rect 9950 7035 9986 7091
rect 9858 6874 9986 7035
rect 9858 6818 9894 6874
rect 9950 6818 9986 6874
rect 9858 6656 9986 6818
rect 9858 6600 9894 6656
rect 9950 6600 9986 6656
rect 9858 6439 9986 6600
rect 9858 6383 9894 6439
rect 9950 6383 9986 6439
rect 9858 6344 9986 6383
rect 6855 6118 6985 6158
rect 6855 6066 6894 6118
rect 6946 6066 6985 6118
rect 6855 6063 6985 6066
rect 5738 5755 5789 5807
rect 5841 5755 5886 5807
rect 704 5605 741 5661
rect 797 5605 952 5661
rect 1008 5605 1162 5661
rect 1218 5605 1373 5661
rect 1429 5605 1584 5661
rect 1640 5605 1795 5661
rect 1851 5605 2006 5661
rect 2062 5605 2216 5661
rect 2272 5605 2427 5661
rect 2483 5605 2639 5661
rect 2695 5605 2850 5661
rect 2906 5605 3060 5661
rect 3116 5605 3271 5661
rect 3327 5605 3482 5661
rect 3538 5605 3693 5661
rect 3749 5605 3904 5661
rect 3960 5605 4114 5661
rect 4170 5605 4325 5661
rect 4381 5605 4418 5661
rect 704 5567 4418 5605
rect 5164 5628 5289 5667
rect 5164 5572 5198 5628
rect 5254 5572 5289 5628
rect 5164 5410 5289 5572
rect 5164 5354 5198 5410
rect 5254 5354 5289 5410
rect 5164 5316 5289 5354
rect 5738 5589 5886 5755
rect 6349 5972 6474 6011
rect 6349 5916 6384 5972
rect 6440 5916 6474 5972
rect 6349 5754 6474 5916
rect 6855 5930 10100 6063
rect 6855 5900 6985 5930
rect 6855 5848 6894 5900
rect 6946 5848 6985 5900
rect 6855 5807 6985 5848
rect 6349 5698 6384 5754
rect 6440 5698 6474 5754
rect 6349 5660 6474 5698
rect 5738 5537 5789 5589
rect 5841 5537 5886 5589
rect 5738 5496 5886 5537
rect 5738 5363 9874 5496
rect 217 4939 5405 4977
rect 217 4883 253 4939
rect 309 4883 464 4939
rect 520 4883 675 4939
rect 731 4883 885 4939
rect 941 4883 1096 4939
rect 1152 4883 1307 4939
rect 1363 4883 1518 4939
rect 1574 4883 1729 4939
rect 1785 4883 1939 4939
rect 1995 4883 2150 4939
rect 2206 4883 2361 4939
rect 2417 4883 2572 4939
rect 2628 4883 2783 4939
rect 2839 4883 2994 4939
rect 3050 4883 3205 4939
rect 3261 4883 3416 4939
rect 3472 4883 3627 4939
rect 3683 4883 3837 4939
rect 3893 4883 4048 4939
rect 4104 4883 4259 4939
rect 4315 4883 4470 4939
rect 4526 4883 4681 4939
rect 4737 4883 4891 4939
rect 4947 4883 5102 4939
rect 5158 4883 5313 4939
rect 5369 4883 5405 4939
rect 217 4721 5405 4883
rect 217 4665 253 4721
rect 309 4665 464 4721
rect 520 4665 675 4721
rect 731 4665 885 4721
rect 941 4665 1096 4721
rect 1152 4665 1307 4721
rect 1363 4665 1518 4721
rect 1574 4665 1729 4721
rect 1785 4665 1939 4721
rect 1995 4665 2150 4721
rect 2206 4665 2361 4721
rect 2417 4665 2572 4721
rect 2628 4665 2783 4721
rect 2839 4665 2994 4721
rect 3050 4665 3205 4721
rect 3261 4665 3416 4721
rect 3472 4665 3627 4721
rect 3683 4665 3837 4721
rect 3893 4665 4048 4721
rect 4104 4665 4259 4721
rect 4315 4665 4470 4721
rect 4526 4665 4681 4721
rect 4737 4665 4891 4721
rect 4947 4665 5102 4721
rect 5158 4665 5313 4721
rect 5369 4665 5405 4721
rect 217 4503 5405 4665
rect 217 4447 253 4503
rect 309 4447 464 4503
rect 520 4447 675 4503
rect 731 4447 885 4503
rect 941 4447 1096 4503
rect 1152 4447 1307 4503
rect 1363 4447 1518 4503
rect 1574 4447 1729 4503
rect 1785 4447 1939 4503
rect 1995 4447 2150 4503
rect 2206 4447 2361 4503
rect 2417 4447 2572 4503
rect 2628 4447 2783 4503
rect 2839 4447 2994 4503
rect 3050 4447 3205 4503
rect 3261 4447 3416 4503
rect 3472 4447 3627 4503
rect 3683 4447 3837 4503
rect 3893 4447 4048 4503
rect 4104 4447 4259 4503
rect 4315 4447 4470 4503
rect 4526 4447 4681 4503
rect 4737 4447 4891 4503
rect 4947 4447 5102 4503
rect 5158 4447 5313 4503
rect 5369 4447 5405 4503
rect 217 4285 5405 4447
rect 217 4229 253 4285
rect 309 4229 464 4285
rect 520 4229 675 4285
rect 731 4229 885 4285
rect 941 4229 1096 4285
rect 1152 4229 1307 4285
rect 1363 4229 1518 4285
rect 1574 4229 1729 4285
rect 1785 4229 1939 4285
rect 1995 4229 2150 4285
rect 2206 4229 2361 4285
rect 2417 4229 2572 4285
rect 2628 4229 2783 4285
rect 2839 4229 2994 4285
rect 3050 4229 3205 4285
rect 3261 4229 3416 4285
rect 3472 4229 3627 4285
rect 3683 4229 3837 4285
rect 3893 4229 4048 4285
rect 4104 4229 4259 4285
rect 4315 4229 4470 4285
rect 4526 4229 4681 4285
rect 4737 4229 4891 4285
rect 4947 4229 5102 4285
rect 5158 4229 5313 4285
rect 5369 4229 5405 4285
rect 217 4191 5405 4229
rect 5738 3599 5886 5363
rect 8585 5208 8925 5249
rect 8585 5156 8623 5208
rect 8675 5156 8835 5208
rect 8887 5156 8925 5208
rect 8585 5115 8925 5156
rect 9745 5201 9874 5363
rect 9971 5201 10100 5930
rect 9745 5161 9875 5201
rect 5325 3558 5886 3599
rect 5325 3506 5362 3558
rect 5414 3506 5574 3558
rect 5626 3506 5886 3558
rect 5325 3466 5886 3506
rect 8024 3065 8100 3075
rect 2514 2732 7606 2742
rect 2514 2676 2524 2732
rect 2580 2676 2656 2732
rect 2712 2676 2788 2732
rect 2844 2676 2920 2732
rect 2976 2676 3052 2732
rect 3108 2676 3184 2732
rect 3240 2676 3316 2732
rect 3372 2676 3448 2732
rect 3504 2676 3580 2732
rect 3636 2676 3712 2732
rect 3768 2676 3844 2732
rect 3900 2676 3976 2732
rect 4032 2676 4108 2732
rect 4164 2676 4240 2732
rect 4296 2676 4372 2732
rect 4428 2676 4504 2732
rect 4560 2676 4636 2732
rect 4692 2676 4768 2732
rect 4824 2676 4900 2732
rect 4956 2676 5032 2732
rect 5088 2676 5164 2732
rect 5220 2676 5296 2732
rect 5352 2676 5428 2732
rect 5484 2676 5560 2732
rect 5616 2676 5692 2732
rect 5748 2676 5824 2732
rect 5880 2676 5956 2732
rect 6012 2676 6088 2732
rect 6144 2676 6220 2732
rect 6276 2676 6352 2732
rect 6408 2676 6484 2732
rect 6540 2676 6616 2732
rect 6672 2676 6748 2732
rect 6804 2676 6880 2732
rect 6936 2676 7012 2732
rect 7068 2676 7144 2732
rect 7200 2676 7276 2732
rect 7332 2676 7408 2732
rect 7464 2676 7540 2732
rect 7596 2676 7606 2732
rect 8024 2697 8034 3065
rect 8090 2697 8100 3065
rect 8024 2687 8100 2697
rect 8472 3065 8548 3075
rect 8472 2697 8482 3065
rect 8538 2697 8548 3065
rect 8472 2687 8548 2697
rect 2514 2600 7606 2676
rect 2514 2544 2524 2600
rect 2580 2544 2656 2600
rect 2712 2544 2788 2600
rect 2844 2544 2920 2600
rect 2976 2544 3052 2600
rect 3108 2544 3184 2600
rect 3240 2544 3316 2600
rect 3372 2544 3448 2600
rect 3504 2544 3580 2600
rect 3636 2544 3712 2600
rect 3768 2544 3844 2600
rect 3900 2544 3976 2600
rect 4032 2544 4108 2600
rect 4164 2544 4240 2600
rect 4296 2544 4372 2600
rect 4428 2544 4504 2600
rect 4560 2544 4636 2600
rect 4692 2544 4768 2600
rect 4824 2544 4900 2600
rect 4956 2544 5032 2600
rect 5088 2544 5164 2600
rect 5220 2544 5296 2600
rect 5352 2544 5428 2600
rect 5484 2544 5560 2600
rect 5616 2544 5692 2600
rect 5748 2544 5824 2600
rect 5880 2544 5956 2600
rect 6012 2544 6088 2600
rect 6144 2544 6220 2600
rect 6276 2544 6352 2600
rect 6408 2544 6484 2600
rect 6540 2544 6616 2600
rect 6672 2544 6748 2600
rect 6804 2544 6880 2600
rect 6936 2544 7012 2600
rect 7068 2544 7144 2600
rect 7200 2544 7276 2600
rect 7332 2544 7408 2600
rect 7464 2544 7540 2600
rect 7596 2544 7606 2600
rect 2514 2468 7606 2544
rect 2514 2412 2524 2468
rect 2580 2412 2656 2468
rect 2712 2412 2788 2468
rect 2844 2412 2920 2468
rect 2976 2412 3052 2468
rect 3108 2412 3184 2468
rect 3240 2412 3316 2468
rect 3372 2412 3448 2468
rect 3504 2412 3580 2468
rect 3636 2412 3712 2468
rect 3768 2412 3844 2468
rect 3900 2412 3976 2468
rect 4032 2412 4108 2468
rect 4164 2412 4240 2468
rect 4296 2412 4372 2468
rect 4428 2412 4504 2468
rect 4560 2412 4636 2468
rect 4692 2412 4768 2468
rect 4824 2412 4900 2468
rect 4956 2412 5032 2468
rect 5088 2412 5164 2468
rect 5220 2412 5296 2468
rect 5352 2412 5428 2468
rect 5484 2412 5560 2468
rect 5616 2412 5692 2468
rect 5748 2412 5824 2468
rect 5880 2412 5956 2468
rect 6012 2412 6088 2468
rect 6144 2412 6220 2468
rect 6276 2412 6352 2468
rect 6408 2412 6484 2468
rect 6540 2412 6616 2468
rect 6672 2412 6748 2468
rect 6804 2412 6880 2468
rect 6936 2412 7012 2468
rect 7068 2412 7144 2468
rect 7200 2412 7276 2468
rect 7332 2412 7408 2468
rect 7464 2412 7540 2468
rect 7596 2412 7606 2468
rect 2514 2336 7606 2412
rect 2514 2280 2524 2336
rect 2580 2280 2656 2336
rect 2712 2280 2788 2336
rect 2844 2280 2920 2336
rect 2976 2280 3052 2336
rect 3108 2280 3184 2336
rect 3240 2280 3316 2336
rect 3372 2280 3448 2336
rect 3504 2280 3580 2336
rect 3636 2280 3712 2336
rect 3768 2280 3844 2336
rect 3900 2280 3976 2336
rect 4032 2280 4108 2336
rect 4164 2280 4240 2336
rect 4296 2280 4372 2336
rect 4428 2280 4504 2336
rect 4560 2280 4636 2336
rect 4692 2280 4768 2336
rect 4824 2280 4900 2336
rect 4956 2280 5032 2336
rect 5088 2280 5164 2336
rect 5220 2280 5296 2336
rect 5352 2280 5428 2336
rect 5484 2280 5560 2336
rect 5616 2280 5692 2336
rect 5748 2280 5824 2336
rect 5880 2280 5956 2336
rect 6012 2280 6088 2336
rect 6144 2280 6220 2336
rect 6276 2280 6352 2336
rect 6408 2280 6484 2336
rect 6540 2280 6616 2336
rect 6672 2280 6748 2336
rect 6804 2280 6880 2336
rect 6936 2280 7012 2336
rect 7068 2280 7144 2336
rect 7200 2280 7276 2336
rect 7332 2280 7408 2336
rect 7464 2280 7540 2336
rect 7596 2280 7606 2336
rect 2514 2270 7606 2280
rect 8689 -253 8822 5115
rect 9745 5109 9784 5161
rect 9836 5109 9875 5161
rect 9745 4943 9875 5109
rect 9745 4891 9784 4943
rect 9836 4891 9875 4943
rect 9745 4850 9875 4891
rect 9971 5161 10101 5201
rect 9971 5109 10010 5161
rect 10062 5109 10101 5161
rect 9971 4943 10101 5109
rect 9971 4891 10010 4943
rect 10062 4891 10101 4943
rect 9971 4850 10101 4891
rect 8944 4703 9283 4741
rect 8944 4647 8979 4703
rect 9035 4647 9191 4703
rect 9247 4647 9283 4703
rect 8944 4485 9283 4647
rect 8944 4429 8979 4485
rect 9035 4429 9191 4485
rect 9247 4429 9283 4485
rect 8944 4267 9283 4429
rect 8944 4211 8979 4267
rect 9035 4211 9191 4267
rect 9247 4211 9283 4267
rect 8944 4049 9283 4211
rect 8944 3993 8979 4049
rect 9035 3993 9191 4049
rect 9247 3993 9283 4049
rect 8944 3955 9283 3993
rect 9416 4736 9545 4775
rect 9416 4680 9452 4736
rect 9508 4680 9545 4736
rect 9416 4519 9545 4680
rect 9416 4463 9452 4519
rect 9508 4463 9545 4519
rect 9416 4301 9545 4463
rect 9416 4245 9452 4301
rect 9508 4245 9545 4301
rect 9416 4083 9545 4245
rect 9416 4027 9452 4083
rect 9508 4027 9545 4083
rect 9416 3866 9545 4027
rect 9416 3810 9452 3866
rect 9508 3810 9545 3866
rect 9416 3648 9545 3810
rect 9416 3592 9452 3648
rect 9508 3592 9545 3648
rect 9416 3431 9545 3592
rect 9416 3375 9452 3431
rect 9508 3375 9545 3431
rect 9416 3213 9545 3375
rect 9416 3157 9452 3213
rect 9508 3157 9545 3213
rect 9416 2995 9545 3157
rect 9416 2939 9452 2995
rect 9508 2939 9545 2995
rect 9416 2778 9545 2939
rect 9416 2722 9452 2778
rect 9508 2722 9545 2778
rect 9416 2560 9545 2722
rect 9416 2504 9452 2560
rect 9508 2504 9545 2560
rect 9416 2342 9545 2504
rect 9416 2286 9452 2342
rect 9508 2286 9545 2342
rect 9416 2125 9545 2286
rect 9416 2069 9452 2125
rect 9508 2069 9545 2125
rect 9416 1907 9545 2069
rect 9416 1851 9452 1907
rect 9508 1851 9545 1907
rect 9416 1689 9545 1851
rect 9416 1633 9452 1689
rect 9508 1633 9545 1689
rect 9416 1472 9545 1633
rect 9416 1416 9452 1472
rect 9508 1416 9545 1472
rect 9416 1254 9545 1416
rect 9416 1198 9452 1254
rect 9508 1198 9545 1254
rect 9416 1037 9545 1198
rect 9416 981 9452 1037
rect 9508 981 9545 1037
rect 9416 819 9545 981
rect 9416 763 9452 819
rect 9508 763 9545 819
rect 9416 601 9545 763
rect 9416 545 9452 601
rect 9508 545 9545 601
rect 9416 384 9545 545
rect 9416 328 9452 384
rect 9508 328 9545 384
rect 9416 289 9545 328
rect 10321 -436 10450 9355
rect 11812 9330 13206 9355
rect 11812 9274 11847 9330
rect 11903 9274 12058 9330
rect 12114 9274 12269 9330
rect 12325 9274 12480 9330
rect 12536 9274 12691 9330
rect 12747 9274 12902 9330
rect 12958 9274 13113 9330
rect 13169 9274 13206 9330
rect 10607 9219 10732 9258
rect 10607 9163 10642 9219
rect 10698 9163 10732 9219
rect 10607 9137 10732 9163
rect 11058 9219 11183 9258
rect 11058 9163 11093 9219
rect 11149 9163 11183 9219
rect 11058 9137 11183 9163
rect 11506 9219 11631 9258
rect 11506 9163 11541 9219
rect 11597 9163 11631 9219
rect 11506 9137 11631 9163
rect 10607 9097 10738 9137
rect 10607 9045 10647 9097
rect 10699 9045 10738 9097
rect 10607 9001 10738 9045
rect 10607 8945 10642 9001
rect 10698 8945 10738 9001
rect 10607 8907 10738 8945
rect 10608 8879 10738 8907
rect 10608 8827 10647 8879
rect 10699 8827 10738 8879
rect 10608 8661 10738 8827
rect 10608 8609 10647 8661
rect 10699 8609 10738 8661
rect 10608 8444 10738 8609
rect 10608 8392 10647 8444
rect 10699 8392 10738 8444
rect 11056 9097 11186 9137
rect 11056 9045 11095 9097
rect 11147 9045 11186 9097
rect 11056 9001 11186 9045
rect 11056 8945 11093 9001
rect 11149 8945 11186 9001
rect 11056 8879 11186 8945
rect 11056 8827 11095 8879
rect 11147 8827 11186 8879
rect 11056 8661 11186 8827
rect 11056 8609 11095 8661
rect 11147 8609 11186 8661
rect 11056 8444 11186 8609
rect 10608 8226 10738 8392
rect 10608 8174 10647 8226
rect 10699 8174 10738 8226
rect 10608 8008 10738 8174
rect 10608 7956 10647 8008
rect 10699 7956 10738 8008
rect 10608 7791 10738 7956
rect 10608 7739 10647 7791
rect 10699 7739 10738 7791
rect 10608 7573 10738 7739
rect 10608 7521 10647 7573
rect 10699 7521 10738 7573
rect 10608 7356 10738 7521
rect 10608 7304 10647 7356
rect 10699 7304 10738 7356
rect 10608 7138 10738 7304
rect 10608 7086 10647 7138
rect 10699 7086 10738 7138
rect 10608 6920 10738 7086
rect 10608 6868 10647 6920
rect 10699 6868 10738 6920
rect 10608 6702 10738 6868
rect 10608 6650 10647 6702
rect 10699 6650 10738 6702
rect 10608 6485 10738 6650
rect 10608 6433 10647 6485
rect 10699 6433 10738 6485
rect 10608 6267 10738 6433
rect 10833 8388 10961 8426
rect 10833 8332 10869 8388
rect 10925 8332 10961 8388
rect 10833 8171 10961 8332
rect 10833 8115 10869 8171
rect 10925 8115 10961 8171
rect 10833 7953 10961 8115
rect 10833 7897 10869 7953
rect 10925 7897 10961 7953
rect 10833 7736 10961 7897
rect 10833 7680 10869 7736
rect 10925 7680 10961 7736
rect 10833 7518 10961 7680
rect 10833 7462 10869 7518
rect 10925 7462 10961 7518
rect 10833 7300 10961 7462
rect 10833 7244 10869 7300
rect 10925 7244 10961 7300
rect 10833 7082 10961 7244
rect 10833 7026 10869 7082
rect 10925 7026 10961 7082
rect 10833 6865 10961 7026
rect 10833 6809 10869 6865
rect 10925 6809 10961 6865
rect 10833 6647 10961 6809
rect 10833 6591 10869 6647
rect 10925 6591 10961 6647
rect 10833 6430 10961 6591
rect 10833 6374 10869 6430
rect 10925 6374 10961 6430
rect 10833 6335 10961 6374
rect 11056 8392 11095 8444
rect 11147 8392 11186 8444
rect 11504 9097 11634 9137
rect 11504 9045 11543 9097
rect 11595 9045 11634 9097
rect 11504 9001 11634 9045
rect 11504 8945 11541 9001
rect 11597 8945 11634 9001
rect 11504 8879 11634 8945
rect 11504 8827 11543 8879
rect 11595 8827 11634 8879
rect 11504 8661 11634 8827
rect 11504 8609 11543 8661
rect 11595 8609 11634 8661
rect 11504 8444 11634 8609
rect 11812 9112 13206 9274
rect 11812 9056 11847 9112
rect 11903 9056 12058 9112
rect 12114 9056 12269 9112
rect 12325 9056 12480 9112
rect 12536 9056 12691 9112
rect 12747 9056 12902 9112
rect 12958 9056 13113 9112
rect 13169 9056 13206 9112
rect 11812 8894 13206 9056
rect 11812 8838 11847 8894
rect 11903 8838 12058 8894
rect 12114 8838 12269 8894
rect 12325 8838 12480 8894
rect 12536 8838 12691 8894
rect 12747 8838 12902 8894
rect 12958 8838 13113 8894
rect 13169 8838 13206 8894
rect 11812 8676 13206 8838
rect 11812 8620 11847 8676
rect 11903 8620 12058 8676
rect 12114 8620 12269 8676
rect 12325 8620 12480 8676
rect 12536 8620 12691 8676
rect 12747 8620 12902 8676
rect 12958 8620 13113 8676
rect 13169 8620 13206 8676
rect 11812 8555 13206 8620
rect 11056 8226 11186 8392
rect 11056 8174 11095 8226
rect 11147 8174 11186 8226
rect 11056 8008 11186 8174
rect 11056 7956 11095 8008
rect 11147 7956 11186 8008
rect 11056 7791 11186 7956
rect 11056 7739 11095 7791
rect 11147 7739 11186 7791
rect 11056 7573 11186 7739
rect 11056 7521 11095 7573
rect 11147 7521 11186 7573
rect 11056 7356 11186 7521
rect 11056 7304 11095 7356
rect 11147 7304 11186 7356
rect 11056 7138 11186 7304
rect 11056 7086 11095 7138
rect 11147 7086 11186 7138
rect 11056 6920 11186 7086
rect 11056 6868 11095 6920
rect 11147 6868 11186 6920
rect 11056 6702 11186 6868
rect 11056 6650 11095 6702
rect 11147 6650 11186 6702
rect 11056 6485 11186 6650
rect 11056 6433 11095 6485
rect 11147 6433 11186 6485
rect 10608 6215 10647 6267
rect 10699 6215 10738 6267
rect 10608 6050 10738 6215
rect 10608 5998 10647 6050
rect 10699 5998 10738 6050
rect 10608 5832 10738 5998
rect 10608 5780 10647 5832
rect 10699 5780 10738 5832
rect 10608 5614 10738 5780
rect 10608 5562 10647 5614
rect 10699 5562 10738 5614
rect 10608 5397 10738 5562
rect 10608 5345 10647 5397
rect 10699 5345 10738 5397
rect 10608 5331 10738 5345
rect 11056 6267 11186 6433
rect 11281 8388 11409 8426
rect 11281 8332 11317 8388
rect 11373 8332 11409 8388
rect 11281 8171 11409 8332
rect 11281 8115 11317 8171
rect 11373 8115 11409 8171
rect 11281 7953 11409 8115
rect 11281 7897 11317 7953
rect 11373 7897 11409 7953
rect 11281 7736 11409 7897
rect 11281 7680 11317 7736
rect 11373 7680 11409 7736
rect 11281 7518 11409 7680
rect 11281 7462 11317 7518
rect 11373 7462 11409 7518
rect 11281 7300 11409 7462
rect 11281 7244 11317 7300
rect 11373 7244 11409 7300
rect 11281 7082 11409 7244
rect 11281 7026 11317 7082
rect 11373 7026 11409 7082
rect 11281 6865 11409 7026
rect 11281 6809 11317 6865
rect 11373 6809 11409 6865
rect 11281 6647 11409 6809
rect 11281 6591 11317 6647
rect 11373 6591 11409 6647
rect 11281 6430 11409 6591
rect 11281 6374 11317 6430
rect 11373 6374 11409 6430
rect 11281 6335 11409 6374
rect 11504 8392 11543 8444
rect 11595 8392 11634 8444
rect 11504 8226 11634 8392
rect 11504 8174 11543 8226
rect 11595 8174 11634 8226
rect 11504 8008 11634 8174
rect 11504 7956 11543 8008
rect 11595 7956 11634 8008
rect 11504 7791 11634 7956
rect 11504 7739 11543 7791
rect 11595 7739 11634 7791
rect 11504 7573 11634 7739
rect 11504 7521 11543 7573
rect 11595 7521 11634 7573
rect 11504 7356 11634 7521
rect 11504 7304 11543 7356
rect 11595 7304 11634 7356
rect 11504 7138 11634 7304
rect 11504 7086 11543 7138
rect 11595 7086 11634 7138
rect 11504 6920 11634 7086
rect 11504 6868 11543 6920
rect 11595 6868 11634 6920
rect 11504 6702 11634 6868
rect 11504 6650 11543 6702
rect 11595 6650 11634 6702
rect 11504 6485 11634 6650
rect 11504 6433 11543 6485
rect 11595 6433 11634 6485
rect 11056 6215 11095 6267
rect 11147 6215 11186 6267
rect 11056 6050 11186 6215
rect 11056 5998 11095 6050
rect 11147 5998 11186 6050
rect 11056 5832 11186 5998
rect 11056 5780 11095 5832
rect 11147 5780 11186 5832
rect 11056 5614 11186 5780
rect 11056 5562 11095 5614
rect 11147 5562 11186 5614
rect 11056 5397 11186 5562
rect 11056 5345 11095 5397
rect 11147 5345 11186 5397
rect 11056 5331 11186 5345
rect 11504 6267 11634 6433
rect 12115 8402 12243 8440
rect 12115 8346 12151 8402
rect 12207 8346 12243 8402
rect 12115 8185 12243 8346
rect 12115 8129 12151 8185
rect 12207 8129 12243 8185
rect 12115 7967 12243 8129
rect 12115 7911 12151 7967
rect 12207 7911 12243 7967
rect 12115 7750 12243 7911
rect 12115 7694 12151 7750
rect 12207 7694 12243 7750
rect 12115 7532 12243 7694
rect 12115 7476 12151 7532
rect 12207 7476 12243 7532
rect 12115 7314 12243 7476
rect 12115 7258 12151 7314
rect 12207 7258 12243 7314
rect 12115 7096 12243 7258
rect 12115 7040 12151 7096
rect 12207 7040 12243 7096
rect 12115 6879 12243 7040
rect 12115 6823 12151 6879
rect 12207 6823 12243 6879
rect 12115 6661 12243 6823
rect 12115 6605 12151 6661
rect 12207 6605 12243 6661
rect 12115 6444 12243 6605
rect 12115 6388 12151 6444
rect 12207 6388 12243 6444
rect 12115 6349 12243 6388
rect 12563 8402 12691 8440
rect 12563 8346 12599 8402
rect 12655 8346 12691 8402
rect 12563 8185 12691 8346
rect 12563 8129 12599 8185
rect 12655 8129 12691 8185
rect 12563 7967 12691 8129
rect 12563 7911 12599 7967
rect 12655 7911 12691 7967
rect 12563 7750 12691 7911
rect 12563 7694 12599 7750
rect 12655 7694 12691 7750
rect 12563 7532 12691 7694
rect 12563 7476 12599 7532
rect 12655 7476 12691 7532
rect 12563 7314 12691 7476
rect 12563 7258 12599 7314
rect 12655 7258 12691 7314
rect 12563 7096 12691 7258
rect 12563 7040 12599 7096
rect 12655 7040 12691 7096
rect 12563 6879 12691 7040
rect 12563 6823 12599 6879
rect 12655 6823 12691 6879
rect 12563 6661 12691 6823
rect 12563 6605 12599 6661
rect 12655 6605 12691 6661
rect 12563 6444 12691 6605
rect 12563 6388 12599 6444
rect 12655 6388 12691 6444
rect 12563 6349 12691 6388
rect 11504 6215 11543 6267
rect 11595 6215 11634 6267
rect 11504 6050 11634 6215
rect 11504 5998 11543 6050
rect 11595 5998 11634 6050
rect 11504 5832 11634 5998
rect 11504 5780 11543 5832
rect 11595 5780 11634 5832
rect 11504 5614 11634 5780
rect 11504 5562 11543 5614
rect 11595 5562 11634 5614
rect 11504 5397 11634 5562
rect 11504 5345 11543 5397
rect 11595 5345 11634 5397
rect 11504 5331 11634 5345
rect 10608 5179 11634 5331
rect 10608 5127 10647 5179
rect 10699 5127 11095 5179
rect 11147 5127 11543 5179
rect 11595 5127 11634 5179
rect 10608 4961 11634 5127
rect 10608 4909 10647 4961
rect 10699 4909 11095 4961
rect 11147 4909 11543 4961
rect 11595 4909 11634 4961
rect 10608 4869 11634 4909
rect 11893 5413 12918 5453
rect 11893 5361 11931 5413
rect 11983 5361 12379 5413
rect 12431 5361 12827 5413
rect 12879 5361 12918 5413
rect 11893 5195 12918 5361
rect 11893 5143 11931 5195
rect 11983 5143 12379 5195
rect 12431 5143 12827 5195
rect 12879 5143 12918 5195
rect 11893 4977 12918 5143
rect 11893 4925 11931 4977
rect 11983 4925 12379 4977
rect 12431 4925 12827 4977
rect 12879 4925 12918 4977
rect 11063 4331 11179 4869
rect 11893 4759 12918 4925
rect 11893 4707 11931 4759
rect 11983 4707 12379 4759
rect 12431 4707 12827 4759
rect 12879 4707 12918 4759
rect 11893 4667 12918 4707
rect 11063 4290 11897 4331
rect 11063 4238 11595 4290
rect 11647 4238 11807 4290
rect 11859 4238 11897 4290
rect 11063 4198 11897 4238
rect 11063 4104 11179 4198
rect 12348 4104 12463 4667
rect 12595 4514 12935 4553
rect 12595 4458 12631 4514
rect 12687 4458 12843 4514
rect 12899 4458 12935 4514
rect 12595 4419 12935 4458
rect 11057 4064 11186 4104
rect 10609 3993 10738 4032
rect 10609 3937 10645 3993
rect 10701 3937 10738 3993
rect 10609 3775 10738 3937
rect 10609 3719 10645 3775
rect 10701 3719 10738 3775
rect 10609 3558 10738 3719
rect 10609 3502 10645 3558
rect 10701 3502 10738 3558
rect 10609 3340 10738 3502
rect 10609 3284 10645 3340
rect 10701 3284 10738 3340
rect 10609 3122 10738 3284
rect 10609 3066 10645 3122
rect 10701 3066 10738 3122
rect 10609 2905 10738 3066
rect 10609 2849 10645 2905
rect 10701 2849 10738 2905
rect 10609 2687 10738 2849
rect 10609 2631 10645 2687
rect 10701 2631 10738 2687
rect 10609 2470 10738 2631
rect 10609 2414 10645 2470
rect 10701 2414 10738 2470
rect 10609 2252 10738 2414
rect 10609 2196 10645 2252
rect 10701 2196 10738 2252
rect 11057 4012 11095 4064
rect 11147 4012 11186 4064
rect 12341 4064 12470 4104
rect 11057 3846 11186 4012
rect 11057 3794 11095 3846
rect 11147 3794 11186 3846
rect 11057 3628 11186 3794
rect 11057 3576 11095 3628
rect 11147 3576 11186 3628
rect 11057 3411 11186 3576
rect 11057 3359 11095 3411
rect 11147 3359 11186 3411
rect 11057 3193 11186 3359
rect 11057 3141 11095 3193
rect 11147 3141 11186 3193
rect 11057 2975 11186 3141
rect 11057 2923 11095 2975
rect 11147 2923 11186 2975
rect 11057 2758 11186 2923
rect 11057 2706 11095 2758
rect 11147 2706 11186 2758
rect 11057 2540 11186 2706
rect 11057 2488 11095 2540
rect 11147 2488 11186 2540
rect 11057 2322 11186 2488
rect 11057 2270 11095 2322
rect 11147 2270 11186 2322
rect 11057 2230 11186 2270
rect 11505 3993 11634 4032
rect 11505 3937 11541 3993
rect 11597 3937 11634 3993
rect 11505 3775 11634 3937
rect 11505 3719 11541 3775
rect 11597 3719 11634 3775
rect 11505 3558 11634 3719
rect 11505 3502 11541 3558
rect 11597 3502 11634 3558
rect 11505 3340 11634 3502
rect 11505 3284 11541 3340
rect 11597 3284 11634 3340
rect 11505 3122 11634 3284
rect 11505 3066 11541 3122
rect 11597 3066 11634 3122
rect 11505 2905 11634 3066
rect 11505 2849 11541 2905
rect 11597 2849 11634 2905
rect 11505 2687 11634 2849
rect 11505 2631 11541 2687
rect 11597 2631 11634 2687
rect 11505 2470 11634 2631
rect 11505 2414 11541 2470
rect 11597 2414 11634 2470
rect 11505 2252 11634 2414
rect 10609 2034 10738 2196
rect 10609 1978 10645 2034
rect 10701 1978 10738 2034
rect 10609 1816 10738 1978
rect 10609 1760 10645 1816
rect 10701 1760 10738 1816
rect 10609 1599 10738 1760
rect 10609 1543 10645 1599
rect 10701 1543 10738 1599
rect 10609 1381 10738 1543
rect 10609 1325 10645 1381
rect 10701 1325 10738 1381
rect 10609 1164 10738 1325
rect 10609 1108 10645 1164
rect 10701 1108 10738 1164
rect 10609 946 10738 1108
rect 10609 890 10645 946
rect 10701 890 10738 946
rect 10609 728 10738 890
rect 10609 672 10645 728
rect 10701 672 10738 728
rect 10609 511 10738 672
rect 10609 455 10645 511
rect 10701 455 10738 511
rect 10609 293 10738 455
rect 10609 237 10645 293
rect 10701 237 10738 293
rect 10609 199 10738 237
rect 11505 2196 11541 2252
rect 11597 2196 11634 2252
rect 11505 2034 11634 2196
rect 11505 1978 11541 2034
rect 11597 1978 11634 2034
rect 11505 1816 11634 1978
rect 11505 1760 11541 1816
rect 11597 1760 11634 1816
rect 11505 1599 11634 1760
rect 11505 1543 11541 1599
rect 11597 1543 11634 1599
rect 11505 1381 11634 1543
rect 11505 1325 11541 1381
rect 11597 1325 11634 1381
rect 11505 1164 11634 1325
rect 11505 1108 11541 1164
rect 11597 1108 11634 1164
rect 11505 946 11634 1108
rect 11505 890 11541 946
rect 11597 890 11634 946
rect 11505 728 11634 890
rect 11505 672 11541 728
rect 11597 672 11634 728
rect 11505 511 11634 672
rect 11505 455 11541 511
rect 11597 455 11634 511
rect 11505 293 11634 455
rect 11505 237 11541 293
rect 11597 237 11634 293
rect 11505 199 11634 237
rect 11893 3993 12022 4032
rect 11893 3937 11929 3993
rect 11985 3937 12022 3993
rect 11893 3775 12022 3937
rect 11893 3719 11929 3775
rect 11985 3719 12022 3775
rect 11893 3558 12022 3719
rect 11893 3502 11929 3558
rect 11985 3502 12022 3558
rect 11893 3340 12022 3502
rect 11893 3284 11929 3340
rect 11985 3284 12022 3340
rect 11893 3122 12022 3284
rect 11893 3066 11929 3122
rect 11985 3066 12022 3122
rect 11893 2905 12022 3066
rect 11893 2849 11929 2905
rect 11985 2849 12022 2905
rect 11893 2687 12022 2849
rect 11893 2631 11929 2687
rect 11985 2631 12022 2687
rect 11893 2470 12022 2631
rect 11893 2414 11929 2470
rect 11985 2414 12022 2470
rect 11893 2252 12022 2414
rect 11893 2196 11929 2252
rect 11985 2196 12022 2252
rect 12341 4012 12379 4064
rect 12431 4012 12470 4064
rect 12341 3846 12470 4012
rect 12341 3794 12379 3846
rect 12431 3794 12470 3846
rect 12341 3628 12470 3794
rect 12341 3576 12379 3628
rect 12431 3576 12470 3628
rect 12341 3411 12470 3576
rect 12341 3359 12379 3411
rect 12431 3359 12470 3411
rect 12341 3193 12470 3359
rect 12341 3141 12379 3193
rect 12431 3141 12470 3193
rect 12341 2975 12470 3141
rect 12341 2923 12379 2975
rect 12431 2923 12470 2975
rect 12341 2758 12470 2923
rect 12341 2706 12379 2758
rect 12431 2706 12470 2758
rect 12341 2540 12470 2706
rect 12341 2488 12379 2540
rect 12431 2488 12470 2540
rect 12341 2322 12470 2488
rect 12341 2270 12379 2322
rect 12431 2270 12470 2322
rect 12341 2230 12470 2270
rect 12789 3993 12918 4032
rect 12789 3937 12825 3993
rect 12881 3937 12918 3993
rect 12789 3775 12918 3937
rect 12789 3719 12825 3775
rect 12881 3719 12918 3775
rect 12789 3558 12918 3719
rect 12789 3502 12825 3558
rect 12881 3502 12918 3558
rect 12789 3340 12918 3502
rect 12789 3284 12825 3340
rect 12881 3284 12918 3340
rect 12789 3122 12918 3284
rect 12789 3066 12825 3122
rect 12881 3066 12918 3122
rect 12789 2905 12918 3066
rect 12789 2849 12825 2905
rect 12881 2849 12918 2905
rect 12789 2687 12918 2849
rect 12789 2631 12825 2687
rect 12881 2631 12918 2687
rect 12789 2470 12918 2631
rect 12789 2414 12825 2470
rect 12881 2414 12918 2470
rect 12789 2252 12918 2414
rect 11893 2034 12022 2196
rect 11893 1978 11929 2034
rect 11985 1978 12022 2034
rect 11893 1816 12022 1978
rect 11893 1760 11929 1816
rect 11985 1760 12022 1816
rect 11893 1599 12022 1760
rect 11893 1543 11929 1599
rect 11985 1543 12022 1599
rect 11893 1381 12022 1543
rect 11893 1325 11929 1381
rect 11985 1325 12022 1381
rect 11893 1164 12022 1325
rect 11893 1108 11929 1164
rect 11985 1108 12022 1164
rect 11893 946 12022 1108
rect 11893 890 11929 946
rect 11985 890 12022 946
rect 11893 728 12022 890
rect 11893 672 11929 728
rect 11985 672 12022 728
rect 11893 511 12022 672
rect 11893 455 11929 511
rect 11985 455 12022 511
rect 11893 293 12022 455
rect 11893 237 11929 293
rect 11985 237 12022 293
rect 11893 199 12022 237
rect 12789 2196 12825 2252
rect 12881 2196 12918 2252
rect 12789 2034 12918 2196
rect 12789 1978 12825 2034
rect 12881 1978 12918 2034
rect 12789 1816 12918 1978
rect 12789 1760 12825 1816
rect 12881 1760 12918 1816
rect 12789 1599 12918 1760
rect 12789 1543 12825 1599
rect 12881 1543 12918 1599
rect 12789 1381 12918 1543
rect 12789 1325 12825 1381
rect 12881 1325 12918 1381
rect 12789 1164 12918 1325
rect 12789 1108 12825 1164
rect 12881 1108 12918 1164
rect 12789 946 12918 1108
rect 12789 890 12825 946
rect 12881 890 12918 946
rect 12789 728 12918 890
rect 12789 672 12825 728
rect 12881 672 12918 728
rect 12789 511 12918 672
rect 12789 455 12825 511
rect 12881 455 12918 511
rect 12789 293 12918 455
rect 12789 237 12825 293
rect 12881 237 12918 293
rect 12789 199 12918 237
rect 13044 -436 13173 8555
rect 13362 8402 13490 8440
rect 13362 8346 13398 8402
rect 13454 8346 13490 8402
rect 13362 8185 13490 8346
rect 13362 8129 13398 8185
rect 13454 8129 13490 8185
rect 13362 7967 13490 8129
rect 13362 7911 13398 7967
rect 13454 7911 13490 7967
rect 13362 7750 13490 7911
rect 13362 7694 13398 7750
rect 13454 7694 13490 7750
rect 13362 7532 13490 7694
rect 13362 7476 13398 7532
rect 13454 7476 13490 7532
rect 13362 7314 13490 7476
rect 13362 7258 13398 7314
rect 13454 7258 13490 7314
rect 13362 7096 13490 7258
rect 13362 7040 13398 7096
rect 13454 7040 13490 7096
rect 13362 6879 13490 7040
rect 13362 6823 13398 6879
rect 13454 6823 13490 6879
rect 13362 6661 13490 6823
rect 13362 6605 13398 6661
rect 13454 6605 13490 6661
rect 13362 6444 13490 6605
rect 13362 6388 13398 6444
rect 13454 6388 13490 6444
rect 13362 6349 13490 6388
rect 13477 3993 13606 4032
rect 13477 3937 13513 3993
rect 13569 3937 13606 3993
rect 13477 3775 13606 3937
rect 13477 3719 13513 3775
rect 13569 3719 13606 3775
rect 13477 3558 13606 3719
rect 13477 3502 13513 3558
rect 13569 3502 13606 3558
rect 13477 3340 13606 3502
rect 13477 3284 13513 3340
rect 13569 3284 13606 3340
rect 13477 3122 13606 3284
rect 13477 3066 13513 3122
rect 13569 3066 13606 3122
rect 13477 2905 13606 3066
rect 13477 2849 13513 2905
rect 13569 2849 13606 2905
rect 13477 2687 13606 2849
rect 13477 2631 13513 2687
rect 13569 2631 13606 2687
rect 13477 2470 13606 2631
rect 13477 2414 13513 2470
rect 13569 2414 13606 2470
rect 13477 2252 13606 2414
rect 13477 2196 13513 2252
rect 13569 2196 13606 2252
rect 13477 2034 13606 2196
rect 13477 1978 13513 2034
rect 13569 1978 13606 2034
rect 13477 1816 13606 1978
rect 13477 1760 13513 1816
rect 13569 1760 13606 1816
rect 13477 1599 13606 1760
rect 13477 1543 13513 1599
rect 13569 1543 13606 1599
rect 13477 1381 13606 1543
rect 13477 1325 13513 1381
rect 13569 1325 13606 1381
rect 13477 1164 13606 1325
rect 13477 1108 13513 1164
rect 13569 1108 13606 1164
rect 13477 946 13606 1108
rect 13477 890 13513 946
rect 13569 890 13606 946
rect 13477 728 13606 890
rect 13477 672 13513 728
rect 13569 672 13606 728
rect 13477 511 13606 672
rect 13477 455 13513 511
rect 13569 455 13606 511
rect 13477 293 13606 455
rect 13477 237 13513 293
rect 13569 237 13606 293
rect 13477 199 13606 237
rect 10215 -477 10555 -436
rect 10215 -529 10253 -477
rect 10305 -529 10465 -477
rect 10517 -529 10555 -477
rect 10215 -695 10555 -529
rect 10215 -747 10253 -695
rect 10305 -747 10465 -695
rect 10517 -747 10555 -695
rect 10215 -787 10555 -747
rect 12938 -477 13278 -436
rect 12938 -529 12976 -477
rect 13028 -529 13188 -477
rect 13240 -529 13278 -477
rect 12938 -695 13278 -529
rect 12938 -747 12976 -695
rect 13028 -747 13188 -695
rect 13240 -747 13278 -695
rect 12938 -787 13278 -747
rect -383 -2046 -43 -2007
rect -383 -2102 -347 -2046
rect -291 -2102 -135 -2046
rect -79 -2102 -43 -2046
rect -383 -2140 -43 -2102
rect -280 -2141 -146 -2140
<< via2 >>
rect 6327 16238 6383 16240
rect 6327 16186 6329 16238
rect 6329 16186 6381 16238
rect 6381 16186 6383 16238
rect 6327 16184 6383 16186
rect 6775 16238 6831 16240
rect 6775 16186 6777 16238
rect 6777 16186 6829 16238
rect 6829 16186 6831 16238
rect 6775 16184 6831 16186
rect 7223 16238 7279 16240
rect 7223 16186 7225 16238
rect 7225 16186 7277 16238
rect 7277 16186 7279 16238
rect 7223 16184 7279 16186
rect 7671 16238 7727 16240
rect 7671 16186 7673 16238
rect 7673 16186 7725 16238
rect 7725 16186 7727 16238
rect 7671 16184 7727 16186
rect 8119 16238 8175 16240
rect 8119 16186 8121 16238
rect 8121 16186 8173 16238
rect 8173 16186 8175 16238
rect 8119 16184 8175 16186
rect 8567 16238 8623 16240
rect 8567 16186 8569 16238
rect 8569 16186 8621 16238
rect 8621 16186 8623 16238
rect 8567 16184 8623 16186
rect 8857 16238 8913 16240
rect 8857 16186 8859 16238
rect 8859 16186 8911 16238
rect 8911 16186 8913 16238
rect 8857 16184 8913 16186
rect 9305 16238 9361 16240
rect 9305 16186 9307 16238
rect 9307 16186 9359 16238
rect 9359 16186 9361 16238
rect 9305 16184 9361 16186
rect 9753 16238 9809 16240
rect 9753 16186 9755 16238
rect 9755 16186 9807 16238
rect 9807 16186 9809 16238
rect 9753 16184 9809 16186
rect 10201 16238 10257 16240
rect 10201 16186 10203 16238
rect 10203 16186 10255 16238
rect 10255 16186 10257 16238
rect 10201 16184 10257 16186
rect 10649 16238 10705 16240
rect 10649 16186 10651 16238
rect 10651 16186 10703 16238
rect 10703 16186 10705 16238
rect 10649 16184 10705 16186
rect 11097 16238 11153 16240
rect 11097 16186 11099 16238
rect 11099 16186 11151 16238
rect 11151 16186 11153 16238
rect 11097 16184 11153 16186
rect 11545 16238 11601 16240
rect 11545 16186 11547 16238
rect 11547 16186 11599 16238
rect 11599 16186 11601 16238
rect 11545 16184 11601 16186
rect 11993 16238 12049 16240
rect 11993 16186 11995 16238
rect 11995 16186 12047 16238
rect 12047 16186 12049 16238
rect 11993 16184 12049 16186
rect 12441 16238 12497 16240
rect 12441 16186 12443 16238
rect 12443 16186 12495 16238
rect 12495 16186 12497 16238
rect 12441 16184 12497 16186
rect 12889 16238 12945 16240
rect 12889 16186 12891 16238
rect 12891 16186 12943 16238
rect 12943 16186 12945 16238
rect 12889 16184 12945 16186
rect 13337 16238 13393 16240
rect 13337 16186 13339 16238
rect 13339 16186 13391 16238
rect 13391 16186 13393 16238
rect 13337 16184 13393 16186
rect 6327 16020 6383 16022
rect 6327 15968 6329 16020
rect 6329 15968 6381 16020
rect 6381 15968 6383 16020
rect 6327 15966 6383 15968
rect 6775 16020 6831 16022
rect 6775 15968 6777 16020
rect 6777 15968 6829 16020
rect 6829 15968 6831 16020
rect 6775 15966 6831 15968
rect 7223 16020 7279 16022
rect 7223 15968 7225 16020
rect 7225 15968 7277 16020
rect 7277 15968 7279 16020
rect 7223 15966 7279 15968
rect 7671 16020 7727 16022
rect 7671 15968 7673 16020
rect 7673 15968 7725 16020
rect 7725 15968 7727 16020
rect 7671 15966 7727 15968
rect 8119 16020 8175 16022
rect 8119 15968 8121 16020
rect 8121 15968 8173 16020
rect 8173 15968 8175 16020
rect 8119 15966 8175 15968
rect 8567 16020 8623 16022
rect 8567 15968 8569 16020
rect 8569 15968 8621 16020
rect 8621 15968 8623 16020
rect 8567 15966 8623 15968
rect 8857 16020 8913 16022
rect 8857 15968 8859 16020
rect 8859 15968 8911 16020
rect 8911 15968 8913 16020
rect 8857 15966 8913 15968
rect 9305 16020 9361 16022
rect 9305 15968 9307 16020
rect 9307 15968 9359 16020
rect 9359 15968 9361 16020
rect 9305 15966 9361 15968
rect 9753 16020 9809 16022
rect 9753 15968 9755 16020
rect 9755 15968 9807 16020
rect 9807 15968 9809 16020
rect 9753 15966 9809 15968
rect 10201 16020 10257 16022
rect 10201 15968 10203 16020
rect 10203 15968 10255 16020
rect 10255 15968 10257 16020
rect 10201 15966 10257 15968
rect 10649 16020 10705 16022
rect 10649 15968 10651 16020
rect 10651 15968 10703 16020
rect 10703 15968 10705 16020
rect 10649 15966 10705 15968
rect 11097 16020 11153 16022
rect 11097 15968 11099 16020
rect 11099 15968 11151 16020
rect 11151 15968 11153 16020
rect 11097 15966 11153 15968
rect 11545 16020 11601 16022
rect 11545 15968 11547 16020
rect 11547 15968 11599 16020
rect 11599 15968 11601 16020
rect 11545 15966 11601 15968
rect 11993 16020 12049 16022
rect 11993 15968 11995 16020
rect 11995 15968 12047 16020
rect 12047 15968 12049 16020
rect 11993 15966 12049 15968
rect 12441 16020 12497 16022
rect 12441 15968 12443 16020
rect 12443 15968 12495 16020
rect 12495 15968 12497 16020
rect 12441 15966 12497 15968
rect 12889 16020 12945 16022
rect 12889 15968 12891 16020
rect 12891 15968 12943 16020
rect 12943 15968 12945 16020
rect 12889 15966 12945 15968
rect 13337 16020 13393 16022
rect 13337 15968 13339 16020
rect 13339 15968 13391 16020
rect 13391 15968 13393 16020
rect 13337 15966 13393 15968
rect 6327 15803 6383 15805
rect 6327 15751 6329 15803
rect 6329 15751 6381 15803
rect 6381 15751 6383 15803
rect 6327 15749 6383 15751
rect 6775 15803 6831 15805
rect 6775 15751 6777 15803
rect 6777 15751 6829 15803
rect 6829 15751 6831 15803
rect 6775 15749 6831 15751
rect 7223 15803 7279 15805
rect 7223 15751 7225 15803
rect 7225 15751 7277 15803
rect 7277 15751 7279 15803
rect 7223 15749 7279 15751
rect 7671 15803 7727 15805
rect 7671 15751 7673 15803
rect 7673 15751 7725 15803
rect 7725 15751 7727 15803
rect 7671 15749 7727 15751
rect 8119 15803 8175 15805
rect 8119 15751 8121 15803
rect 8121 15751 8173 15803
rect 8173 15751 8175 15803
rect 8119 15749 8175 15751
rect 8567 15803 8623 15805
rect 8567 15751 8569 15803
rect 8569 15751 8621 15803
rect 8621 15751 8623 15803
rect 8567 15749 8623 15751
rect 8857 15803 8913 15805
rect 8857 15751 8859 15803
rect 8859 15751 8911 15803
rect 8911 15751 8913 15803
rect 8857 15749 8913 15751
rect 9305 15803 9361 15805
rect 9305 15751 9307 15803
rect 9307 15751 9359 15803
rect 9359 15751 9361 15803
rect 9305 15749 9361 15751
rect 9753 15803 9809 15805
rect 9753 15751 9755 15803
rect 9755 15751 9807 15803
rect 9807 15751 9809 15803
rect 9753 15749 9809 15751
rect 10201 15803 10257 15805
rect 10201 15751 10203 15803
rect 10203 15751 10255 15803
rect 10255 15751 10257 15803
rect 10201 15749 10257 15751
rect 10649 15803 10705 15805
rect 10649 15751 10651 15803
rect 10651 15751 10703 15803
rect 10703 15751 10705 15803
rect 10649 15749 10705 15751
rect 11097 15803 11153 15805
rect 11097 15751 11099 15803
rect 11099 15751 11151 15803
rect 11151 15751 11153 15803
rect 11097 15749 11153 15751
rect 11545 15803 11601 15805
rect 11545 15751 11547 15803
rect 11547 15751 11599 15803
rect 11599 15751 11601 15803
rect 11545 15749 11601 15751
rect 11993 15803 12049 15805
rect 11993 15751 11995 15803
rect 11995 15751 12047 15803
rect 12047 15751 12049 15803
rect 11993 15749 12049 15751
rect 12441 15803 12497 15805
rect 12441 15751 12443 15803
rect 12443 15751 12495 15803
rect 12495 15751 12497 15803
rect 12441 15749 12497 15751
rect 12889 15803 12945 15805
rect 12889 15751 12891 15803
rect 12891 15751 12943 15803
rect 12943 15751 12945 15803
rect 12889 15749 12945 15751
rect 13337 15803 13393 15805
rect 13337 15751 13339 15803
rect 13339 15751 13391 15803
rect 13391 15751 13393 15803
rect 13337 15749 13393 15751
rect 6327 15585 6383 15587
rect 6327 15533 6329 15585
rect 6329 15533 6381 15585
rect 6381 15533 6383 15585
rect 6327 15531 6383 15533
rect 6775 15585 6831 15587
rect 6775 15533 6777 15585
rect 6777 15533 6829 15585
rect 6829 15533 6831 15585
rect 6775 15531 6831 15533
rect 7223 15585 7279 15587
rect 7223 15533 7225 15585
rect 7225 15533 7277 15585
rect 7277 15533 7279 15585
rect 7223 15531 7279 15533
rect 7671 15585 7727 15587
rect 7671 15533 7673 15585
rect 7673 15533 7725 15585
rect 7725 15533 7727 15585
rect 7671 15531 7727 15533
rect 8119 15585 8175 15587
rect 8119 15533 8121 15585
rect 8121 15533 8173 15585
rect 8173 15533 8175 15585
rect 8119 15531 8175 15533
rect 8567 15585 8623 15587
rect 8567 15533 8569 15585
rect 8569 15533 8621 15585
rect 8621 15533 8623 15585
rect 8567 15531 8623 15533
rect 8857 15585 8913 15587
rect 8857 15533 8859 15585
rect 8859 15533 8911 15585
rect 8911 15533 8913 15585
rect 8857 15531 8913 15533
rect 9305 15585 9361 15587
rect 9305 15533 9307 15585
rect 9307 15533 9359 15585
rect 9359 15533 9361 15585
rect 9305 15531 9361 15533
rect 9753 15585 9809 15587
rect 9753 15533 9755 15585
rect 9755 15533 9807 15585
rect 9807 15533 9809 15585
rect 9753 15531 9809 15533
rect 10201 15585 10257 15587
rect 10201 15533 10203 15585
rect 10203 15533 10255 15585
rect 10255 15533 10257 15585
rect 10201 15531 10257 15533
rect 10649 15585 10705 15587
rect 10649 15533 10651 15585
rect 10651 15533 10703 15585
rect 10703 15533 10705 15585
rect 10649 15531 10705 15533
rect 11097 15585 11153 15587
rect 11097 15533 11099 15585
rect 11099 15533 11151 15585
rect 11151 15533 11153 15585
rect 11097 15531 11153 15533
rect 11545 15585 11601 15587
rect 11545 15533 11547 15585
rect 11547 15533 11599 15585
rect 11599 15533 11601 15585
rect 11545 15531 11601 15533
rect 11993 15585 12049 15587
rect 11993 15533 11995 15585
rect 11995 15533 12047 15585
rect 12047 15533 12049 15585
rect 11993 15531 12049 15533
rect 12441 15585 12497 15587
rect 12441 15533 12443 15585
rect 12443 15533 12495 15585
rect 12495 15533 12497 15585
rect 12441 15531 12497 15533
rect 12889 15585 12945 15587
rect 12889 15533 12891 15585
rect 12891 15533 12943 15585
rect 12943 15533 12945 15585
rect 12889 15531 12945 15533
rect 13337 15585 13393 15587
rect 13337 15533 13339 15585
rect 13339 15533 13391 15585
rect 13391 15533 13393 15585
rect 13337 15531 13393 15533
rect 6327 15367 6383 15369
rect 6327 15315 6329 15367
rect 6329 15315 6381 15367
rect 6381 15315 6383 15367
rect 6327 15313 6383 15315
rect 6775 15367 6831 15369
rect 6775 15315 6777 15367
rect 6777 15315 6829 15367
rect 6829 15315 6831 15367
rect 6775 15313 6831 15315
rect 7223 15367 7279 15369
rect 7223 15315 7225 15367
rect 7225 15315 7277 15367
rect 7277 15315 7279 15367
rect 7223 15313 7279 15315
rect 7671 15367 7727 15369
rect 7671 15315 7673 15367
rect 7673 15315 7725 15367
rect 7725 15315 7727 15367
rect 7671 15313 7727 15315
rect 8119 15367 8175 15369
rect 8119 15315 8121 15367
rect 8121 15315 8173 15367
rect 8173 15315 8175 15367
rect 8119 15313 8175 15315
rect 8567 15367 8623 15369
rect 8567 15315 8569 15367
rect 8569 15315 8621 15367
rect 8621 15315 8623 15367
rect 8567 15313 8623 15315
rect 8857 15367 8913 15369
rect 8857 15315 8859 15367
rect 8859 15315 8911 15367
rect 8911 15315 8913 15367
rect 8857 15313 8913 15315
rect 9305 15367 9361 15369
rect 9305 15315 9307 15367
rect 9307 15315 9359 15367
rect 9359 15315 9361 15367
rect 9305 15313 9361 15315
rect 9753 15367 9809 15369
rect 9753 15315 9755 15367
rect 9755 15315 9807 15367
rect 9807 15315 9809 15367
rect 9753 15313 9809 15315
rect 10201 15367 10257 15369
rect 10201 15315 10203 15367
rect 10203 15315 10255 15367
rect 10255 15315 10257 15367
rect 10201 15313 10257 15315
rect 10649 15367 10705 15369
rect 10649 15315 10651 15367
rect 10651 15315 10703 15367
rect 10703 15315 10705 15367
rect 10649 15313 10705 15315
rect 11097 15367 11153 15369
rect 11097 15315 11099 15367
rect 11099 15315 11151 15367
rect 11151 15315 11153 15367
rect 11097 15313 11153 15315
rect 11545 15367 11601 15369
rect 11545 15315 11547 15367
rect 11547 15315 11599 15367
rect 11599 15315 11601 15367
rect 11545 15313 11601 15315
rect 11993 15367 12049 15369
rect 11993 15315 11995 15367
rect 11995 15315 12047 15367
rect 12047 15315 12049 15367
rect 11993 15313 12049 15315
rect 12441 15367 12497 15369
rect 12441 15315 12443 15367
rect 12443 15315 12495 15367
rect 12495 15315 12497 15367
rect 12441 15313 12497 15315
rect 12889 15367 12945 15369
rect 12889 15315 12891 15367
rect 12891 15315 12943 15367
rect 12943 15315 12945 15367
rect 12889 15313 12945 15315
rect 13337 15367 13393 15369
rect 13337 15315 13339 15367
rect 13339 15315 13391 15367
rect 13391 15315 13393 15367
rect 13337 15313 13393 15315
rect 6327 15149 6383 15151
rect 6327 15097 6329 15149
rect 6329 15097 6381 15149
rect 6381 15097 6383 15149
rect 6327 15095 6383 15097
rect 6775 15149 6831 15151
rect 6775 15097 6777 15149
rect 6777 15097 6829 15149
rect 6829 15097 6831 15149
rect 6775 15095 6831 15097
rect 7223 15149 7279 15151
rect 7223 15097 7225 15149
rect 7225 15097 7277 15149
rect 7277 15097 7279 15149
rect 7223 15095 7279 15097
rect 7671 15149 7727 15151
rect 7671 15097 7673 15149
rect 7673 15097 7725 15149
rect 7725 15097 7727 15149
rect 7671 15095 7727 15097
rect 8119 15149 8175 15151
rect 8119 15097 8121 15149
rect 8121 15097 8173 15149
rect 8173 15097 8175 15149
rect 8119 15095 8175 15097
rect 8567 15149 8623 15151
rect 8567 15097 8569 15149
rect 8569 15097 8621 15149
rect 8621 15097 8623 15149
rect 8567 15095 8623 15097
rect 8857 15149 8913 15151
rect 8857 15097 8859 15149
rect 8859 15097 8911 15149
rect 8911 15097 8913 15149
rect 8857 15095 8913 15097
rect 9305 15149 9361 15151
rect 9305 15097 9307 15149
rect 9307 15097 9359 15149
rect 9359 15097 9361 15149
rect 9305 15095 9361 15097
rect 9753 15149 9809 15151
rect 9753 15097 9755 15149
rect 9755 15097 9807 15149
rect 9807 15097 9809 15149
rect 9753 15095 9809 15097
rect 10201 15149 10257 15151
rect 10201 15097 10203 15149
rect 10203 15097 10255 15149
rect 10255 15097 10257 15149
rect 10201 15095 10257 15097
rect 10649 15149 10705 15151
rect 10649 15097 10651 15149
rect 10651 15097 10703 15149
rect 10703 15097 10705 15149
rect 10649 15095 10705 15097
rect 11097 15149 11153 15151
rect 11097 15097 11099 15149
rect 11099 15097 11151 15149
rect 11151 15097 11153 15149
rect 11097 15095 11153 15097
rect 11545 15149 11601 15151
rect 11545 15097 11547 15149
rect 11547 15097 11599 15149
rect 11599 15097 11601 15149
rect 11545 15095 11601 15097
rect 11993 15149 12049 15151
rect 11993 15097 11995 15149
rect 11995 15097 12047 15149
rect 12047 15097 12049 15149
rect 11993 15095 12049 15097
rect 12441 15149 12497 15151
rect 12441 15097 12443 15149
rect 12443 15097 12495 15149
rect 12495 15097 12497 15149
rect 12441 15095 12497 15097
rect 12889 15149 12945 15151
rect 12889 15097 12891 15149
rect 12891 15097 12943 15149
rect 12943 15097 12945 15149
rect 12889 15095 12945 15097
rect 13337 15149 13393 15151
rect 13337 15097 13339 15149
rect 13339 15097 13391 15149
rect 13391 15097 13393 15149
rect 13337 15095 13393 15097
rect 6327 14932 6383 14934
rect 6327 14880 6329 14932
rect 6329 14880 6381 14932
rect 6381 14880 6383 14932
rect 6327 14878 6383 14880
rect 6775 14932 6831 14934
rect 6775 14880 6777 14932
rect 6777 14880 6829 14932
rect 6829 14880 6831 14932
rect 6775 14878 6831 14880
rect 7223 14932 7279 14934
rect 7223 14880 7225 14932
rect 7225 14880 7277 14932
rect 7277 14880 7279 14932
rect 7223 14878 7279 14880
rect 7671 14932 7727 14934
rect 7671 14880 7673 14932
rect 7673 14880 7725 14932
rect 7725 14880 7727 14932
rect 7671 14878 7727 14880
rect 8119 14932 8175 14934
rect 8119 14880 8121 14932
rect 8121 14880 8173 14932
rect 8173 14880 8175 14932
rect 8119 14878 8175 14880
rect 8567 14932 8623 14934
rect 8567 14880 8569 14932
rect 8569 14880 8621 14932
rect 8621 14880 8623 14932
rect 8567 14878 8623 14880
rect 8857 14932 8913 14934
rect 8857 14880 8859 14932
rect 8859 14880 8911 14932
rect 8911 14880 8913 14932
rect 8857 14878 8913 14880
rect 9305 14932 9361 14934
rect 9305 14880 9307 14932
rect 9307 14880 9359 14932
rect 9359 14880 9361 14932
rect 9305 14878 9361 14880
rect 9753 14932 9809 14934
rect 9753 14880 9755 14932
rect 9755 14880 9807 14932
rect 9807 14880 9809 14932
rect 9753 14878 9809 14880
rect 10201 14932 10257 14934
rect 10201 14880 10203 14932
rect 10203 14880 10255 14932
rect 10255 14880 10257 14932
rect 10201 14878 10257 14880
rect 10649 14932 10705 14934
rect 10649 14880 10651 14932
rect 10651 14880 10703 14932
rect 10703 14880 10705 14932
rect 10649 14878 10705 14880
rect 11097 14932 11153 14934
rect 11097 14880 11099 14932
rect 11099 14880 11151 14932
rect 11151 14880 11153 14932
rect 11097 14878 11153 14880
rect 11545 14932 11601 14934
rect 11545 14880 11547 14932
rect 11547 14880 11599 14932
rect 11599 14880 11601 14932
rect 11545 14878 11601 14880
rect 11993 14932 12049 14934
rect 11993 14880 11995 14932
rect 11995 14880 12047 14932
rect 12047 14880 12049 14932
rect 11993 14878 12049 14880
rect 12441 14932 12497 14934
rect 12441 14880 12443 14932
rect 12443 14880 12495 14932
rect 12495 14880 12497 14932
rect 12441 14878 12497 14880
rect 12889 14932 12945 14934
rect 12889 14880 12891 14932
rect 12891 14880 12943 14932
rect 12943 14880 12945 14932
rect 12889 14878 12945 14880
rect 13337 14932 13393 14934
rect 13337 14880 13339 14932
rect 13339 14880 13391 14932
rect 13391 14880 13393 14932
rect 13337 14878 13393 14880
rect 6327 14714 6383 14716
rect 6327 14662 6329 14714
rect 6329 14662 6381 14714
rect 6381 14662 6383 14714
rect 6327 14660 6383 14662
rect 6775 14714 6831 14716
rect 6775 14662 6777 14714
rect 6777 14662 6829 14714
rect 6829 14662 6831 14714
rect 6775 14660 6831 14662
rect 7223 14714 7279 14716
rect 7223 14662 7225 14714
rect 7225 14662 7277 14714
rect 7277 14662 7279 14714
rect 7223 14660 7279 14662
rect 7671 14714 7727 14716
rect 7671 14662 7673 14714
rect 7673 14662 7725 14714
rect 7725 14662 7727 14714
rect 7671 14660 7727 14662
rect 8119 14714 8175 14716
rect 8119 14662 8121 14714
rect 8121 14662 8173 14714
rect 8173 14662 8175 14714
rect 8119 14660 8175 14662
rect 8567 14714 8623 14716
rect 8567 14662 8569 14714
rect 8569 14662 8621 14714
rect 8621 14662 8623 14714
rect 8567 14660 8623 14662
rect 8857 14714 8913 14716
rect 8857 14662 8859 14714
rect 8859 14662 8911 14714
rect 8911 14662 8913 14714
rect 8857 14660 8913 14662
rect 9305 14714 9361 14716
rect 9305 14662 9307 14714
rect 9307 14662 9359 14714
rect 9359 14662 9361 14714
rect 9305 14660 9361 14662
rect 9753 14714 9809 14716
rect 9753 14662 9755 14714
rect 9755 14662 9807 14714
rect 9807 14662 9809 14714
rect 9753 14660 9809 14662
rect 10201 14714 10257 14716
rect 10201 14662 10203 14714
rect 10203 14662 10255 14714
rect 10255 14662 10257 14714
rect 10201 14660 10257 14662
rect 10649 14714 10705 14716
rect 10649 14662 10651 14714
rect 10651 14662 10703 14714
rect 10703 14662 10705 14714
rect 10649 14660 10705 14662
rect 11097 14714 11153 14716
rect 11097 14662 11099 14714
rect 11099 14662 11151 14714
rect 11151 14662 11153 14714
rect 11097 14660 11153 14662
rect 11545 14714 11601 14716
rect 11545 14662 11547 14714
rect 11547 14662 11599 14714
rect 11599 14662 11601 14714
rect 11545 14660 11601 14662
rect 11993 14714 12049 14716
rect 11993 14662 11995 14714
rect 11995 14662 12047 14714
rect 12047 14662 12049 14714
rect 11993 14660 12049 14662
rect 12441 14714 12497 14716
rect 12441 14662 12443 14714
rect 12443 14662 12495 14714
rect 12495 14662 12497 14714
rect 12441 14660 12497 14662
rect 12889 14714 12945 14716
rect 12889 14662 12891 14714
rect 12891 14662 12943 14714
rect 12943 14662 12945 14714
rect 12889 14660 12945 14662
rect 13337 14714 13393 14716
rect 13337 14662 13339 14714
rect 13339 14662 13391 14714
rect 13391 14662 13393 14714
rect 13337 14660 13393 14662
rect 6312 11293 6368 11295
rect 6312 11241 6314 11293
rect 6314 11241 6366 11293
rect 6366 11241 6368 11293
rect 6312 11239 6368 11241
rect 6312 11075 6368 11077
rect 6312 11023 6314 11075
rect 6314 11023 6366 11075
rect 6366 11023 6368 11075
rect 6312 11021 6368 11023
rect 6312 10858 6368 10860
rect 6312 10806 6314 10858
rect 6314 10806 6366 10858
rect 6366 10806 6368 10858
rect 6312 10804 6368 10806
rect 6312 10640 6368 10642
rect 6312 10588 6314 10640
rect 6314 10588 6366 10640
rect 6366 10588 6368 10640
rect 6312 10586 6368 10588
rect 6312 10422 6368 10424
rect 6312 10370 6314 10422
rect 6314 10370 6366 10422
rect 6366 10370 6368 10422
rect 6312 10368 6368 10370
rect 6312 10205 6368 10207
rect 6312 10153 6314 10205
rect 6314 10153 6366 10205
rect 6366 10153 6368 10205
rect 6312 10151 6368 10153
rect 6312 9987 6368 9989
rect 6312 9935 6314 9987
rect 6314 9935 6366 9987
rect 6366 9935 6368 9987
rect 6312 9933 6368 9935
rect 7068 10262 7124 10264
rect 7068 10210 7070 10262
rect 7070 10210 7122 10262
rect 7122 10210 7124 10262
rect 7068 10208 7124 10210
rect 7068 10044 7124 10046
rect 7068 9992 7070 10044
rect 7070 9992 7122 10044
rect 7122 9992 7124 10044
rect 7068 9990 7124 9992
rect 7068 9826 7124 9828
rect 7068 9774 7070 9826
rect 7070 9774 7122 9826
rect 7122 9774 7124 9826
rect 7068 9772 7124 9774
rect 7068 9608 7124 9610
rect 7068 9556 7070 9608
rect 7070 9556 7122 9608
rect 7122 9556 7124 9608
rect 7068 9554 7124 9556
rect 7515 10262 7571 10264
rect 7515 10210 7517 10262
rect 7517 10210 7569 10262
rect 7569 10210 7571 10262
rect 7515 10208 7571 10210
rect 7515 10044 7571 10046
rect 7515 9992 7517 10044
rect 7517 9992 7569 10044
rect 7569 9992 7571 10044
rect 7515 9990 7571 9992
rect 7515 9826 7571 9828
rect 7515 9774 7517 9826
rect 7517 9774 7569 9826
rect 7569 9774 7571 9826
rect 7515 9772 7571 9774
rect 7515 9608 7571 9610
rect 7515 9556 7517 9608
rect 7517 9556 7569 9608
rect 7569 9556 7571 9608
rect 7515 9554 7571 9556
rect 8015 10474 8071 10476
rect 8015 10422 8017 10474
rect 8017 10422 8069 10474
rect 8069 10422 8071 10474
rect 8015 10420 8071 10422
rect 8227 10474 8283 10476
rect 8227 10422 8229 10474
rect 8229 10422 8281 10474
rect 8281 10422 8283 10474
rect 8227 10420 8283 10422
rect 8015 10257 8071 10259
rect 8015 10205 8017 10257
rect 8017 10205 8069 10257
rect 8069 10205 8071 10257
rect 8015 10203 8071 10205
rect 8227 10257 8283 10259
rect 8227 10205 8229 10257
rect 8229 10205 8281 10257
rect 8281 10205 8283 10257
rect 8227 10203 8283 10205
rect 8015 10039 8071 10041
rect 8015 9987 8017 10039
rect 8017 9987 8069 10039
rect 8069 9987 8071 10039
rect 8015 9985 8071 9987
rect 8227 10039 8283 10041
rect 8227 9987 8229 10039
rect 8229 9987 8281 10039
rect 8281 9987 8283 10039
rect 8227 9985 8283 9987
rect 8015 9821 8071 9823
rect 8015 9769 8017 9821
rect 8017 9769 8069 9821
rect 8069 9769 8071 9821
rect 8015 9767 8071 9769
rect 8227 9821 8283 9823
rect 8227 9769 8229 9821
rect 8229 9769 8281 9821
rect 8281 9769 8283 9821
rect 8227 9767 8283 9769
rect 8015 9604 8071 9606
rect 8015 9552 8017 9604
rect 8017 9552 8069 9604
rect 8069 9552 8071 9604
rect 8015 9550 8071 9552
rect 8227 9604 8283 9606
rect 8227 9552 8229 9604
rect 8229 9552 8281 9604
rect 8281 9552 8283 9604
rect 8227 9550 8283 9552
rect 8859 10593 8915 10595
rect 8859 10541 8861 10593
rect 8861 10541 8913 10593
rect 8913 10541 8915 10593
rect 8859 10539 8915 10541
rect 8859 10375 8915 10377
rect 8859 10323 8861 10375
rect 8861 10323 8913 10375
rect 8913 10323 8915 10375
rect 8859 10321 8915 10323
rect 8859 10157 8915 10159
rect 8859 10105 8861 10157
rect 8861 10105 8913 10157
rect 8913 10105 8915 10157
rect 8859 10103 8915 10105
rect 8859 9939 8915 9941
rect 8859 9887 8861 9939
rect 8861 9887 8913 9939
rect 8913 9887 8915 9939
rect 8859 9885 8915 9887
rect 9307 10593 9363 10595
rect 9307 10541 9309 10593
rect 9309 10541 9361 10593
rect 9361 10541 9363 10593
rect 9307 10539 9363 10541
rect 9307 10375 9363 10377
rect 9307 10323 9309 10375
rect 9309 10323 9361 10375
rect 9361 10323 9363 10375
rect 9307 10321 9363 10323
rect 9307 10157 9363 10159
rect 9307 10105 9309 10157
rect 9309 10105 9361 10157
rect 9361 10105 9363 10157
rect 9307 10103 9363 10105
rect 9307 9939 9363 9941
rect 9307 9887 9309 9939
rect 9309 9887 9361 9939
rect 9361 9887 9363 9939
rect 9307 9885 9363 9887
rect 9755 10593 9811 10595
rect 9755 10541 9757 10593
rect 9757 10541 9809 10593
rect 9809 10541 9811 10593
rect 9755 10539 9811 10541
rect 9755 10375 9811 10377
rect 9755 10323 9757 10375
rect 9757 10323 9809 10375
rect 9809 10323 9811 10375
rect 9755 10321 9811 10323
rect 9755 10157 9811 10159
rect 9755 10105 9757 10157
rect 9757 10105 9809 10157
rect 9809 10105 9811 10157
rect 9755 10103 9811 10105
rect 9755 9939 9811 9941
rect 9755 9887 9757 9939
rect 9757 9887 9809 9939
rect 9809 9887 9811 9939
rect 9755 9885 9811 9887
rect 10203 10593 10259 10595
rect 10203 10541 10205 10593
rect 10205 10541 10257 10593
rect 10257 10541 10259 10593
rect 10203 10539 10259 10541
rect 10203 10375 10259 10377
rect 10203 10323 10205 10375
rect 10205 10323 10257 10375
rect 10257 10323 10259 10375
rect 10203 10321 10259 10323
rect 10203 10157 10259 10159
rect 10203 10105 10205 10157
rect 10205 10105 10257 10157
rect 10257 10105 10259 10157
rect 10203 10103 10259 10105
rect 10203 9939 10259 9941
rect 10203 9887 10205 9939
rect 10205 9887 10257 9939
rect 10257 9887 10259 9939
rect 10203 9885 10259 9887
rect 10651 10593 10707 10595
rect 10651 10541 10653 10593
rect 10653 10541 10705 10593
rect 10705 10541 10707 10593
rect 10651 10539 10707 10541
rect 10651 10375 10707 10377
rect 10651 10323 10653 10375
rect 10653 10323 10705 10375
rect 10705 10323 10707 10375
rect 10651 10321 10707 10323
rect 10651 10157 10707 10159
rect 10651 10105 10653 10157
rect 10653 10105 10705 10157
rect 10705 10105 10707 10157
rect 10651 10103 10707 10105
rect 10651 9939 10707 9941
rect 10651 9887 10653 9939
rect 10653 9887 10705 9939
rect 10705 9887 10707 9939
rect 10651 9885 10707 9887
rect 11099 10593 11155 10595
rect 11099 10541 11101 10593
rect 11101 10541 11153 10593
rect 11153 10541 11155 10593
rect 11099 10539 11155 10541
rect 11099 10375 11155 10377
rect 11099 10323 11101 10375
rect 11101 10323 11153 10375
rect 11153 10323 11155 10375
rect 11099 10321 11155 10323
rect 11099 10157 11155 10159
rect 11099 10105 11101 10157
rect 11101 10105 11153 10157
rect 11153 10105 11155 10157
rect 11099 10103 11155 10105
rect 11099 9939 11155 9941
rect 11099 9887 11101 9939
rect 11101 9887 11153 9939
rect 11153 9887 11155 9939
rect 11099 9885 11155 9887
rect 11547 10593 11603 10595
rect 11547 10541 11549 10593
rect 11549 10541 11601 10593
rect 11601 10541 11603 10593
rect 11547 10539 11603 10541
rect 11547 10375 11603 10377
rect 11547 10323 11549 10375
rect 11549 10323 11601 10375
rect 11601 10323 11603 10375
rect 11547 10321 11603 10323
rect 11547 10157 11603 10159
rect 11547 10105 11549 10157
rect 11549 10105 11601 10157
rect 11601 10105 11603 10157
rect 11547 10103 11603 10105
rect 11547 9939 11603 9941
rect 11547 9887 11549 9939
rect 11549 9887 11601 9939
rect 11601 9887 11603 9939
rect 11547 9885 11603 9887
rect 11995 10593 12051 10595
rect 11995 10541 11997 10593
rect 11997 10541 12049 10593
rect 12049 10541 12051 10593
rect 11995 10539 12051 10541
rect 11995 10375 12051 10377
rect 11995 10323 11997 10375
rect 11997 10323 12049 10375
rect 12049 10323 12051 10375
rect 11995 10321 12051 10323
rect 11995 10157 12051 10159
rect 11995 10105 11997 10157
rect 11997 10105 12049 10157
rect 12049 10105 12051 10157
rect 11995 10103 12051 10105
rect 11995 9939 12051 9941
rect 11995 9887 11997 9939
rect 11997 9887 12049 9939
rect 12049 9887 12051 9939
rect 11995 9885 12051 9887
rect 12443 10593 12499 10595
rect 12443 10541 12445 10593
rect 12445 10541 12497 10593
rect 12497 10541 12499 10593
rect 12443 10539 12499 10541
rect 12443 10375 12499 10377
rect 12443 10323 12445 10375
rect 12445 10323 12497 10375
rect 12497 10323 12499 10375
rect 12443 10321 12499 10323
rect 12443 10157 12499 10159
rect 12443 10105 12445 10157
rect 12445 10105 12497 10157
rect 12497 10105 12499 10157
rect 12443 10103 12499 10105
rect 12443 9939 12499 9941
rect 12443 9887 12445 9939
rect 12445 9887 12497 9939
rect 12497 9887 12499 9939
rect 12443 9885 12499 9887
rect 12891 10593 12947 10595
rect 12891 10541 12893 10593
rect 12893 10541 12945 10593
rect 12945 10541 12947 10593
rect 12891 10539 12947 10541
rect 12891 10375 12947 10377
rect 12891 10323 12893 10375
rect 12893 10323 12945 10375
rect 12945 10323 12947 10375
rect 12891 10321 12947 10323
rect 12891 10157 12947 10159
rect 12891 10105 12893 10157
rect 12893 10105 12945 10157
rect 12945 10105 12947 10157
rect 12891 10103 12947 10105
rect 12891 9939 12947 9941
rect 12891 9887 12893 9939
rect 12893 9887 12945 9939
rect 12945 9887 12947 9939
rect 12891 9885 12947 9887
rect 13337 10593 13393 10595
rect 13337 10541 13339 10593
rect 13339 10541 13391 10593
rect 13391 10541 13393 10593
rect 13337 10539 13393 10541
rect 13337 10375 13393 10377
rect 13337 10323 13339 10375
rect 13339 10323 13391 10375
rect 13391 10323 13393 10375
rect 13337 10321 13393 10323
rect 13337 10157 13393 10159
rect 13337 10105 13339 10157
rect 13339 10105 13391 10157
rect 13391 10105 13393 10157
rect 13337 10103 13393 10105
rect 13337 9939 13393 9941
rect 13337 9887 13339 9939
rect 13339 9887 13391 9939
rect 13391 9887 13393 9939
rect 13337 9885 13393 9887
rect 13638 10627 13694 10629
rect 13638 10575 13640 10627
rect 13640 10575 13692 10627
rect 13692 10575 13694 10627
rect 13638 10573 13694 10575
rect 13638 10409 13694 10411
rect 13638 10357 13640 10409
rect 13640 10357 13692 10409
rect 13692 10357 13694 10409
rect 13638 10355 13694 10357
rect 13638 10191 13694 10193
rect 13638 10139 13640 10191
rect 13640 10139 13692 10191
rect 13692 10139 13694 10191
rect 13638 10137 13694 10139
rect 13638 9973 13694 9975
rect 13638 9921 13640 9973
rect 13640 9921 13692 9973
rect 13692 9921 13694 9973
rect 13638 9919 13694 9921
rect 6584 9163 6640 9219
rect 6796 9163 6852 9219
rect 6584 8945 6640 9001
rect 6796 8945 6852 9001
rect 4647 8704 4703 8760
rect 4859 8704 4915 8760
rect 455 8258 511 8260
rect 455 8206 457 8258
rect 457 8206 509 8258
rect 509 8206 511 8258
rect 455 8204 511 8206
rect 666 8258 722 8260
rect 666 8206 668 8258
rect 668 8206 720 8258
rect 720 8206 722 8258
rect 666 8204 722 8206
rect 876 8258 932 8260
rect 876 8206 878 8258
rect 878 8206 930 8258
rect 930 8206 932 8258
rect 876 8204 932 8206
rect 1087 8258 1143 8260
rect 1087 8206 1089 8258
rect 1089 8206 1141 8258
rect 1141 8206 1143 8258
rect 1087 8204 1143 8206
rect 1298 8258 1354 8260
rect 1298 8206 1300 8258
rect 1300 8206 1352 8258
rect 1352 8206 1354 8258
rect 1298 8204 1354 8206
rect 1509 8258 1565 8260
rect 1509 8206 1511 8258
rect 1511 8206 1563 8258
rect 1563 8206 1565 8258
rect 1509 8204 1565 8206
rect 1720 8258 1776 8260
rect 1720 8206 1722 8258
rect 1722 8206 1774 8258
rect 1774 8206 1776 8258
rect 1720 8204 1776 8206
rect 1930 8258 1986 8260
rect 1930 8206 1932 8258
rect 1932 8206 1984 8258
rect 1984 8206 1986 8258
rect 1930 8204 1986 8206
rect 2141 8258 2197 8260
rect 2141 8206 2143 8258
rect 2143 8206 2195 8258
rect 2195 8206 2197 8258
rect 2141 8204 2197 8206
rect 2353 8258 2409 8260
rect 2353 8206 2355 8258
rect 2355 8206 2407 8258
rect 2407 8206 2409 8258
rect 2353 8204 2409 8206
rect 2564 8258 2620 8260
rect 2564 8206 2566 8258
rect 2566 8206 2618 8258
rect 2618 8206 2620 8258
rect 2564 8204 2620 8206
rect 2774 8258 2830 8260
rect 2774 8206 2776 8258
rect 2776 8206 2828 8258
rect 2828 8206 2830 8258
rect 2774 8204 2830 8206
rect 2985 8258 3041 8260
rect 2985 8206 2987 8258
rect 2987 8206 3039 8258
rect 3039 8206 3041 8258
rect 2985 8204 3041 8206
rect 3196 8258 3252 8260
rect 3196 8206 3198 8258
rect 3198 8206 3250 8258
rect 3250 8206 3252 8258
rect 3196 8204 3252 8206
rect 3407 8258 3463 8260
rect 3407 8206 3409 8258
rect 3409 8206 3461 8258
rect 3461 8206 3463 8258
rect 3407 8204 3463 8206
rect 3618 8258 3674 8260
rect 3618 8206 3620 8258
rect 3620 8206 3672 8258
rect 3672 8206 3674 8258
rect 3618 8204 3674 8206
rect 3828 8258 3884 8260
rect 3828 8206 3830 8258
rect 3830 8206 3882 8258
rect 3882 8206 3884 8258
rect 3828 8204 3884 8206
rect 4039 8258 4095 8260
rect 4039 8206 4041 8258
rect 4041 8206 4093 8258
rect 4093 8206 4095 8258
rect 4039 8204 4095 8206
rect 455 8040 511 8042
rect 455 7988 457 8040
rect 457 7988 509 8040
rect 509 7988 511 8040
rect 455 7986 511 7988
rect 666 8040 722 8042
rect 666 7988 668 8040
rect 668 7988 720 8040
rect 720 7988 722 8040
rect 666 7986 722 7988
rect 876 8040 932 8042
rect 876 7988 878 8040
rect 878 7988 930 8040
rect 930 7988 932 8040
rect 876 7986 932 7988
rect 1087 8040 1143 8042
rect 1087 7988 1089 8040
rect 1089 7988 1141 8040
rect 1141 7988 1143 8040
rect 1087 7986 1143 7988
rect 1298 8040 1354 8042
rect 1298 7988 1300 8040
rect 1300 7988 1352 8040
rect 1352 7988 1354 8040
rect 1298 7986 1354 7988
rect 1509 8040 1565 8042
rect 1509 7988 1511 8040
rect 1511 7988 1563 8040
rect 1563 7988 1565 8040
rect 1509 7986 1565 7988
rect 1720 8040 1776 8042
rect 1720 7988 1722 8040
rect 1722 7988 1774 8040
rect 1774 7988 1776 8040
rect 1720 7986 1776 7988
rect 1930 8040 1986 8042
rect 1930 7988 1932 8040
rect 1932 7988 1984 8040
rect 1984 7988 1986 8040
rect 1930 7986 1986 7988
rect 2141 8040 2197 8042
rect 2141 7988 2143 8040
rect 2143 7988 2195 8040
rect 2195 7988 2197 8040
rect 2141 7986 2197 7988
rect 2353 8040 2409 8042
rect 2353 7988 2355 8040
rect 2355 7988 2407 8040
rect 2407 7988 2409 8040
rect 2353 7986 2409 7988
rect 2564 8040 2620 8042
rect 2564 7988 2566 8040
rect 2566 7988 2618 8040
rect 2618 7988 2620 8040
rect 2564 7986 2620 7988
rect 2774 8040 2830 8042
rect 2774 7988 2776 8040
rect 2776 7988 2828 8040
rect 2828 7988 2830 8040
rect 2774 7986 2830 7988
rect 2985 8040 3041 8042
rect 2985 7988 2987 8040
rect 2987 7988 3039 8040
rect 3039 7988 3041 8040
rect 2985 7986 3041 7988
rect 3196 8040 3252 8042
rect 3196 7988 3198 8040
rect 3198 7988 3250 8040
rect 3250 7988 3252 8040
rect 3196 7986 3252 7988
rect 3407 8040 3463 8042
rect 3407 7988 3409 8040
rect 3409 7988 3461 8040
rect 3461 7988 3463 8040
rect 3407 7986 3463 7988
rect 3618 8040 3674 8042
rect 3618 7988 3620 8040
rect 3620 7988 3672 8040
rect 3672 7988 3674 8040
rect 3618 7986 3674 7988
rect 3828 8040 3884 8042
rect 3828 7988 3830 8040
rect 3830 7988 3882 8040
rect 3882 7988 3884 8040
rect 3828 7986 3884 7988
rect 4039 8040 4095 8042
rect 4039 7988 4041 8040
rect 4041 7988 4093 8040
rect 4093 7988 4095 8040
rect 4039 7986 4095 7988
rect 455 7822 511 7824
rect 455 7770 457 7822
rect 457 7770 509 7822
rect 509 7770 511 7822
rect 455 7768 511 7770
rect 666 7822 722 7824
rect 666 7770 668 7822
rect 668 7770 720 7822
rect 720 7770 722 7822
rect 666 7768 722 7770
rect 876 7822 932 7824
rect 876 7770 878 7822
rect 878 7770 930 7822
rect 930 7770 932 7822
rect 876 7768 932 7770
rect 1087 7822 1143 7824
rect 1087 7770 1089 7822
rect 1089 7770 1141 7822
rect 1141 7770 1143 7822
rect 1087 7768 1143 7770
rect 1298 7822 1354 7824
rect 1298 7770 1300 7822
rect 1300 7770 1352 7822
rect 1352 7770 1354 7822
rect 1298 7768 1354 7770
rect 1509 7822 1565 7824
rect 1509 7770 1511 7822
rect 1511 7770 1563 7822
rect 1563 7770 1565 7822
rect 1509 7768 1565 7770
rect 1720 7822 1776 7824
rect 1720 7770 1722 7822
rect 1722 7770 1774 7822
rect 1774 7770 1776 7822
rect 1720 7768 1776 7770
rect 1930 7822 1986 7824
rect 1930 7770 1932 7822
rect 1932 7770 1984 7822
rect 1984 7770 1986 7822
rect 1930 7768 1986 7770
rect 2141 7822 2197 7824
rect 2141 7770 2143 7822
rect 2143 7770 2195 7822
rect 2195 7770 2197 7822
rect 2141 7768 2197 7770
rect 2353 7822 2409 7824
rect 2353 7770 2355 7822
rect 2355 7770 2407 7822
rect 2407 7770 2409 7822
rect 2353 7768 2409 7770
rect 2564 7822 2620 7824
rect 2564 7770 2566 7822
rect 2566 7770 2618 7822
rect 2618 7770 2620 7822
rect 2564 7768 2620 7770
rect 2774 7822 2830 7824
rect 2774 7770 2776 7822
rect 2776 7770 2828 7822
rect 2828 7770 2830 7822
rect 2774 7768 2830 7770
rect 2985 7822 3041 7824
rect 2985 7770 2987 7822
rect 2987 7770 3039 7822
rect 3039 7770 3041 7822
rect 2985 7768 3041 7770
rect 3196 7822 3252 7824
rect 3196 7770 3198 7822
rect 3198 7770 3250 7822
rect 3250 7770 3252 7822
rect 3196 7768 3252 7770
rect 3407 7822 3463 7824
rect 3407 7770 3409 7822
rect 3409 7770 3461 7822
rect 3461 7770 3463 7822
rect 3407 7768 3463 7770
rect 3618 7822 3674 7824
rect 3618 7770 3620 7822
rect 3620 7770 3672 7822
rect 3672 7770 3674 7822
rect 3618 7768 3674 7770
rect 3828 7822 3884 7824
rect 3828 7770 3830 7822
rect 3830 7770 3882 7822
rect 3882 7770 3884 7822
rect 3828 7768 3884 7770
rect 4039 7822 4095 7824
rect 4039 7770 4041 7822
rect 4041 7770 4093 7822
rect 4093 7770 4095 7822
rect 4039 7768 4095 7770
rect -283 7340 -227 7396
rect -71 7340 -15 7396
rect 741 6861 797 6863
rect 741 6809 743 6861
rect 743 6809 795 6861
rect 795 6809 797 6861
rect 741 6807 797 6809
rect 952 6861 1008 6863
rect 952 6809 954 6861
rect 954 6809 1006 6861
rect 1006 6809 1008 6861
rect 952 6807 1008 6809
rect 1162 6861 1218 6863
rect 1162 6809 1164 6861
rect 1164 6809 1216 6861
rect 1216 6809 1218 6861
rect 1162 6807 1218 6809
rect 1373 6861 1429 6863
rect 1373 6809 1375 6861
rect 1375 6809 1427 6861
rect 1427 6809 1429 6861
rect 1373 6807 1429 6809
rect 1584 6861 1640 6863
rect 1584 6809 1586 6861
rect 1586 6809 1638 6861
rect 1638 6809 1640 6861
rect 1584 6807 1640 6809
rect 1795 6861 1851 6863
rect 1795 6809 1797 6861
rect 1797 6809 1849 6861
rect 1849 6809 1851 6861
rect 1795 6807 1851 6809
rect 2006 6861 2062 6863
rect 2006 6809 2008 6861
rect 2008 6809 2060 6861
rect 2060 6809 2062 6861
rect 2006 6807 2062 6809
rect 2216 6861 2272 6863
rect 2216 6809 2218 6861
rect 2218 6809 2270 6861
rect 2270 6809 2272 6861
rect 2216 6807 2272 6809
rect 2427 6861 2483 6863
rect 2427 6809 2429 6861
rect 2429 6809 2481 6861
rect 2481 6809 2483 6861
rect 2427 6807 2483 6809
rect 2639 6861 2695 6863
rect 2639 6809 2641 6861
rect 2641 6809 2693 6861
rect 2693 6809 2695 6861
rect 2639 6807 2695 6809
rect 2850 6861 2906 6863
rect 2850 6809 2852 6861
rect 2852 6809 2904 6861
rect 2904 6809 2906 6861
rect 2850 6807 2906 6809
rect 3060 6861 3116 6863
rect 3060 6809 3062 6861
rect 3062 6809 3114 6861
rect 3114 6809 3116 6861
rect 3060 6807 3116 6809
rect 3271 6861 3327 6863
rect 3271 6809 3273 6861
rect 3273 6809 3325 6861
rect 3325 6809 3327 6861
rect 3271 6807 3327 6809
rect 3482 6861 3538 6863
rect 3482 6809 3484 6861
rect 3484 6809 3536 6861
rect 3536 6809 3538 6861
rect 3482 6807 3538 6809
rect 3693 6861 3749 6863
rect 3693 6809 3695 6861
rect 3695 6809 3747 6861
rect 3747 6809 3749 6861
rect 3693 6807 3749 6809
rect 3904 6861 3960 6863
rect 3904 6809 3906 6861
rect 3906 6809 3958 6861
rect 3958 6809 3960 6861
rect 3904 6807 3960 6809
rect 4114 6861 4170 6863
rect 4114 6809 4116 6861
rect 4116 6809 4168 6861
rect 4168 6809 4170 6861
rect 4114 6807 4170 6809
rect 4325 6861 4381 6863
rect 4325 6809 4327 6861
rect 4327 6809 4379 6861
rect 4379 6809 4381 6861
rect 4325 6807 4381 6809
rect 741 6643 797 6645
rect 741 6591 743 6643
rect 743 6591 795 6643
rect 795 6591 797 6643
rect 741 6589 797 6591
rect 952 6643 1008 6645
rect 952 6591 954 6643
rect 954 6591 1006 6643
rect 1006 6591 1008 6643
rect 952 6589 1008 6591
rect 1162 6643 1218 6645
rect 1162 6591 1164 6643
rect 1164 6591 1216 6643
rect 1216 6591 1218 6643
rect 1162 6589 1218 6591
rect 1373 6643 1429 6645
rect 1373 6591 1375 6643
rect 1375 6591 1427 6643
rect 1427 6591 1429 6643
rect 1373 6589 1429 6591
rect 1584 6643 1640 6645
rect 1584 6591 1586 6643
rect 1586 6591 1638 6643
rect 1638 6591 1640 6643
rect 1584 6589 1640 6591
rect 1795 6643 1851 6645
rect 1795 6591 1797 6643
rect 1797 6591 1849 6643
rect 1849 6591 1851 6643
rect 1795 6589 1851 6591
rect 2006 6643 2062 6645
rect 2006 6591 2008 6643
rect 2008 6591 2060 6643
rect 2060 6591 2062 6643
rect 2006 6589 2062 6591
rect 2216 6643 2272 6645
rect 2216 6591 2218 6643
rect 2218 6591 2270 6643
rect 2270 6591 2272 6643
rect 2216 6589 2272 6591
rect 2427 6643 2483 6645
rect 2427 6591 2429 6643
rect 2429 6591 2481 6643
rect 2481 6591 2483 6643
rect 2427 6589 2483 6591
rect 2639 6643 2695 6645
rect 2639 6591 2641 6643
rect 2641 6591 2693 6643
rect 2693 6591 2695 6643
rect 2639 6589 2695 6591
rect 2850 6643 2906 6645
rect 2850 6591 2852 6643
rect 2852 6591 2904 6643
rect 2904 6591 2906 6643
rect 2850 6589 2906 6591
rect 3060 6643 3116 6645
rect 3060 6591 3062 6643
rect 3062 6591 3114 6643
rect 3114 6591 3116 6643
rect 3060 6589 3116 6591
rect 3271 6643 3327 6645
rect 3271 6591 3273 6643
rect 3273 6591 3325 6643
rect 3325 6591 3327 6643
rect 3271 6589 3327 6591
rect 3482 6643 3538 6645
rect 3482 6591 3484 6643
rect 3484 6591 3536 6643
rect 3536 6591 3538 6643
rect 3482 6589 3538 6591
rect 3693 6643 3749 6645
rect 3693 6591 3695 6643
rect 3695 6591 3747 6643
rect 3747 6591 3749 6643
rect 3693 6589 3749 6591
rect 3904 6643 3960 6645
rect 3904 6591 3906 6643
rect 3906 6591 3958 6643
rect 3958 6591 3960 6643
rect 3904 6589 3960 6591
rect 4114 6643 4170 6645
rect 4114 6591 4116 6643
rect 4116 6591 4168 6643
rect 4168 6591 4170 6643
rect 4114 6589 4170 6591
rect 4325 6643 4381 6645
rect 4325 6591 4327 6643
rect 4327 6591 4379 6643
rect 4379 6591 4381 6643
rect 4325 6589 4381 6591
rect 5409 8471 5465 8527
rect 5621 8471 5677 8527
rect 7723 8471 7779 8527
rect 7935 8471 7991 8527
rect 7116 8153 7172 8155
rect 7116 8101 7118 8153
rect 7118 8101 7170 8153
rect 7170 8101 7172 8153
rect 7116 8099 7172 8101
rect 7116 7935 7172 7937
rect 7116 7883 7118 7935
rect 7118 7883 7170 7935
rect 7170 7883 7172 7935
rect 7116 7881 7172 7883
rect 8975 8395 9031 8397
rect 8975 8343 8977 8395
rect 8977 8343 9029 8395
rect 9029 8343 9031 8395
rect 8975 8341 9031 8343
rect 9187 8395 9243 8397
rect 9187 8343 9189 8395
rect 9189 8343 9241 8395
rect 9241 8343 9243 8395
rect 9187 8341 9243 8343
rect 8975 8178 9031 8180
rect 8975 8126 8977 8178
rect 8977 8126 9029 8178
rect 9029 8126 9031 8178
rect 8975 8124 9031 8126
rect 9187 8178 9243 8180
rect 9187 8126 9189 8178
rect 9189 8126 9241 8178
rect 9241 8126 9243 8178
rect 9187 8124 9243 8126
rect 8975 7960 9031 7962
rect 8975 7908 8977 7960
rect 8977 7908 9029 7960
rect 9029 7908 9031 7960
rect 8975 7906 9031 7908
rect 9187 7960 9243 7962
rect 9187 7908 9189 7960
rect 9189 7908 9241 7960
rect 9241 7908 9243 7960
rect 9187 7906 9243 7908
rect 8975 7743 9031 7745
rect 8975 7691 8977 7743
rect 8977 7691 9029 7743
rect 9029 7691 9031 7743
rect 8975 7689 9031 7691
rect 9187 7743 9243 7745
rect 9187 7691 9189 7743
rect 9189 7691 9241 7743
rect 9241 7691 9243 7743
rect 9187 7689 9243 7691
rect 4974 7065 5030 7067
rect 4974 7013 4976 7065
rect 4976 7013 5028 7065
rect 5028 7013 5030 7065
rect 4974 7011 5030 7013
rect 4974 6847 5030 6849
rect 4974 6795 4976 6847
rect 4976 6795 5028 6847
rect 5028 6795 5030 6847
rect 4974 6793 5030 6795
rect 4974 6629 5030 6631
rect 4974 6577 4976 6629
rect 4976 6577 5028 6629
rect 5028 6577 5030 6629
rect 4974 6575 5030 6577
rect 5677 7340 5733 7396
rect 5889 7340 5945 7396
rect 741 5877 797 5879
rect 741 5825 743 5877
rect 743 5825 795 5877
rect 795 5825 797 5877
rect 741 5823 797 5825
rect 952 5877 1008 5879
rect 952 5825 954 5877
rect 954 5825 1006 5877
rect 1006 5825 1008 5877
rect 952 5823 1008 5825
rect 1162 5877 1218 5879
rect 1162 5825 1164 5877
rect 1164 5825 1216 5877
rect 1216 5825 1218 5877
rect 1162 5823 1218 5825
rect 1373 5877 1429 5879
rect 1373 5825 1375 5877
rect 1375 5825 1427 5877
rect 1427 5825 1429 5877
rect 1373 5823 1429 5825
rect 1584 5877 1640 5879
rect 1584 5825 1586 5877
rect 1586 5825 1638 5877
rect 1638 5825 1640 5877
rect 1584 5823 1640 5825
rect 1795 5877 1851 5879
rect 1795 5825 1797 5877
rect 1797 5825 1849 5877
rect 1849 5825 1851 5877
rect 1795 5823 1851 5825
rect 2006 5877 2062 5879
rect 2006 5825 2008 5877
rect 2008 5825 2060 5877
rect 2060 5825 2062 5877
rect 2006 5823 2062 5825
rect 2216 5877 2272 5879
rect 2216 5825 2218 5877
rect 2218 5825 2270 5877
rect 2270 5825 2272 5877
rect 2216 5823 2272 5825
rect 2427 5877 2483 5879
rect 2427 5825 2429 5877
rect 2429 5825 2481 5877
rect 2481 5825 2483 5877
rect 2427 5823 2483 5825
rect 2639 5877 2695 5879
rect 2639 5825 2641 5877
rect 2641 5825 2693 5877
rect 2693 5825 2695 5877
rect 2639 5823 2695 5825
rect 2850 5877 2906 5879
rect 2850 5825 2852 5877
rect 2852 5825 2904 5877
rect 2904 5825 2906 5877
rect 2850 5823 2906 5825
rect 3060 5877 3116 5879
rect 3060 5825 3062 5877
rect 3062 5825 3114 5877
rect 3114 5825 3116 5877
rect 3060 5823 3116 5825
rect 3271 5877 3327 5879
rect 3271 5825 3273 5877
rect 3273 5825 3325 5877
rect 3325 5825 3327 5877
rect 3271 5823 3327 5825
rect 3482 5877 3538 5879
rect 3482 5825 3484 5877
rect 3484 5825 3536 5877
rect 3536 5825 3538 5877
rect 3482 5823 3538 5825
rect 3693 5877 3749 5879
rect 3693 5825 3695 5877
rect 3695 5825 3747 5877
rect 3747 5825 3749 5877
rect 3693 5823 3749 5825
rect 3904 5877 3960 5879
rect 3904 5825 3906 5877
rect 3906 5825 3958 5877
rect 3958 5825 3960 5877
rect 3904 5823 3960 5825
rect 4114 5877 4170 5879
rect 4114 5825 4116 5877
rect 4116 5825 4168 5877
rect 4168 5825 4170 5877
rect 4114 5823 4170 5825
rect 4325 5877 4381 5879
rect 4325 5825 4327 5877
rect 4327 5825 4379 5877
rect 4379 5825 4381 5877
rect 4325 5823 4381 5825
rect 8975 7525 9031 7527
rect 8975 7473 8977 7525
rect 8977 7473 9029 7525
rect 9029 7473 9031 7525
rect 8975 7471 9031 7473
rect 9187 7525 9243 7527
rect 9187 7473 9189 7525
rect 9189 7473 9241 7525
rect 9241 7473 9243 7525
rect 9187 7471 9243 7473
rect 8975 7307 9031 7309
rect 8975 7255 8977 7307
rect 8977 7255 9029 7307
rect 9029 7255 9031 7307
rect 8975 7253 9031 7255
rect 9187 7307 9243 7309
rect 9187 7255 9189 7307
rect 9189 7255 9241 7307
rect 9241 7255 9243 7307
rect 9187 7253 9243 7255
rect 7116 7075 7172 7077
rect 7116 7023 7118 7075
rect 7118 7023 7170 7075
rect 7170 7023 7172 7075
rect 7116 7021 7172 7023
rect 6384 6857 6440 6859
rect 6384 6805 6386 6857
rect 6386 6805 6438 6857
rect 6438 6805 6440 6857
rect 6384 6803 6440 6805
rect 6384 6639 6440 6641
rect 6384 6587 6386 6639
rect 6386 6587 6438 6639
rect 6438 6587 6440 6639
rect 6384 6585 6440 6587
rect 6384 6421 6440 6423
rect 6384 6369 6386 6421
rect 6386 6369 6438 6421
rect 6438 6369 6440 6421
rect 6384 6367 6440 6369
rect 7116 6857 7172 6859
rect 7116 6805 7118 6857
rect 7118 6805 7170 6857
rect 7170 6805 7172 6857
rect 7116 6803 7172 6805
rect 7116 6639 7172 6641
rect 7116 6587 7118 6639
rect 7118 6587 7170 6639
rect 7170 6587 7172 6639
rect 7116 6585 7172 6587
rect 7116 6421 7172 6423
rect 7116 6369 7118 6421
rect 7118 6369 7170 6421
rect 7170 6369 7172 6421
rect 7116 6367 7172 6369
rect 8975 7089 9031 7091
rect 8975 7037 8977 7089
rect 8977 7037 9029 7089
rect 9029 7037 9031 7089
rect 8975 7035 9031 7037
rect 9187 7089 9243 7091
rect 9187 7037 9189 7089
rect 9189 7037 9241 7089
rect 9241 7037 9243 7089
rect 9187 7035 9243 7037
rect 8975 6872 9031 6874
rect 8975 6820 8977 6872
rect 8977 6820 9029 6872
rect 9029 6820 9031 6872
rect 8975 6818 9031 6820
rect 9187 6872 9243 6874
rect 9187 6820 9189 6872
rect 9189 6820 9241 6872
rect 9241 6820 9243 6872
rect 9187 6818 9243 6820
rect 8975 6654 9031 6656
rect 8975 6602 8977 6654
rect 8977 6602 9029 6654
rect 9029 6602 9031 6654
rect 8975 6600 9031 6602
rect 9187 6654 9243 6656
rect 9187 6602 9189 6654
rect 9189 6602 9241 6654
rect 9241 6602 9243 6654
rect 9187 6600 9243 6602
rect 8975 6437 9031 6439
rect 8975 6385 8977 6437
rect 8977 6385 9029 6437
rect 9029 6385 9031 6437
rect 8975 6383 9031 6385
rect 9187 6437 9243 6439
rect 9187 6385 9189 6437
rect 9189 6385 9241 6437
rect 9241 6385 9243 6437
rect 9187 6383 9243 6385
rect 9446 8395 9502 8397
rect 9446 8343 9448 8395
rect 9448 8343 9500 8395
rect 9500 8343 9502 8395
rect 9446 8341 9502 8343
rect 9446 8178 9502 8180
rect 9446 8126 9448 8178
rect 9448 8126 9500 8178
rect 9500 8126 9502 8178
rect 9446 8124 9502 8126
rect 9446 7960 9502 7962
rect 9446 7908 9448 7960
rect 9448 7908 9500 7960
rect 9500 7908 9502 7960
rect 9446 7906 9502 7908
rect 9446 7743 9502 7745
rect 9446 7691 9448 7743
rect 9448 7691 9500 7743
rect 9500 7691 9502 7743
rect 9446 7689 9502 7691
rect 9446 7525 9502 7527
rect 9446 7473 9448 7525
rect 9448 7473 9500 7525
rect 9500 7473 9502 7525
rect 9446 7471 9502 7473
rect 9446 7307 9502 7309
rect 9446 7255 9448 7307
rect 9448 7255 9500 7307
rect 9500 7255 9502 7307
rect 9446 7253 9502 7255
rect 9446 7089 9502 7091
rect 9446 7037 9448 7089
rect 9448 7037 9500 7089
rect 9500 7037 9502 7089
rect 9446 7035 9502 7037
rect 9446 6872 9502 6874
rect 9446 6820 9448 6872
rect 9448 6820 9500 6872
rect 9500 6820 9502 6872
rect 9446 6818 9502 6820
rect 9446 6654 9502 6656
rect 9446 6602 9448 6654
rect 9448 6602 9500 6654
rect 9500 6602 9502 6654
rect 9446 6600 9502 6602
rect 9446 6437 9502 6439
rect 9446 6385 9448 6437
rect 9448 6385 9500 6437
rect 9500 6385 9502 6437
rect 9446 6383 9502 6385
rect 9894 8395 9950 8397
rect 9894 8343 9896 8395
rect 9896 8343 9948 8395
rect 9948 8343 9950 8395
rect 9894 8341 9950 8343
rect 9894 8178 9950 8180
rect 9894 8126 9896 8178
rect 9896 8126 9948 8178
rect 9948 8126 9950 8178
rect 9894 8124 9950 8126
rect 9894 7960 9950 7962
rect 9894 7908 9896 7960
rect 9896 7908 9948 7960
rect 9948 7908 9950 7960
rect 9894 7906 9950 7908
rect 9894 7743 9950 7745
rect 9894 7691 9896 7743
rect 9896 7691 9948 7743
rect 9948 7691 9950 7743
rect 9894 7689 9950 7691
rect 9894 7525 9950 7527
rect 9894 7473 9896 7525
rect 9896 7473 9948 7525
rect 9948 7473 9950 7525
rect 9894 7471 9950 7473
rect 9894 7307 9950 7309
rect 9894 7255 9896 7307
rect 9896 7255 9948 7307
rect 9948 7255 9950 7307
rect 9894 7253 9950 7255
rect 9894 7089 9950 7091
rect 9894 7037 9896 7089
rect 9896 7037 9948 7089
rect 9948 7037 9950 7089
rect 9894 7035 9950 7037
rect 9894 6872 9950 6874
rect 9894 6820 9896 6872
rect 9896 6820 9948 6872
rect 9948 6820 9950 6872
rect 9894 6818 9950 6820
rect 9894 6654 9950 6656
rect 9894 6602 9896 6654
rect 9896 6602 9948 6654
rect 9948 6602 9950 6654
rect 9894 6600 9950 6602
rect 9894 6437 9950 6439
rect 9894 6385 9896 6437
rect 9896 6385 9948 6437
rect 9948 6385 9950 6437
rect 9894 6383 9950 6385
rect 741 5659 797 5661
rect 741 5607 743 5659
rect 743 5607 795 5659
rect 795 5607 797 5659
rect 741 5605 797 5607
rect 952 5659 1008 5661
rect 952 5607 954 5659
rect 954 5607 1006 5659
rect 1006 5607 1008 5659
rect 952 5605 1008 5607
rect 1162 5659 1218 5661
rect 1162 5607 1164 5659
rect 1164 5607 1216 5659
rect 1216 5607 1218 5659
rect 1162 5605 1218 5607
rect 1373 5659 1429 5661
rect 1373 5607 1375 5659
rect 1375 5607 1427 5659
rect 1427 5607 1429 5659
rect 1373 5605 1429 5607
rect 1584 5659 1640 5661
rect 1584 5607 1586 5659
rect 1586 5607 1638 5659
rect 1638 5607 1640 5659
rect 1584 5605 1640 5607
rect 1795 5659 1851 5661
rect 1795 5607 1797 5659
rect 1797 5607 1849 5659
rect 1849 5607 1851 5659
rect 1795 5605 1851 5607
rect 2006 5659 2062 5661
rect 2006 5607 2008 5659
rect 2008 5607 2060 5659
rect 2060 5607 2062 5659
rect 2006 5605 2062 5607
rect 2216 5659 2272 5661
rect 2216 5607 2218 5659
rect 2218 5607 2270 5659
rect 2270 5607 2272 5659
rect 2216 5605 2272 5607
rect 2427 5659 2483 5661
rect 2427 5607 2429 5659
rect 2429 5607 2481 5659
rect 2481 5607 2483 5659
rect 2427 5605 2483 5607
rect 2639 5659 2695 5661
rect 2639 5607 2641 5659
rect 2641 5607 2693 5659
rect 2693 5607 2695 5659
rect 2639 5605 2695 5607
rect 2850 5659 2906 5661
rect 2850 5607 2852 5659
rect 2852 5607 2904 5659
rect 2904 5607 2906 5659
rect 2850 5605 2906 5607
rect 3060 5659 3116 5661
rect 3060 5607 3062 5659
rect 3062 5607 3114 5659
rect 3114 5607 3116 5659
rect 3060 5605 3116 5607
rect 3271 5659 3327 5661
rect 3271 5607 3273 5659
rect 3273 5607 3325 5659
rect 3325 5607 3327 5659
rect 3271 5605 3327 5607
rect 3482 5659 3538 5661
rect 3482 5607 3484 5659
rect 3484 5607 3536 5659
rect 3536 5607 3538 5659
rect 3482 5605 3538 5607
rect 3693 5659 3749 5661
rect 3693 5607 3695 5659
rect 3695 5607 3747 5659
rect 3747 5607 3749 5659
rect 3693 5605 3749 5607
rect 3904 5659 3960 5661
rect 3904 5607 3906 5659
rect 3906 5607 3958 5659
rect 3958 5607 3960 5659
rect 3904 5605 3960 5607
rect 4114 5659 4170 5661
rect 4114 5607 4116 5659
rect 4116 5607 4168 5659
rect 4168 5607 4170 5659
rect 4114 5605 4170 5607
rect 4325 5659 4381 5661
rect 4325 5607 4327 5659
rect 4327 5607 4379 5659
rect 4379 5607 4381 5659
rect 4325 5605 4381 5607
rect 5198 5626 5254 5628
rect 5198 5574 5200 5626
rect 5200 5574 5252 5626
rect 5252 5574 5254 5626
rect 5198 5572 5254 5574
rect 5198 5408 5254 5410
rect 5198 5356 5200 5408
rect 5200 5356 5252 5408
rect 5252 5356 5254 5408
rect 5198 5354 5254 5356
rect 6384 5970 6440 5972
rect 6384 5918 6386 5970
rect 6386 5918 6438 5970
rect 6438 5918 6440 5970
rect 6384 5916 6440 5918
rect 6384 5752 6440 5754
rect 6384 5700 6386 5752
rect 6386 5700 6438 5752
rect 6438 5700 6440 5752
rect 6384 5698 6440 5700
rect 253 4937 309 4939
rect 253 4885 255 4937
rect 255 4885 307 4937
rect 307 4885 309 4937
rect 253 4883 309 4885
rect 464 4937 520 4939
rect 464 4885 466 4937
rect 466 4885 518 4937
rect 518 4885 520 4937
rect 464 4883 520 4885
rect 675 4937 731 4939
rect 675 4885 677 4937
rect 677 4885 729 4937
rect 729 4885 731 4937
rect 675 4883 731 4885
rect 885 4937 941 4939
rect 885 4885 887 4937
rect 887 4885 939 4937
rect 939 4885 941 4937
rect 885 4883 941 4885
rect 1096 4937 1152 4939
rect 1096 4885 1098 4937
rect 1098 4885 1150 4937
rect 1150 4885 1152 4937
rect 1096 4883 1152 4885
rect 1307 4937 1363 4939
rect 1307 4885 1309 4937
rect 1309 4885 1361 4937
rect 1361 4885 1363 4937
rect 1307 4883 1363 4885
rect 1518 4937 1574 4939
rect 1518 4885 1520 4937
rect 1520 4885 1572 4937
rect 1572 4885 1574 4937
rect 1518 4883 1574 4885
rect 1729 4937 1785 4939
rect 1729 4885 1731 4937
rect 1731 4885 1783 4937
rect 1783 4885 1785 4937
rect 1729 4883 1785 4885
rect 1939 4937 1995 4939
rect 1939 4885 1941 4937
rect 1941 4885 1993 4937
rect 1993 4885 1995 4937
rect 1939 4883 1995 4885
rect 2150 4937 2206 4939
rect 2150 4885 2152 4937
rect 2152 4885 2204 4937
rect 2204 4885 2206 4937
rect 2150 4883 2206 4885
rect 2361 4937 2417 4939
rect 2361 4885 2363 4937
rect 2363 4885 2415 4937
rect 2415 4885 2417 4937
rect 2361 4883 2417 4885
rect 2572 4937 2628 4939
rect 2572 4885 2574 4937
rect 2574 4885 2626 4937
rect 2626 4885 2628 4937
rect 2572 4883 2628 4885
rect 2783 4937 2839 4939
rect 2783 4885 2785 4937
rect 2785 4885 2837 4937
rect 2837 4885 2839 4937
rect 2783 4883 2839 4885
rect 2994 4937 3050 4939
rect 2994 4885 2996 4937
rect 2996 4885 3048 4937
rect 3048 4885 3050 4937
rect 2994 4883 3050 4885
rect 3205 4937 3261 4939
rect 3205 4885 3207 4937
rect 3207 4885 3259 4937
rect 3259 4885 3261 4937
rect 3205 4883 3261 4885
rect 3416 4937 3472 4939
rect 3416 4885 3418 4937
rect 3418 4885 3470 4937
rect 3470 4885 3472 4937
rect 3416 4883 3472 4885
rect 3627 4937 3683 4939
rect 3627 4885 3629 4937
rect 3629 4885 3681 4937
rect 3681 4885 3683 4937
rect 3627 4883 3683 4885
rect 3837 4937 3893 4939
rect 3837 4885 3839 4937
rect 3839 4885 3891 4937
rect 3891 4885 3893 4937
rect 3837 4883 3893 4885
rect 4048 4937 4104 4939
rect 4048 4885 4050 4937
rect 4050 4885 4102 4937
rect 4102 4885 4104 4937
rect 4048 4883 4104 4885
rect 4259 4937 4315 4939
rect 4259 4885 4261 4937
rect 4261 4885 4313 4937
rect 4313 4885 4315 4937
rect 4259 4883 4315 4885
rect 4470 4937 4526 4939
rect 4470 4885 4472 4937
rect 4472 4885 4524 4937
rect 4524 4885 4526 4937
rect 4470 4883 4526 4885
rect 4681 4937 4737 4939
rect 4681 4885 4683 4937
rect 4683 4885 4735 4937
rect 4735 4885 4737 4937
rect 4681 4883 4737 4885
rect 4891 4937 4947 4939
rect 4891 4885 4893 4937
rect 4893 4885 4945 4937
rect 4945 4885 4947 4937
rect 4891 4883 4947 4885
rect 5102 4937 5158 4939
rect 5102 4885 5104 4937
rect 5104 4885 5156 4937
rect 5156 4885 5158 4937
rect 5102 4883 5158 4885
rect 5313 4937 5369 4939
rect 5313 4885 5315 4937
rect 5315 4885 5367 4937
rect 5367 4885 5369 4937
rect 5313 4883 5369 4885
rect 253 4719 309 4721
rect 253 4667 255 4719
rect 255 4667 307 4719
rect 307 4667 309 4719
rect 253 4665 309 4667
rect 464 4719 520 4721
rect 464 4667 466 4719
rect 466 4667 518 4719
rect 518 4667 520 4719
rect 464 4665 520 4667
rect 675 4719 731 4721
rect 675 4667 677 4719
rect 677 4667 729 4719
rect 729 4667 731 4719
rect 675 4665 731 4667
rect 885 4719 941 4721
rect 885 4667 887 4719
rect 887 4667 939 4719
rect 939 4667 941 4719
rect 885 4665 941 4667
rect 1096 4719 1152 4721
rect 1096 4667 1098 4719
rect 1098 4667 1150 4719
rect 1150 4667 1152 4719
rect 1096 4665 1152 4667
rect 1307 4719 1363 4721
rect 1307 4667 1309 4719
rect 1309 4667 1361 4719
rect 1361 4667 1363 4719
rect 1307 4665 1363 4667
rect 1518 4719 1574 4721
rect 1518 4667 1520 4719
rect 1520 4667 1572 4719
rect 1572 4667 1574 4719
rect 1518 4665 1574 4667
rect 1729 4719 1785 4721
rect 1729 4667 1731 4719
rect 1731 4667 1783 4719
rect 1783 4667 1785 4719
rect 1729 4665 1785 4667
rect 1939 4719 1995 4721
rect 1939 4667 1941 4719
rect 1941 4667 1993 4719
rect 1993 4667 1995 4719
rect 1939 4665 1995 4667
rect 2150 4719 2206 4721
rect 2150 4667 2152 4719
rect 2152 4667 2204 4719
rect 2204 4667 2206 4719
rect 2150 4665 2206 4667
rect 2361 4719 2417 4721
rect 2361 4667 2363 4719
rect 2363 4667 2415 4719
rect 2415 4667 2417 4719
rect 2361 4665 2417 4667
rect 2572 4719 2628 4721
rect 2572 4667 2574 4719
rect 2574 4667 2626 4719
rect 2626 4667 2628 4719
rect 2572 4665 2628 4667
rect 2783 4719 2839 4721
rect 2783 4667 2785 4719
rect 2785 4667 2837 4719
rect 2837 4667 2839 4719
rect 2783 4665 2839 4667
rect 2994 4719 3050 4721
rect 2994 4667 2996 4719
rect 2996 4667 3048 4719
rect 3048 4667 3050 4719
rect 2994 4665 3050 4667
rect 3205 4719 3261 4721
rect 3205 4667 3207 4719
rect 3207 4667 3259 4719
rect 3259 4667 3261 4719
rect 3205 4665 3261 4667
rect 3416 4719 3472 4721
rect 3416 4667 3418 4719
rect 3418 4667 3470 4719
rect 3470 4667 3472 4719
rect 3416 4665 3472 4667
rect 3627 4719 3683 4721
rect 3627 4667 3629 4719
rect 3629 4667 3681 4719
rect 3681 4667 3683 4719
rect 3627 4665 3683 4667
rect 3837 4719 3893 4721
rect 3837 4667 3839 4719
rect 3839 4667 3891 4719
rect 3891 4667 3893 4719
rect 3837 4665 3893 4667
rect 4048 4719 4104 4721
rect 4048 4667 4050 4719
rect 4050 4667 4102 4719
rect 4102 4667 4104 4719
rect 4048 4665 4104 4667
rect 4259 4719 4315 4721
rect 4259 4667 4261 4719
rect 4261 4667 4313 4719
rect 4313 4667 4315 4719
rect 4259 4665 4315 4667
rect 4470 4719 4526 4721
rect 4470 4667 4472 4719
rect 4472 4667 4524 4719
rect 4524 4667 4526 4719
rect 4470 4665 4526 4667
rect 4681 4719 4737 4721
rect 4681 4667 4683 4719
rect 4683 4667 4735 4719
rect 4735 4667 4737 4719
rect 4681 4665 4737 4667
rect 4891 4719 4947 4721
rect 4891 4667 4893 4719
rect 4893 4667 4945 4719
rect 4945 4667 4947 4719
rect 4891 4665 4947 4667
rect 5102 4719 5158 4721
rect 5102 4667 5104 4719
rect 5104 4667 5156 4719
rect 5156 4667 5158 4719
rect 5102 4665 5158 4667
rect 5313 4719 5369 4721
rect 5313 4667 5315 4719
rect 5315 4667 5367 4719
rect 5367 4667 5369 4719
rect 5313 4665 5369 4667
rect 253 4501 309 4503
rect 253 4449 255 4501
rect 255 4449 307 4501
rect 307 4449 309 4501
rect 253 4447 309 4449
rect 464 4501 520 4503
rect 464 4449 466 4501
rect 466 4449 518 4501
rect 518 4449 520 4501
rect 464 4447 520 4449
rect 675 4501 731 4503
rect 675 4449 677 4501
rect 677 4449 729 4501
rect 729 4449 731 4501
rect 675 4447 731 4449
rect 885 4501 941 4503
rect 885 4449 887 4501
rect 887 4449 939 4501
rect 939 4449 941 4501
rect 885 4447 941 4449
rect 1096 4501 1152 4503
rect 1096 4449 1098 4501
rect 1098 4449 1150 4501
rect 1150 4449 1152 4501
rect 1096 4447 1152 4449
rect 1307 4501 1363 4503
rect 1307 4449 1309 4501
rect 1309 4449 1361 4501
rect 1361 4449 1363 4501
rect 1307 4447 1363 4449
rect 1518 4501 1574 4503
rect 1518 4449 1520 4501
rect 1520 4449 1572 4501
rect 1572 4449 1574 4501
rect 1518 4447 1574 4449
rect 1729 4501 1785 4503
rect 1729 4449 1731 4501
rect 1731 4449 1783 4501
rect 1783 4449 1785 4501
rect 1729 4447 1785 4449
rect 1939 4501 1995 4503
rect 1939 4449 1941 4501
rect 1941 4449 1993 4501
rect 1993 4449 1995 4501
rect 1939 4447 1995 4449
rect 2150 4501 2206 4503
rect 2150 4449 2152 4501
rect 2152 4449 2204 4501
rect 2204 4449 2206 4501
rect 2150 4447 2206 4449
rect 2361 4501 2417 4503
rect 2361 4449 2363 4501
rect 2363 4449 2415 4501
rect 2415 4449 2417 4501
rect 2361 4447 2417 4449
rect 2572 4501 2628 4503
rect 2572 4449 2574 4501
rect 2574 4449 2626 4501
rect 2626 4449 2628 4501
rect 2572 4447 2628 4449
rect 2783 4501 2839 4503
rect 2783 4449 2785 4501
rect 2785 4449 2837 4501
rect 2837 4449 2839 4501
rect 2783 4447 2839 4449
rect 2994 4501 3050 4503
rect 2994 4449 2996 4501
rect 2996 4449 3048 4501
rect 3048 4449 3050 4501
rect 2994 4447 3050 4449
rect 3205 4501 3261 4503
rect 3205 4449 3207 4501
rect 3207 4449 3259 4501
rect 3259 4449 3261 4501
rect 3205 4447 3261 4449
rect 3416 4501 3472 4503
rect 3416 4449 3418 4501
rect 3418 4449 3470 4501
rect 3470 4449 3472 4501
rect 3416 4447 3472 4449
rect 3627 4501 3683 4503
rect 3627 4449 3629 4501
rect 3629 4449 3681 4501
rect 3681 4449 3683 4501
rect 3627 4447 3683 4449
rect 3837 4501 3893 4503
rect 3837 4449 3839 4501
rect 3839 4449 3891 4501
rect 3891 4449 3893 4501
rect 3837 4447 3893 4449
rect 4048 4501 4104 4503
rect 4048 4449 4050 4501
rect 4050 4449 4102 4501
rect 4102 4449 4104 4501
rect 4048 4447 4104 4449
rect 4259 4501 4315 4503
rect 4259 4449 4261 4501
rect 4261 4449 4313 4501
rect 4313 4449 4315 4501
rect 4259 4447 4315 4449
rect 4470 4501 4526 4503
rect 4470 4449 4472 4501
rect 4472 4449 4524 4501
rect 4524 4449 4526 4501
rect 4470 4447 4526 4449
rect 4681 4501 4737 4503
rect 4681 4449 4683 4501
rect 4683 4449 4735 4501
rect 4735 4449 4737 4501
rect 4681 4447 4737 4449
rect 4891 4501 4947 4503
rect 4891 4449 4893 4501
rect 4893 4449 4945 4501
rect 4945 4449 4947 4501
rect 4891 4447 4947 4449
rect 5102 4501 5158 4503
rect 5102 4449 5104 4501
rect 5104 4449 5156 4501
rect 5156 4449 5158 4501
rect 5102 4447 5158 4449
rect 5313 4501 5369 4503
rect 5313 4449 5315 4501
rect 5315 4449 5367 4501
rect 5367 4449 5369 4501
rect 5313 4447 5369 4449
rect 253 4283 309 4285
rect 253 4231 255 4283
rect 255 4231 307 4283
rect 307 4231 309 4283
rect 253 4229 309 4231
rect 464 4283 520 4285
rect 464 4231 466 4283
rect 466 4231 518 4283
rect 518 4231 520 4283
rect 464 4229 520 4231
rect 675 4283 731 4285
rect 675 4231 677 4283
rect 677 4231 729 4283
rect 729 4231 731 4283
rect 675 4229 731 4231
rect 885 4283 941 4285
rect 885 4231 887 4283
rect 887 4231 939 4283
rect 939 4231 941 4283
rect 885 4229 941 4231
rect 1096 4283 1152 4285
rect 1096 4231 1098 4283
rect 1098 4231 1150 4283
rect 1150 4231 1152 4283
rect 1096 4229 1152 4231
rect 1307 4283 1363 4285
rect 1307 4231 1309 4283
rect 1309 4231 1361 4283
rect 1361 4231 1363 4283
rect 1307 4229 1363 4231
rect 1518 4283 1574 4285
rect 1518 4231 1520 4283
rect 1520 4231 1572 4283
rect 1572 4231 1574 4283
rect 1518 4229 1574 4231
rect 1729 4283 1785 4285
rect 1729 4231 1731 4283
rect 1731 4231 1783 4283
rect 1783 4231 1785 4283
rect 1729 4229 1785 4231
rect 1939 4283 1995 4285
rect 1939 4231 1941 4283
rect 1941 4231 1993 4283
rect 1993 4231 1995 4283
rect 1939 4229 1995 4231
rect 2150 4283 2206 4285
rect 2150 4231 2152 4283
rect 2152 4231 2204 4283
rect 2204 4231 2206 4283
rect 2150 4229 2206 4231
rect 2361 4283 2417 4285
rect 2361 4231 2363 4283
rect 2363 4231 2415 4283
rect 2415 4231 2417 4283
rect 2361 4229 2417 4231
rect 2572 4283 2628 4285
rect 2572 4231 2574 4283
rect 2574 4231 2626 4283
rect 2626 4231 2628 4283
rect 2572 4229 2628 4231
rect 2783 4283 2839 4285
rect 2783 4231 2785 4283
rect 2785 4231 2837 4283
rect 2837 4231 2839 4283
rect 2783 4229 2839 4231
rect 2994 4283 3050 4285
rect 2994 4231 2996 4283
rect 2996 4231 3048 4283
rect 3048 4231 3050 4283
rect 2994 4229 3050 4231
rect 3205 4283 3261 4285
rect 3205 4231 3207 4283
rect 3207 4231 3259 4283
rect 3259 4231 3261 4283
rect 3205 4229 3261 4231
rect 3416 4283 3472 4285
rect 3416 4231 3418 4283
rect 3418 4231 3470 4283
rect 3470 4231 3472 4283
rect 3416 4229 3472 4231
rect 3627 4283 3683 4285
rect 3627 4231 3629 4283
rect 3629 4231 3681 4283
rect 3681 4231 3683 4283
rect 3627 4229 3683 4231
rect 3837 4283 3893 4285
rect 3837 4231 3839 4283
rect 3839 4231 3891 4283
rect 3891 4231 3893 4283
rect 3837 4229 3893 4231
rect 4048 4283 4104 4285
rect 4048 4231 4050 4283
rect 4050 4231 4102 4283
rect 4102 4231 4104 4283
rect 4048 4229 4104 4231
rect 4259 4283 4315 4285
rect 4259 4231 4261 4283
rect 4261 4231 4313 4283
rect 4313 4231 4315 4283
rect 4259 4229 4315 4231
rect 4470 4283 4526 4285
rect 4470 4231 4472 4283
rect 4472 4231 4524 4283
rect 4524 4231 4526 4283
rect 4470 4229 4526 4231
rect 4681 4283 4737 4285
rect 4681 4231 4683 4283
rect 4683 4231 4735 4283
rect 4735 4231 4737 4283
rect 4681 4229 4737 4231
rect 4891 4283 4947 4285
rect 4891 4231 4893 4283
rect 4893 4231 4945 4283
rect 4945 4231 4947 4283
rect 4891 4229 4947 4231
rect 5102 4283 5158 4285
rect 5102 4231 5104 4283
rect 5104 4231 5156 4283
rect 5156 4231 5158 4283
rect 5102 4229 5158 4231
rect 5313 4283 5369 4285
rect 5313 4231 5315 4283
rect 5315 4231 5367 4283
rect 5367 4231 5369 4283
rect 5313 4229 5369 4231
rect 2524 2730 2580 2732
rect 2524 2678 2526 2730
rect 2526 2678 2578 2730
rect 2578 2678 2580 2730
rect 2524 2676 2580 2678
rect 2656 2730 2712 2732
rect 2656 2678 2658 2730
rect 2658 2678 2710 2730
rect 2710 2678 2712 2730
rect 2656 2676 2712 2678
rect 2788 2730 2844 2732
rect 2788 2678 2790 2730
rect 2790 2678 2842 2730
rect 2842 2678 2844 2730
rect 2788 2676 2844 2678
rect 2920 2730 2976 2732
rect 2920 2678 2922 2730
rect 2922 2678 2974 2730
rect 2974 2678 2976 2730
rect 2920 2676 2976 2678
rect 3052 2730 3108 2732
rect 3052 2678 3054 2730
rect 3054 2678 3106 2730
rect 3106 2678 3108 2730
rect 3052 2676 3108 2678
rect 3184 2730 3240 2732
rect 3184 2678 3186 2730
rect 3186 2678 3238 2730
rect 3238 2678 3240 2730
rect 3184 2676 3240 2678
rect 3316 2730 3372 2732
rect 3316 2678 3318 2730
rect 3318 2678 3370 2730
rect 3370 2678 3372 2730
rect 3316 2676 3372 2678
rect 3448 2730 3504 2732
rect 3448 2678 3450 2730
rect 3450 2678 3502 2730
rect 3502 2678 3504 2730
rect 3448 2676 3504 2678
rect 3580 2730 3636 2732
rect 3580 2678 3582 2730
rect 3582 2678 3634 2730
rect 3634 2678 3636 2730
rect 3580 2676 3636 2678
rect 3712 2730 3768 2732
rect 3712 2678 3714 2730
rect 3714 2678 3766 2730
rect 3766 2678 3768 2730
rect 3712 2676 3768 2678
rect 3844 2730 3900 2732
rect 3844 2678 3846 2730
rect 3846 2678 3898 2730
rect 3898 2678 3900 2730
rect 3844 2676 3900 2678
rect 3976 2730 4032 2732
rect 3976 2678 3978 2730
rect 3978 2678 4030 2730
rect 4030 2678 4032 2730
rect 3976 2676 4032 2678
rect 4108 2730 4164 2732
rect 4108 2678 4110 2730
rect 4110 2678 4162 2730
rect 4162 2678 4164 2730
rect 4108 2676 4164 2678
rect 4240 2730 4296 2732
rect 4240 2678 4242 2730
rect 4242 2678 4294 2730
rect 4294 2678 4296 2730
rect 4240 2676 4296 2678
rect 4372 2730 4428 2732
rect 4372 2678 4374 2730
rect 4374 2678 4426 2730
rect 4426 2678 4428 2730
rect 4372 2676 4428 2678
rect 4504 2730 4560 2732
rect 4504 2678 4506 2730
rect 4506 2678 4558 2730
rect 4558 2678 4560 2730
rect 4504 2676 4560 2678
rect 4636 2730 4692 2732
rect 4636 2678 4638 2730
rect 4638 2678 4690 2730
rect 4690 2678 4692 2730
rect 4636 2676 4692 2678
rect 4768 2730 4824 2732
rect 4768 2678 4770 2730
rect 4770 2678 4822 2730
rect 4822 2678 4824 2730
rect 4768 2676 4824 2678
rect 4900 2730 4956 2732
rect 4900 2678 4902 2730
rect 4902 2678 4954 2730
rect 4954 2678 4956 2730
rect 4900 2676 4956 2678
rect 5032 2730 5088 2732
rect 5032 2678 5034 2730
rect 5034 2678 5086 2730
rect 5086 2678 5088 2730
rect 5032 2676 5088 2678
rect 5164 2730 5220 2732
rect 5164 2678 5166 2730
rect 5166 2678 5218 2730
rect 5218 2678 5220 2730
rect 5164 2676 5220 2678
rect 5296 2730 5352 2732
rect 5296 2678 5298 2730
rect 5298 2678 5350 2730
rect 5350 2678 5352 2730
rect 5296 2676 5352 2678
rect 5428 2730 5484 2732
rect 5428 2678 5430 2730
rect 5430 2678 5482 2730
rect 5482 2678 5484 2730
rect 5428 2676 5484 2678
rect 5560 2730 5616 2732
rect 5560 2678 5562 2730
rect 5562 2678 5614 2730
rect 5614 2678 5616 2730
rect 5560 2676 5616 2678
rect 5692 2730 5748 2732
rect 5692 2678 5694 2730
rect 5694 2678 5746 2730
rect 5746 2678 5748 2730
rect 5692 2676 5748 2678
rect 5824 2730 5880 2732
rect 5824 2678 5826 2730
rect 5826 2678 5878 2730
rect 5878 2678 5880 2730
rect 5824 2676 5880 2678
rect 5956 2730 6012 2732
rect 5956 2678 5958 2730
rect 5958 2678 6010 2730
rect 6010 2678 6012 2730
rect 5956 2676 6012 2678
rect 6088 2730 6144 2732
rect 6088 2678 6090 2730
rect 6090 2678 6142 2730
rect 6142 2678 6144 2730
rect 6088 2676 6144 2678
rect 6220 2730 6276 2732
rect 6220 2678 6222 2730
rect 6222 2678 6274 2730
rect 6274 2678 6276 2730
rect 6220 2676 6276 2678
rect 6352 2730 6408 2732
rect 6352 2678 6354 2730
rect 6354 2678 6406 2730
rect 6406 2678 6408 2730
rect 6352 2676 6408 2678
rect 6484 2730 6540 2732
rect 6484 2678 6486 2730
rect 6486 2678 6538 2730
rect 6538 2678 6540 2730
rect 6484 2676 6540 2678
rect 6616 2730 6672 2732
rect 6616 2678 6618 2730
rect 6618 2678 6670 2730
rect 6670 2678 6672 2730
rect 6616 2676 6672 2678
rect 6748 2730 6804 2732
rect 6748 2678 6750 2730
rect 6750 2678 6802 2730
rect 6802 2678 6804 2730
rect 6748 2676 6804 2678
rect 6880 2730 6936 2732
rect 6880 2678 6882 2730
rect 6882 2678 6934 2730
rect 6934 2678 6936 2730
rect 6880 2676 6936 2678
rect 7012 2730 7068 2732
rect 7012 2678 7014 2730
rect 7014 2678 7066 2730
rect 7066 2678 7068 2730
rect 7012 2676 7068 2678
rect 7144 2730 7200 2732
rect 7144 2678 7146 2730
rect 7146 2678 7198 2730
rect 7198 2678 7200 2730
rect 7144 2676 7200 2678
rect 7276 2730 7332 2732
rect 7276 2678 7278 2730
rect 7278 2678 7330 2730
rect 7330 2678 7332 2730
rect 7276 2676 7332 2678
rect 7408 2730 7464 2732
rect 7408 2678 7410 2730
rect 7410 2678 7462 2730
rect 7462 2678 7464 2730
rect 7408 2676 7464 2678
rect 7540 2730 7596 2732
rect 7540 2678 7542 2730
rect 7542 2678 7594 2730
rect 7594 2678 7596 2730
rect 7540 2676 7596 2678
rect 8034 3063 8090 3065
rect 8034 2699 8036 3063
rect 8036 2699 8088 3063
rect 8088 2699 8090 3063
rect 8034 2697 8090 2699
rect 8482 3063 8538 3065
rect 8482 2699 8484 3063
rect 8484 2699 8536 3063
rect 8536 2699 8538 3063
rect 8482 2697 8538 2699
rect 2524 2598 2580 2600
rect 2524 2546 2526 2598
rect 2526 2546 2578 2598
rect 2578 2546 2580 2598
rect 2524 2544 2580 2546
rect 2656 2598 2712 2600
rect 2656 2546 2658 2598
rect 2658 2546 2710 2598
rect 2710 2546 2712 2598
rect 2656 2544 2712 2546
rect 2788 2598 2844 2600
rect 2788 2546 2790 2598
rect 2790 2546 2842 2598
rect 2842 2546 2844 2598
rect 2788 2544 2844 2546
rect 2920 2598 2976 2600
rect 2920 2546 2922 2598
rect 2922 2546 2974 2598
rect 2974 2546 2976 2598
rect 2920 2544 2976 2546
rect 3052 2598 3108 2600
rect 3052 2546 3054 2598
rect 3054 2546 3106 2598
rect 3106 2546 3108 2598
rect 3052 2544 3108 2546
rect 3184 2598 3240 2600
rect 3184 2546 3186 2598
rect 3186 2546 3238 2598
rect 3238 2546 3240 2598
rect 3184 2544 3240 2546
rect 3316 2598 3372 2600
rect 3316 2546 3318 2598
rect 3318 2546 3370 2598
rect 3370 2546 3372 2598
rect 3316 2544 3372 2546
rect 3448 2598 3504 2600
rect 3448 2546 3450 2598
rect 3450 2546 3502 2598
rect 3502 2546 3504 2598
rect 3448 2544 3504 2546
rect 3580 2598 3636 2600
rect 3580 2546 3582 2598
rect 3582 2546 3634 2598
rect 3634 2546 3636 2598
rect 3580 2544 3636 2546
rect 3712 2598 3768 2600
rect 3712 2546 3714 2598
rect 3714 2546 3766 2598
rect 3766 2546 3768 2598
rect 3712 2544 3768 2546
rect 3844 2598 3900 2600
rect 3844 2546 3846 2598
rect 3846 2546 3898 2598
rect 3898 2546 3900 2598
rect 3844 2544 3900 2546
rect 3976 2598 4032 2600
rect 3976 2546 3978 2598
rect 3978 2546 4030 2598
rect 4030 2546 4032 2598
rect 3976 2544 4032 2546
rect 4108 2598 4164 2600
rect 4108 2546 4110 2598
rect 4110 2546 4162 2598
rect 4162 2546 4164 2598
rect 4108 2544 4164 2546
rect 4240 2598 4296 2600
rect 4240 2546 4242 2598
rect 4242 2546 4294 2598
rect 4294 2546 4296 2598
rect 4240 2544 4296 2546
rect 4372 2598 4428 2600
rect 4372 2546 4374 2598
rect 4374 2546 4426 2598
rect 4426 2546 4428 2598
rect 4372 2544 4428 2546
rect 4504 2598 4560 2600
rect 4504 2546 4506 2598
rect 4506 2546 4558 2598
rect 4558 2546 4560 2598
rect 4504 2544 4560 2546
rect 4636 2598 4692 2600
rect 4636 2546 4638 2598
rect 4638 2546 4690 2598
rect 4690 2546 4692 2598
rect 4636 2544 4692 2546
rect 4768 2598 4824 2600
rect 4768 2546 4770 2598
rect 4770 2546 4822 2598
rect 4822 2546 4824 2598
rect 4768 2544 4824 2546
rect 4900 2598 4956 2600
rect 4900 2546 4902 2598
rect 4902 2546 4954 2598
rect 4954 2546 4956 2598
rect 4900 2544 4956 2546
rect 5032 2598 5088 2600
rect 5032 2546 5034 2598
rect 5034 2546 5086 2598
rect 5086 2546 5088 2598
rect 5032 2544 5088 2546
rect 5164 2598 5220 2600
rect 5164 2546 5166 2598
rect 5166 2546 5218 2598
rect 5218 2546 5220 2598
rect 5164 2544 5220 2546
rect 5296 2598 5352 2600
rect 5296 2546 5298 2598
rect 5298 2546 5350 2598
rect 5350 2546 5352 2598
rect 5296 2544 5352 2546
rect 5428 2598 5484 2600
rect 5428 2546 5430 2598
rect 5430 2546 5482 2598
rect 5482 2546 5484 2598
rect 5428 2544 5484 2546
rect 5560 2598 5616 2600
rect 5560 2546 5562 2598
rect 5562 2546 5614 2598
rect 5614 2546 5616 2598
rect 5560 2544 5616 2546
rect 5692 2598 5748 2600
rect 5692 2546 5694 2598
rect 5694 2546 5746 2598
rect 5746 2546 5748 2598
rect 5692 2544 5748 2546
rect 5824 2598 5880 2600
rect 5824 2546 5826 2598
rect 5826 2546 5878 2598
rect 5878 2546 5880 2598
rect 5824 2544 5880 2546
rect 5956 2598 6012 2600
rect 5956 2546 5958 2598
rect 5958 2546 6010 2598
rect 6010 2546 6012 2598
rect 5956 2544 6012 2546
rect 6088 2598 6144 2600
rect 6088 2546 6090 2598
rect 6090 2546 6142 2598
rect 6142 2546 6144 2598
rect 6088 2544 6144 2546
rect 6220 2598 6276 2600
rect 6220 2546 6222 2598
rect 6222 2546 6274 2598
rect 6274 2546 6276 2598
rect 6220 2544 6276 2546
rect 6352 2598 6408 2600
rect 6352 2546 6354 2598
rect 6354 2546 6406 2598
rect 6406 2546 6408 2598
rect 6352 2544 6408 2546
rect 6484 2598 6540 2600
rect 6484 2546 6486 2598
rect 6486 2546 6538 2598
rect 6538 2546 6540 2598
rect 6484 2544 6540 2546
rect 6616 2598 6672 2600
rect 6616 2546 6618 2598
rect 6618 2546 6670 2598
rect 6670 2546 6672 2598
rect 6616 2544 6672 2546
rect 6748 2598 6804 2600
rect 6748 2546 6750 2598
rect 6750 2546 6802 2598
rect 6802 2546 6804 2598
rect 6748 2544 6804 2546
rect 6880 2598 6936 2600
rect 6880 2546 6882 2598
rect 6882 2546 6934 2598
rect 6934 2546 6936 2598
rect 6880 2544 6936 2546
rect 7012 2598 7068 2600
rect 7012 2546 7014 2598
rect 7014 2546 7066 2598
rect 7066 2546 7068 2598
rect 7012 2544 7068 2546
rect 7144 2598 7200 2600
rect 7144 2546 7146 2598
rect 7146 2546 7198 2598
rect 7198 2546 7200 2598
rect 7144 2544 7200 2546
rect 7276 2598 7332 2600
rect 7276 2546 7278 2598
rect 7278 2546 7330 2598
rect 7330 2546 7332 2598
rect 7276 2544 7332 2546
rect 7408 2598 7464 2600
rect 7408 2546 7410 2598
rect 7410 2546 7462 2598
rect 7462 2546 7464 2598
rect 7408 2544 7464 2546
rect 7540 2598 7596 2600
rect 7540 2546 7542 2598
rect 7542 2546 7594 2598
rect 7594 2546 7596 2598
rect 7540 2544 7596 2546
rect 2524 2466 2580 2468
rect 2524 2414 2526 2466
rect 2526 2414 2578 2466
rect 2578 2414 2580 2466
rect 2524 2412 2580 2414
rect 2656 2466 2712 2468
rect 2656 2414 2658 2466
rect 2658 2414 2710 2466
rect 2710 2414 2712 2466
rect 2656 2412 2712 2414
rect 2788 2466 2844 2468
rect 2788 2414 2790 2466
rect 2790 2414 2842 2466
rect 2842 2414 2844 2466
rect 2788 2412 2844 2414
rect 2920 2466 2976 2468
rect 2920 2414 2922 2466
rect 2922 2414 2974 2466
rect 2974 2414 2976 2466
rect 2920 2412 2976 2414
rect 3052 2466 3108 2468
rect 3052 2414 3054 2466
rect 3054 2414 3106 2466
rect 3106 2414 3108 2466
rect 3052 2412 3108 2414
rect 3184 2466 3240 2468
rect 3184 2414 3186 2466
rect 3186 2414 3238 2466
rect 3238 2414 3240 2466
rect 3184 2412 3240 2414
rect 3316 2466 3372 2468
rect 3316 2414 3318 2466
rect 3318 2414 3370 2466
rect 3370 2414 3372 2466
rect 3316 2412 3372 2414
rect 3448 2466 3504 2468
rect 3448 2414 3450 2466
rect 3450 2414 3502 2466
rect 3502 2414 3504 2466
rect 3448 2412 3504 2414
rect 3580 2466 3636 2468
rect 3580 2414 3582 2466
rect 3582 2414 3634 2466
rect 3634 2414 3636 2466
rect 3580 2412 3636 2414
rect 3712 2466 3768 2468
rect 3712 2414 3714 2466
rect 3714 2414 3766 2466
rect 3766 2414 3768 2466
rect 3712 2412 3768 2414
rect 3844 2466 3900 2468
rect 3844 2414 3846 2466
rect 3846 2414 3898 2466
rect 3898 2414 3900 2466
rect 3844 2412 3900 2414
rect 3976 2466 4032 2468
rect 3976 2414 3978 2466
rect 3978 2414 4030 2466
rect 4030 2414 4032 2466
rect 3976 2412 4032 2414
rect 4108 2466 4164 2468
rect 4108 2414 4110 2466
rect 4110 2414 4162 2466
rect 4162 2414 4164 2466
rect 4108 2412 4164 2414
rect 4240 2466 4296 2468
rect 4240 2414 4242 2466
rect 4242 2414 4294 2466
rect 4294 2414 4296 2466
rect 4240 2412 4296 2414
rect 4372 2466 4428 2468
rect 4372 2414 4374 2466
rect 4374 2414 4426 2466
rect 4426 2414 4428 2466
rect 4372 2412 4428 2414
rect 4504 2466 4560 2468
rect 4504 2414 4506 2466
rect 4506 2414 4558 2466
rect 4558 2414 4560 2466
rect 4504 2412 4560 2414
rect 4636 2466 4692 2468
rect 4636 2414 4638 2466
rect 4638 2414 4690 2466
rect 4690 2414 4692 2466
rect 4636 2412 4692 2414
rect 4768 2466 4824 2468
rect 4768 2414 4770 2466
rect 4770 2414 4822 2466
rect 4822 2414 4824 2466
rect 4768 2412 4824 2414
rect 4900 2466 4956 2468
rect 4900 2414 4902 2466
rect 4902 2414 4954 2466
rect 4954 2414 4956 2466
rect 4900 2412 4956 2414
rect 5032 2466 5088 2468
rect 5032 2414 5034 2466
rect 5034 2414 5086 2466
rect 5086 2414 5088 2466
rect 5032 2412 5088 2414
rect 5164 2466 5220 2468
rect 5164 2414 5166 2466
rect 5166 2414 5218 2466
rect 5218 2414 5220 2466
rect 5164 2412 5220 2414
rect 5296 2466 5352 2468
rect 5296 2414 5298 2466
rect 5298 2414 5350 2466
rect 5350 2414 5352 2466
rect 5296 2412 5352 2414
rect 5428 2466 5484 2468
rect 5428 2414 5430 2466
rect 5430 2414 5482 2466
rect 5482 2414 5484 2466
rect 5428 2412 5484 2414
rect 5560 2466 5616 2468
rect 5560 2414 5562 2466
rect 5562 2414 5614 2466
rect 5614 2414 5616 2466
rect 5560 2412 5616 2414
rect 5692 2466 5748 2468
rect 5692 2414 5694 2466
rect 5694 2414 5746 2466
rect 5746 2414 5748 2466
rect 5692 2412 5748 2414
rect 5824 2466 5880 2468
rect 5824 2414 5826 2466
rect 5826 2414 5878 2466
rect 5878 2414 5880 2466
rect 5824 2412 5880 2414
rect 5956 2466 6012 2468
rect 5956 2414 5958 2466
rect 5958 2414 6010 2466
rect 6010 2414 6012 2466
rect 5956 2412 6012 2414
rect 6088 2466 6144 2468
rect 6088 2414 6090 2466
rect 6090 2414 6142 2466
rect 6142 2414 6144 2466
rect 6088 2412 6144 2414
rect 6220 2466 6276 2468
rect 6220 2414 6222 2466
rect 6222 2414 6274 2466
rect 6274 2414 6276 2466
rect 6220 2412 6276 2414
rect 6352 2466 6408 2468
rect 6352 2414 6354 2466
rect 6354 2414 6406 2466
rect 6406 2414 6408 2466
rect 6352 2412 6408 2414
rect 6484 2466 6540 2468
rect 6484 2414 6486 2466
rect 6486 2414 6538 2466
rect 6538 2414 6540 2466
rect 6484 2412 6540 2414
rect 6616 2466 6672 2468
rect 6616 2414 6618 2466
rect 6618 2414 6670 2466
rect 6670 2414 6672 2466
rect 6616 2412 6672 2414
rect 6748 2466 6804 2468
rect 6748 2414 6750 2466
rect 6750 2414 6802 2466
rect 6802 2414 6804 2466
rect 6748 2412 6804 2414
rect 6880 2466 6936 2468
rect 6880 2414 6882 2466
rect 6882 2414 6934 2466
rect 6934 2414 6936 2466
rect 6880 2412 6936 2414
rect 7012 2466 7068 2468
rect 7012 2414 7014 2466
rect 7014 2414 7066 2466
rect 7066 2414 7068 2466
rect 7012 2412 7068 2414
rect 7144 2466 7200 2468
rect 7144 2414 7146 2466
rect 7146 2414 7198 2466
rect 7198 2414 7200 2466
rect 7144 2412 7200 2414
rect 7276 2466 7332 2468
rect 7276 2414 7278 2466
rect 7278 2414 7330 2466
rect 7330 2414 7332 2466
rect 7276 2412 7332 2414
rect 7408 2466 7464 2468
rect 7408 2414 7410 2466
rect 7410 2414 7462 2466
rect 7462 2414 7464 2466
rect 7408 2412 7464 2414
rect 7540 2466 7596 2468
rect 7540 2414 7542 2466
rect 7542 2414 7594 2466
rect 7594 2414 7596 2466
rect 7540 2412 7596 2414
rect 2524 2334 2580 2336
rect 2524 2282 2526 2334
rect 2526 2282 2578 2334
rect 2578 2282 2580 2334
rect 2524 2280 2580 2282
rect 2656 2334 2712 2336
rect 2656 2282 2658 2334
rect 2658 2282 2710 2334
rect 2710 2282 2712 2334
rect 2656 2280 2712 2282
rect 2788 2334 2844 2336
rect 2788 2282 2790 2334
rect 2790 2282 2842 2334
rect 2842 2282 2844 2334
rect 2788 2280 2844 2282
rect 2920 2334 2976 2336
rect 2920 2282 2922 2334
rect 2922 2282 2974 2334
rect 2974 2282 2976 2334
rect 2920 2280 2976 2282
rect 3052 2334 3108 2336
rect 3052 2282 3054 2334
rect 3054 2282 3106 2334
rect 3106 2282 3108 2334
rect 3052 2280 3108 2282
rect 3184 2334 3240 2336
rect 3184 2282 3186 2334
rect 3186 2282 3238 2334
rect 3238 2282 3240 2334
rect 3184 2280 3240 2282
rect 3316 2334 3372 2336
rect 3316 2282 3318 2334
rect 3318 2282 3370 2334
rect 3370 2282 3372 2334
rect 3316 2280 3372 2282
rect 3448 2334 3504 2336
rect 3448 2282 3450 2334
rect 3450 2282 3502 2334
rect 3502 2282 3504 2334
rect 3448 2280 3504 2282
rect 3580 2334 3636 2336
rect 3580 2282 3582 2334
rect 3582 2282 3634 2334
rect 3634 2282 3636 2334
rect 3580 2280 3636 2282
rect 3712 2334 3768 2336
rect 3712 2282 3714 2334
rect 3714 2282 3766 2334
rect 3766 2282 3768 2334
rect 3712 2280 3768 2282
rect 3844 2334 3900 2336
rect 3844 2282 3846 2334
rect 3846 2282 3898 2334
rect 3898 2282 3900 2334
rect 3844 2280 3900 2282
rect 3976 2334 4032 2336
rect 3976 2282 3978 2334
rect 3978 2282 4030 2334
rect 4030 2282 4032 2334
rect 3976 2280 4032 2282
rect 4108 2334 4164 2336
rect 4108 2282 4110 2334
rect 4110 2282 4162 2334
rect 4162 2282 4164 2334
rect 4108 2280 4164 2282
rect 4240 2334 4296 2336
rect 4240 2282 4242 2334
rect 4242 2282 4294 2334
rect 4294 2282 4296 2334
rect 4240 2280 4296 2282
rect 4372 2334 4428 2336
rect 4372 2282 4374 2334
rect 4374 2282 4426 2334
rect 4426 2282 4428 2334
rect 4372 2280 4428 2282
rect 4504 2334 4560 2336
rect 4504 2282 4506 2334
rect 4506 2282 4558 2334
rect 4558 2282 4560 2334
rect 4504 2280 4560 2282
rect 4636 2334 4692 2336
rect 4636 2282 4638 2334
rect 4638 2282 4690 2334
rect 4690 2282 4692 2334
rect 4636 2280 4692 2282
rect 4768 2334 4824 2336
rect 4768 2282 4770 2334
rect 4770 2282 4822 2334
rect 4822 2282 4824 2334
rect 4768 2280 4824 2282
rect 4900 2334 4956 2336
rect 4900 2282 4902 2334
rect 4902 2282 4954 2334
rect 4954 2282 4956 2334
rect 4900 2280 4956 2282
rect 5032 2334 5088 2336
rect 5032 2282 5034 2334
rect 5034 2282 5086 2334
rect 5086 2282 5088 2334
rect 5032 2280 5088 2282
rect 5164 2334 5220 2336
rect 5164 2282 5166 2334
rect 5166 2282 5218 2334
rect 5218 2282 5220 2334
rect 5164 2280 5220 2282
rect 5296 2334 5352 2336
rect 5296 2282 5298 2334
rect 5298 2282 5350 2334
rect 5350 2282 5352 2334
rect 5296 2280 5352 2282
rect 5428 2334 5484 2336
rect 5428 2282 5430 2334
rect 5430 2282 5482 2334
rect 5482 2282 5484 2334
rect 5428 2280 5484 2282
rect 5560 2334 5616 2336
rect 5560 2282 5562 2334
rect 5562 2282 5614 2334
rect 5614 2282 5616 2334
rect 5560 2280 5616 2282
rect 5692 2334 5748 2336
rect 5692 2282 5694 2334
rect 5694 2282 5746 2334
rect 5746 2282 5748 2334
rect 5692 2280 5748 2282
rect 5824 2334 5880 2336
rect 5824 2282 5826 2334
rect 5826 2282 5878 2334
rect 5878 2282 5880 2334
rect 5824 2280 5880 2282
rect 5956 2334 6012 2336
rect 5956 2282 5958 2334
rect 5958 2282 6010 2334
rect 6010 2282 6012 2334
rect 5956 2280 6012 2282
rect 6088 2334 6144 2336
rect 6088 2282 6090 2334
rect 6090 2282 6142 2334
rect 6142 2282 6144 2334
rect 6088 2280 6144 2282
rect 6220 2334 6276 2336
rect 6220 2282 6222 2334
rect 6222 2282 6274 2334
rect 6274 2282 6276 2334
rect 6220 2280 6276 2282
rect 6352 2334 6408 2336
rect 6352 2282 6354 2334
rect 6354 2282 6406 2334
rect 6406 2282 6408 2334
rect 6352 2280 6408 2282
rect 6484 2334 6540 2336
rect 6484 2282 6486 2334
rect 6486 2282 6538 2334
rect 6538 2282 6540 2334
rect 6484 2280 6540 2282
rect 6616 2334 6672 2336
rect 6616 2282 6618 2334
rect 6618 2282 6670 2334
rect 6670 2282 6672 2334
rect 6616 2280 6672 2282
rect 6748 2334 6804 2336
rect 6748 2282 6750 2334
rect 6750 2282 6802 2334
rect 6802 2282 6804 2334
rect 6748 2280 6804 2282
rect 6880 2334 6936 2336
rect 6880 2282 6882 2334
rect 6882 2282 6934 2334
rect 6934 2282 6936 2334
rect 6880 2280 6936 2282
rect 7012 2334 7068 2336
rect 7012 2282 7014 2334
rect 7014 2282 7066 2334
rect 7066 2282 7068 2334
rect 7012 2280 7068 2282
rect 7144 2334 7200 2336
rect 7144 2282 7146 2334
rect 7146 2282 7198 2334
rect 7198 2282 7200 2334
rect 7144 2280 7200 2282
rect 7276 2334 7332 2336
rect 7276 2282 7278 2334
rect 7278 2282 7330 2334
rect 7330 2282 7332 2334
rect 7276 2280 7332 2282
rect 7408 2334 7464 2336
rect 7408 2282 7410 2334
rect 7410 2282 7462 2334
rect 7462 2282 7464 2334
rect 7408 2280 7464 2282
rect 7540 2334 7596 2336
rect 7540 2282 7542 2334
rect 7542 2282 7594 2334
rect 7594 2282 7596 2334
rect 7540 2280 7596 2282
rect 8979 4701 9035 4703
rect 8979 4649 8981 4701
rect 8981 4649 9033 4701
rect 9033 4649 9035 4701
rect 8979 4647 9035 4649
rect 9191 4701 9247 4703
rect 9191 4649 9193 4701
rect 9193 4649 9245 4701
rect 9245 4649 9247 4701
rect 9191 4647 9247 4649
rect 8979 4483 9035 4485
rect 8979 4431 8981 4483
rect 8981 4431 9033 4483
rect 9033 4431 9035 4483
rect 8979 4429 9035 4431
rect 9191 4483 9247 4485
rect 9191 4431 9193 4483
rect 9193 4431 9245 4483
rect 9245 4431 9247 4483
rect 9191 4429 9247 4431
rect 8979 4265 9035 4267
rect 8979 4213 8981 4265
rect 8981 4213 9033 4265
rect 9033 4213 9035 4265
rect 8979 4211 9035 4213
rect 9191 4265 9247 4267
rect 9191 4213 9193 4265
rect 9193 4213 9245 4265
rect 9245 4213 9247 4265
rect 9191 4211 9247 4213
rect 8979 4047 9035 4049
rect 8979 3995 8981 4047
rect 8981 3995 9033 4047
rect 9033 3995 9035 4047
rect 8979 3993 9035 3995
rect 9191 4047 9247 4049
rect 9191 3995 9193 4047
rect 9193 3995 9245 4047
rect 9245 3995 9247 4047
rect 9191 3993 9247 3995
rect 9452 4734 9508 4736
rect 9452 4682 9454 4734
rect 9454 4682 9506 4734
rect 9506 4682 9508 4734
rect 9452 4680 9508 4682
rect 9452 4517 9508 4519
rect 9452 4465 9454 4517
rect 9454 4465 9506 4517
rect 9506 4465 9508 4517
rect 9452 4463 9508 4465
rect 9452 4299 9508 4301
rect 9452 4247 9454 4299
rect 9454 4247 9506 4299
rect 9506 4247 9508 4299
rect 9452 4245 9508 4247
rect 9452 4081 9508 4083
rect 9452 4029 9454 4081
rect 9454 4029 9506 4081
rect 9506 4029 9508 4081
rect 9452 4027 9508 4029
rect 9452 3864 9508 3866
rect 9452 3812 9454 3864
rect 9454 3812 9506 3864
rect 9506 3812 9508 3864
rect 9452 3810 9508 3812
rect 9452 3646 9508 3648
rect 9452 3594 9454 3646
rect 9454 3594 9506 3646
rect 9506 3594 9508 3646
rect 9452 3592 9508 3594
rect 9452 3429 9508 3431
rect 9452 3377 9454 3429
rect 9454 3377 9506 3429
rect 9506 3377 9508 3429
rect 9452 3375 9508 3377
rect 9452 3211 9508 3213
rect 9452 3159 9454 3211
rect 9454 3159 9506 3211
rect 9506 3159 9508 3211
rect 9452 3157 9508 3159
rect 9452 2993 9508 2995
rect 9452 2941 9454 2993
rect 9454 2941 9506 2993
rect 9506 2941 9508 2993
rect 9452 2939 9508 2941
rect 9452 2776 9508 2778
rect 9452 2724 9454 2776
rect 9454 2724 9506 2776
rect 9506 2724 9508 2776
rect 9452 2722 9508 2724
rect 9452 2558 9508 2560
rect 9452 2506 9454 2558
rect 9454 2506 9506 2558
rect 9506 2506 9508 2558
rect 9452 2504 9508 2506
rect 9452 2340 9508 2342
rect 9452 2288 9454 2340
rect 9454 2288 9506 2340
rect 9506 2288 9508 2340
rect 9452 2286 9508 2288
rect 9452 2123 9508 2125
rect 9452 2071 9454 2123
rect 9454 2071 9506 2123
rect 9506 2071 9508 2123
rect 9452 2069 9508 2071
rect 9452 1905 9508 1907
rect 9452 1853 9454 1905
rect 9454 1853 9506 1905
rect 9506 1853 9508 1905
rect 9452 1851 9508 1853
rect 9452 1687 9508 1689
rect 9452 1635 9454 1687
rect 9454 1635 9506 1687
rect 9506 1635 9508 1687
rect 9452 1633 9508 1635
rect 9452 1470 9508 1472
rect 9452 1418 9454 1470
rect 9454 1418 9506 1470
rect 9506 1418 9508 1470
rect 9452 1416 9508 1418
rect 9452 1252 9508 1254
rect 9452 1200 9454 1252
rect 9454 1200 9506 1252
rect 9506 1200 9508 1252
rect 9452 1198 9508 1200
rect 9452 1035 9508 1037
rect 9452 983 9454 1035
rect 9454 983 9506 1035
rect 9506 983 9508 1035
rect 9452 981 9508 983
rect 9452 817 9508 819
rect 9452 765 9454 817
rect 9454 765 9506 817
rect 9506 765 9508 817
rect 9452 763 9508 765
rect 9452 599 9508 601
rect 9452 547 9454 599
rect 9454 547 9506 599
rect 9506 547 9508 599
rect 9452 545 9508 547
rect 9452 382 9508 384
rect 9452 330 9454 382
rect 9454 330 9506 382
rect 9506 330 9508 382
rect 9452 328 9508 330
rect 11847 9274 11903 9330
rect 12058 9274 12114 9330
rect 12269 9274 12325 9330
rect 12480 9274 12536 9330
rect 12691 9274 12747 9330
rect 12902 9274 12958 9330
rect 13113 9274 13169 9330
rect 10642 9163 10698 9219
rect 11093 9163 11149 9219
rect 11541 9163 11597 9219
rect 10642 8945 10698 9001
rect 11093 8945 11149 9001
rect 10869 8386 10925 8388
rect 10869 8334 10871 8386
rect 10871 8334 10923 8386
rect 10923 8334 10925 8386
rect 10869 8332 10925 8334
rect 10869 8169 10925 8171
rect 10869 8117 10871 8169
rect 10871 8117 10923 8169
rect 10923 8117 10925 8169
rect 10869 8115 10925 8117
rect 10869 7951 10925 7953
rect 10869 7899 10871 7951
rect 10871 7899 10923 7951
rect 10923 7899 10925 7951
rect 10869 7897 10925 7899
rect 10869 7734 10925 7736
rect 10869 7682 10871 7734
rect 10871 7682 10923 7734
rect 10923 7682 10925 7734
rect 10869 7680 10925 7682
rect 10869 7516 10925 7518
rect 10869 7464 10871 7516
rect 10871 7464 10923 7516
rect 10923 7464 10925 7516
rect 10869 7462 10925 7464
rect 10869 7298 10925 7300
rect 10869 7246 10871 7298
rect 10871 7246 10923 7298
rect 10923 7246 10925 7298
rect 10869 7244 10925 7246
rect 10869 7080 10925 7082
rect 10869 7028 10871 7080
rect 10871 7028 10923 7080
rect 10923 7028 10925 7080
rect 10869 7026 10925 7028
rect 10869 6863 10925 6865
rect 10869 6811 10871 6863
rect 10871 6811 10923 6863
rect 10923 6811 10925 6863
rect 10869 6809 10925 6811
rect 10869 6645 10925 6647
rect 10869 6593 10871 6645
rect 10871 6593 10923 6645
rect 10923 6593 10925 6645
rect 10869 6591 10925 6593
rect 10869 6428 10925 6430
rect 10869 6376 10871 6428
rect 10871 6376 10923 6428
rect 10923 6376 10925 6428
rect 10869 6374 10925 6376
rect 11541 8945 11597 9001
rect 11847 9056 11903 9112
rect 12058 9056 12114 9112
rect 12269 9056 12325 9112
rect 12480 9056 12536 9112
rect 12691 9056 12747 9112
rect 12902 9056 12958 9112
rect 13113 9056 13169 9112
rect 11847 8838 11903 8894
rect 12058 8838 12114 8894
rect 12269 8838 12325 8894
rect 12480 8838 12536 8894
rect 12691 8838 12747 8894
rect 12902 8838 12958 8894
rect 13113 8838 13169 8894
rect 11847 8620 11903 8676
rect 12058 8620 12114 8676
rect 12269 8620 12325 8676
rect 12480 8620 12536 8676
rect 12691 8620 12747 8676
rect 12902 8620 12958 8676
rect 13113 8620 13169 8676
rect 11317 8386 11373 8388
rect 11317 8334 11319 8386
rect 11319 8334 11371 8386
rect 11371 8334 11373 8386
rect 11317 8332 11373 8334
rect 11317 8169 11373 8171
rect 11317 8117 11319 8169
rect 11319 8117 11371 8169
rect 11371 8117 11373 8169
rect 11317 8115 11373 8117
rect 11317 7951 11373 7953
rect 11317 7899 11319 7951
rect 11319 7899 11371 7951
rect 11371 7899 11373 7951
rect 11317 7897 11373 7899
rect 11317 7734 11373 7736
rect 11317 7682 11319 7734
rect 11319 7682 11371 7734
rect 11371 7682 11373 7734
rect 11317 7680 11373 7682
rect 11317 7516 11373 7518
rect 11317 7464 11319 7516
rect 11319 7464 11371 7516
rect 11371 7464 11373 7516
rect 11317 7462 11373 7464
rect 11317 7298 11373 7300
rect 11317 7246 11319 7298
rect 11319 7246 11371 7298
rect 11371 7246 11373 7298
rect 11317 7244 11373 7246
rect 11317 7080 11373 7082
rect 11317 7028 11319 7080
rect 11319 7028 11371 7080
rect 11371 7028 11373 7080
rect 11317 7026 11373 7028
rect 11317 6863 11373 6865
rect 11317 6811 11319 6863
rect 11319 6811 11371 6863
rect 11371 6811 11373 6863
rect 11317 6809 11373 6811
rect 11317 6645 11373 6647
rect 11317 6593 11319 6645
rect 11319 6593 11371 6645
rect 11371 6593 11373 6645
rect 11317 6591 11373 6593
rect 11317 6428 11373 6430
rect 11317 6376 11319 6428
rect 11319 6376 11371 6428
rect 11371 6376 11373 6428
rect 11317 6374 11373 6376
rect 12151 8400 12207 8402
rect 12151 8348 12153 8400
rect 12153 8348 12205 8400
rect 12205 8348 12207 8400
rect 12151 8346 12207 8348
rect 12151 8183 12207 8185
rect 12151 8131 12153 8183
rect 12153 8131 12205 8183
rect 12205 8131 12207 8183
rect 12151 8129 12207 8131
rect 12151 7965 12207 7967
rect 12151 7913 12153 7965
rect 12153 7913 12205 7965
rect 12205 7913 12207 7965
rect 12151 7911 12207 7913
rect 12151 7748 12207 7750
rect 12151 7696 12153 7748
rect 12153 7696 12205 7748
rect 12205 7696 12207 7748
rect 12151 7694 12207 7696
rect 12151 7530 12207 7532
rect 12151 7478 12153 7530
rect 12153 7478 12205 7530
rect 12205 7478 12207 7530
rect 12151 7476 12207 7478
rect 12151 7312 12207 7314
rect 12151 7260 12153 7312
rect 12153 7260 12205 7312
rect 12205 7260 12207 7312
rect 12151 7258 12207 7260
rect 12151 7094 12207 7096
rect 12151 7042 12153 7094
rect 12153 7042 12205 7094
rect 12205 7042 12207 7094
rect 12151 7040 12207 7042
rect 12151 6877 12207 6879
rect 12151 6825 12153 6877
rect 12153 6825 12205 6877
rect 12205 6825 12207 6877
rect 12151 6823 12207 6825
rect 12151 6659 12207 6661
rect 12151 6607 12153 6659
rect 12153 6607 12205 6659
rect 12205 6607 12207 6659
rect 12151 6605 12207 6607
rect 12151 6442 12207 6444
rect 12151 6390 12153 6442
rect 12153 6390 12205 6442
rect 12205 6390 12207 6442
rect 12151 6388 12207 6390
rect 12599 8400 12655 8402
rect 12599 8348 12601 8400
rect 12601 8348 12653 8400
rect 12653 8348 12655 8400
rect 12599 8346 12655 8348
rect 12599 8183 12655 8185
rect 12599 8131 12601 8183
rect 12601 8131 12653 8183
rect 12653 8131 12655 8183
rect 12599 8129 12655 8131
rect 12599 7965 12655 7967
rect 12599 7913 12601 7965
rect 12601 7913 12653 7965
rect 12653 7913 12655 7965
rect 12599 7911 12655 7913
rect 12599 7748 12655 7750
rect 12599 7696 12601 7748
rect 12601 7696 12653 7748
rect 12653 7696 12655 7748
rect 12599 7694 12655 7696
rect 12599 7530 12655 7532
rect 12599 7478 12601 7530
rect 12601 7478 12653 7530
rect 12653 7478 12655 7530
rect 12599 7476 12655 7478
rect 12599 7312 12655 7314
rect 12599 7260 12601 7312
rect 12601 7260 12653 7312
rect 12653 7260 12655 7312
rect 12599 7258 12655 7260
rect 12599 7094 12655 7096
rect 12599 7042 12601 7094
rect 12601 7042 12653 7094
rect 12653 7042 12655 7094
rect 12599 7040 12655 7042
rect 12599 6877 12655 6879
rect 12599 6825 12601 6877
rect 12601 6825 12653 6877
rect 12653 6825 12655 6877
rect 12599 6823 12655 6825
rect 12599 6659 12655 6661
rect 12599 6607 12601 6659
rect 12601 6607 12653 6659
rect 12653 6607 12655 6659
rect 12599 6605 12655 6607
rect 12599 6442 12655 6444
rect 12599 6390 12601 6442
rect 12601 6390 12653 6442
rect 12653 6390 12655 6442
rect 12599 6388 12655 6390
rect 12631 4512 12687 4514
rect 12631 4460 12633 4512
rect 12633 4460 12685 4512
rect 12685 4460 12687 4512
rect 12631 4458 12687 4460
rect 12843 4512 12899 4514
rect 12843 4460 12845 4512
rect 12845 4460 12897 4512
rect 12897 4460 12899 4512
rect 12843 4458 12899 4460
rect 10645 3991 10701 3993
rect 10645 3939 10647 3991
rect 10647 3939 10699 3991
rect 10699 3939 10701 3991
rect 10645 3937 10701 3939
rect 10645 3773 10701 3775
rect 10645 3721 10647 3773
rect 10647 3721 10699 3773
rect 10699 3721 10701 3773
rect 10645 3719 10701 3721
rect 10645 3556 10701 3558
rect 10645 3504 10647 3556
rect 10647 3504 10699 3556
rect 10699 3504 10701 3556
rect 10645 3502 10701 3504
rect 10645 3338 10701 3340
rect 10645 3286 10647 3338
rect 10647 3286 10699 3338
rect 10699 3286 10701 3338
rect 10645 3284 10701 3286
rect 10645 3120 10701 3122
rect 10645 3068 10647 3120
rect 10647 3068 10699 3120
rect 10699 3068 10701 3120
rect 10645 3066 10701 3068
rect 10645 2903 10701 2905
rect 10645 2851 10647 2903
rect 10647 2851 10699 2903
rect 10699 2851 10701 2903
rect 10645 2849 10701 2851
rect 10645 2685 10701 2687
rect 10645 2633 10647 2685
rect 10647 2633 10699 2685
rect 10699 2633 10701 2685
rect 10645 2631 10701 2633
rect 10645 2468 10701 2470
rect 10645 2416 10647 2468
rect 10647 2416 10699 2468
rect 10699 2416 10701 2468
rect 10645 2414 10701 2416
rect 10645 2250 10701 2252
rect 10645 2198 10647 2250
rect 10647 2198 10699 2250
rect 10699 2198 10701 2250
rect 10645 2196 10701 2198
rect 11541 3991 11597 3993
rect 11541 3939 11543 3991
rect 11543 3939 11595 3991
rect 11595 3939 11597 3991
rect 11541 3937 11597 3939
rect 11541 3773 11597 3775
rect 11541 3721 11543 3773
rect 11543 3721 11595 3773
rect 11595 3721 11597 3773
rect 11541 3719 11597 3721
rect 11541 3556 11597 3558
rect 11541 3504 11543 3556
rect 11543 3504 11595 3556
rect 11595 3504 11597 3556
rect 11541 3502 11597 3504
rect 11541 3338 11597 3340
rect 11541 3286 11543 3338
rect 11543 3286 11595 3338
rect 11595 3286 11597 3338
rect 11541 3284 11597 3286
rect 11541 3120 11597 3122
rect 11541 3068 11543 3120
rect 11543 3068 11595 3120
rect 11595 3068 11597 3120
rect 11541 3066 11597 3068
rect 11541 2903 11597 2905
rect 11541 2851 11543 2903
rect 11543 2851 11595 2903
rect 11595 2851 11597 2903
rect 11541 2849 11597 2851
rect 11541 2685 11597 2687
rect 11541 2633 11543 2685
rect 11543 2633 11595 2685
rect 11595 2633 11597 2685
rect 11541 2631 11597 2633
rect 11541 2468 11597 2470
rect 11541 2416 11543 2468
rect 11543 2416 11595 2468
rect 11595 2416 11597 2468
rect 11541 2414 11597 2416
rect 10645 2032 10701 2034
rect 10645 1980 10647 2032
rect 10647 1980 10699 2032
rect 10699 1980 10701 2032
rect 10645 1978 10701 1980
rect 10645 1814 10701 1816
rect 10645 1762 10647 1814
rect 10647 1762 10699 1814
rect 10699 1762 10701 1814
rect 10645 1760 10701 1762
rect 10645 1597 10701 1599
rect 10645 1545 10647 1597
rect 10647 1545 10699 1597
rect 10699 1545 10701 1597
rect 10645 1543 10701 1545
rect 10645 1379 10701 1381
rect 10645 1327 10647 1379
rect 10647 1327 10699 1379
rect 10699 1327 10701 1379
rect 10645 1325 10701 1327
rect 10645 1162 10701 1164
rect 10645 1110 10647 1162
rect 10647 1110 10699 1162
rect 10699 1110 10701 1162
rect 10645 1108 10701 1110
rect 10645 944 10701 946
rect 10645 892 10647 944
rect 10647 892 10699 944
rect 10699 892 10701 944
rect 10645 890 10701 892
rect 10645 726 10701 728
rect 10645 674 10647 726
rect 10647 674 10699 726
rect 10699 674 10701 726
rect 10645 672 10701 674
rect 10645 509 10701 511
rect 10645 457 10647 509
rect 10647 457 10699 509
rect 10699 457 10701 509
rect 10645 455 10701 457
rect 10645 291 10701 293
rect 10645 239 10647 291
rect 10647 239 10699 291
rect 10699 239 10701 291
rect 10645 237 10701 239
rect 11541 2250 11597 2252
rect 11541 2198 11543 2250
rect 11543 2198 11595 2250
rect 11595 2198 11597 2250
rect 11541 2196 11597 2198
rect 11541 2032 11597 2034
rect 11541 1980 11543 2032
rect 11543 1980 11595 2032
rect 11595 1980 11597 2032
rect 11541 1978 11597 1980
rect 11541 1814 11597 1816
rect 11541 1762 11543 1814
rect 11543 1762 11595 1814
rect 11595 1762 11597 1814
rect 11541 1760 11597 1762
rect 11541 1597 11597 1599
rect 11541 1545 11543 1597
rect 11543 1545 11595 1597
rect 11595 1545 11597 1597
rect 11541 1543 11597 1545
rect 11541 1379 11597 1381
rect 11541 1327 11543 1379
rect 11543 1327 11595 1379
rect 11595 1327 11597 1379
rect 11541 1325 11597 1327
rect 11541 1162 11597 1164
rect 11541 1110 11543 1162
rect 11543 1110 11595 1162
rect 11595 1110 11597 1162
rect 11541 1108 11597 1110
rect 11541 944 11597 946
rect 11541 892 11543 944
rect 11543 892 11595 944
rect 11595 892 11597 944
rect 11541 890 11597 892
rect 11541 726 11597 728
rect 11541 674 11543 726
rect 11543 674 11595 726
rect 11595 674 11597 726
rect 11541 672 11597 674
rect 11541 509 11597 511
rect 11541 457 11543 509
rect 11543 457 11595 509
rect 11595 457 11597 509
rect 11541 455 11597 457
rect 11541 291 11597 293
rect 11541 239 11543 291
rect 11543 239 11595 291
rect 11595 239 11597 291
rect 11541 237 11597 239
rect 11929 3991 11985 3993
rect 11929 3939 11931 3991
rect 11931 3939 11983 3991
rect 11983 3939 11985 3991
rect 11929 3937 11985 3939
rect 11929 3773 11985 3775
rect 11929 3721 11931 3773
rect 11931 3721 11983 3773
rect 11983 3721 11985 3773
rect 11929 3719 11985 3721
rect 11929 3556 11985 3558
rect 11929 3504 11931 3556
rect 11931 3504 11983 3556
rect 11983 3504 11985 3556
rect 11929 3502 11985 3504
rect 11929 3338 11985 3340
rect 11929 3286 11931 3338
rect 11931 3286 11983 3338
rect 11983 3286 11985 3338
rect 11929 3284 11985 3286
rect 11929 3120 11985 3122
rect 11929 3068 11931 3120
rect 11931 3068 11983 3120
rect 11983 3068 11985 3120
rect 11929 3066 11985 3068
rect 11929 2903 11985 2905
rect 11929 2851 11931 2903
rect 11931 2851 11983 2903
rect 11983 2851 11985 2903
rect 11929 2849 11985 2851
rect 11929 2685 11985 2687
rect 11929 2633 11931 2685
rect 11931 2633 11983 2685
rect 11983 2633 11985 2685
rect 11929 2631 11985 2633
rect 11929 2468 11985 2470
rect 11929 2416 11931 2468
rect 11931 2416 11983 2468
rect 11983 2416 11985 2468
rect 11929 2414 11985 2416
rect 11929 2250 11985 2252
rect 11929 2198 11931 2250
rect 11931 2198 11983 2250
rect 11983 2198 11985 2250
rect 11929 2196 11985 2198
rect 12825 3991 12881 3993
rect 12825 3939 12827 3991
rect 12827 3939 12879 3991
rect 12879 3939 12881 3991
rect 12825 3937 12881 3939
rect 12825 3773 12881 3775
rect 12825 3721 12827 3773
rect 12827 3721 12879 3773
rect 12879 3721 12881 3773
rect 12825 3719 12881 3721
rect 12825 3556 12881 3558
rect 12825 3504 12827 3556
rect 12827 3504 12879 3556
rect 12879 3504 12881 3556
rect 12825 3502 12881 3504
rect 12825 3338 12881 3340
rect 12825 3286 12827 3338
rect 12827 3286 12879 3338
rect 12879 3286 12881 3338
rect 12825 3284 12881 3286
rect 12825 3120 12881 3122
rect 12825 3068 12827 3120
rect 12827 3068 12879 3120
rect 12879 3068 12881 3120
rect 12825 3066 12881 3068
rect 12825 2903 12881 2905
rect 12825 2851 12827 2903
rect 12827 2851 12879 2903
rect 12879 2851 12881 2903
rect 12825 2849 12881 2851
rect 12825 2685 12881 2687
rect 12825 2633 12827 2685
rect 12827 2633 12879 2685
rect 12879 2633 12881 2685
rect 12825 2631 12881 2633
rect 12825 2468 12881 2470
rect 12825 2416 12827 2468
rect 12827 2416 12879 2468
rect 12879 2416 12881 2468
rect 12825 2414 12881 2416
rect 11929 2032 11985 2034
rect 11929 1980 11931 2032
rect 11931 1980 11983 2032
rect 11983 1980 11985 2032
rect 11929 1978 11985 1980
rect 11929 1814 11985 1816
rect 11929 1762 11931 1814
rect 11931 1762 11983 1814
rect 11983 1762 11985 1814
rect 11929 1760 11985 1762
rect 11929 1597 11985 1599
rect 11929 1545 11931 1597
rect 11931 1545 11983 1597
rect 11983 1545 11985 1597
rect 11929 1543 11985 1545
rect 11929 1379 11985 1381
rect 11929 1327 11931 1379
rect 11931 1327 11983 1379
rect 11983 1327 11985 1379
rect 11929 1325 11985 1327
rect 11929 1162 11985 1164
rect 11929 1110 11931 1162
rect 11931 1110 11983 1162
rect 11983 1110 11985 1162
rect 11929 1108 11985 1110
rect 11929 944 11985 946
rect 11929 892 11931 944
rect 11931 892 11983 944
rect 11983 892 11985 944
rect 11929 890 11985 892
rect 11929 726 11985 728
rect 11929 674 11931 726
rect 11931 674 11983 726
rect 11983 674 11985 726
rect 11929 672 11985 674
rect 11929 509 11985 511
rect 11929 457 11931 509
rect 11931 457 11983 509
rect 11983 457 11985 509
rect 11929 455 11985 457
rect 11929 291 11985 293
rect 11929 239 11931 291
rect 11931 239 11983 291
rect 11983 239 11985 291
rect 11929 237 11985 239
rect 12825 2250 12881 2252
rect 12825 2198 12827 2250
rect 12827 2198 12879 2250
rect 12879 2198 12881 2250
rect 12825 2196 12881 2198
rect 12825 2032 12881 2034
rect 12825 1980 12827 2032
rect 12827 1980 12879 2032
rect 12879 1980 12881 2032
rect 12825 1978 12881 1980
rect 12825 1814 12881 1816
rect 12825 1762 12827 1814
rect 12827 1762 12879 1814
rect 12879 1762 12881 1814
rect 12825 1760 12881 1762
rect 12825 1597 12881 1599
rect 12825 1545 12827 1597
rect 12827 1545 12879 1597
rect 12879 1545 12881 1597
rect 12825 1543 12881 1545
rect 12825 1379 12881 1381
rect 12825 1327 12827 1379
rect 12827 1327 12879 1379
rect 12879 1327 12881 1379
rect 12825 1325 12881 1327
rect 12825 1162 12881 1164
rect 12825 1110 12827 1162
rect 12827 1110 12879 1162
rect 12879 1110 12881 1162
rect 12825 1108 12881 1110
rect 12825 944 12881 946
rect 12825 892 12827 944
rect 12827 892 12879 944
rect 12879 892 12881 944
rect 12825 890 12881 892
rect 12825 726 12881 728
rect 12825 674 12827 726
rect 12827 674 12879 726
rect 12879 674 12881 726
rect 12825 672 12881 674
rect 12825 509 12881 511
rect 12825 457 12827 509
rect 12827 457 12879 509
rect 12879 457 12881 509
rect 12825 455 12881 457
rect 12825 291 12881 293
rect 12825 239 12827 291
rect 12827 239 12879 291
rect 12879 239 12881 291
rect 12825 237 12881 239
rect 13398 8400 13454 8402
rect 13398 8348 13400 8400
rect 13400 8348 13452 8400
rect 13452 8348 13454 8400
rect 13398 8346 13454 8348
rect 13398 8183 13454 8185
rect 13398 8131 13400 8183
rect 13400 8131 13452 8183
rect 13452 8131 13454 8183
rect 13398 8129 13454 8131
rect 13398 7965 13454 7967
rect 13398 7913 13400 7965
rect 13400 7913 13452 7965
rect 13452 7913 13454 7965
rect 13398 7911 13454 7913
rect 13398 7748 13454 7750
rect 13398 7696 13400 7748
rect 13400 7696 13452 7748
rect 13452 7696 13454 7748
rect 13398 7694 13454 7696
rect 13398 7530 13454 7532
rect 13398 7478 13400 7530
rect 13400 7478 13452 7530
rect 13452 7478 13454 7530
rect 13398 7476 13454 7478
rect 13398 7312 13454 7314
rect 13398 7260 13400 7312
rect 13400 7260 13452 7312
rect 13452 7260 13454 7312
rect 13398 7258 13454 7260
rect 13398 7094 13454 7096
rect 13398 7042 13400 7094
rect 13400 7042 13452 7094
rect 13452 7042 13454 7094
rect 13398 7040 13454 7042
rect 13398 6877 13454 6879
rect 13398 6825 13400 6877
rect 13400 6825 13452 6877
rect 13452 6825 13454 6877
rect 13398 6823 13454 6825
rect 13398 6659 13454 6661
rect 13398 6607 13400 6659
rect 13400 6607 13452 6659
rect 13452 6607 13454 6659
rect 13398 6605 13454 6607
rect 13398 6442 13454 6444
rect 13398 6390 13400 6442
rect 13400 6390 13452 6442
rect 13452 6390 13454 6442
rect 13398 6388 13454 6390
rect 13513 3991 13569 3993
rect 13513 3939 13515 3991
rect 13515 3939 13567 3991
rect 13567 3939 13569 3991
rect 13513 3937 13569 3939
rect 13513 3773 13569 3775
rect 13513 3721 13515 3773
rect 13515 3721 13567 3773
rect 13567 3721 13569 3773
rect 13513 3719 13569 3721
rect 13513 3556 13569 3558
rect 13513 3504 13515 3556
rect 13515 3504 13567 3556
rect 13567 3504 13569 3556
rect 13513 3502 13569 3504
rect 13513 3338 13569 3340
rect 13513 3286 13515 3338
rect 13515 3286 13567 3338
rect 13567 3286 13569 3338
rect 13513 3284 13569 3286
rect 13513 3120 13569 3122
rect 13513 3068 13515 3120
rect 13515 3068 13567 3120
rect 13567 3068 13569 3120
rect 13513 3066 13569 3068
rect 13513 2903 13569 2905
rect 13513 2851 13515 2903
rect 13515 2851 13567 2903
rect 13567 2851 13569 2903
rect 13513 2849 13569 2851
rect 13513 2685 13569 2687
rect 13513 2633 13515 2685
rect 13515 2633 13567 2685
rect 13567 2633 13569 2685
rect 13513 2631 13569 2633
rect 13513 2468 13569 2470
rect 13513 2416 13515 2468
rect 13515 2416 13567 2468
rect 13567 2416 13569 2468
rect 13513 2414 13569 2416
rect 13513 2250 13569 2252
rect 13513 2198 13515 2250
rect 13515 2198 13567 2250
rect 13567 2198 13569 2250
rect 13513 2196 13569 2198
rect 13513 2032 13569 2034
rect 13513 1980 13515 2032
rect 13515 1980 13567 2032
rect 13567 1980 13569 2032
rect 13513 1978 13569 1980
rect 13513 1814 13569 1816
rect 13513 1762 13515 1814
rect 13515 1762 13567 1814
rect 13567 1762 13569 1814
rect 13513 1760 13569 1762
rect 13513 1597 13569 1599
rect 13513 1545 13515 1597
rect 13515 1545 13567 1597
rect 13567 1545 13569 1597
rect 13513 1543 13569 1545
rect 13513 1379 13569 1381
rect 13513 1327 13515 1379
rect 13515 1327 13567 1379
rect 13567 1327 13569 1379
rect 13513 1325 13569 1327
rect 13513 1162 13569 1164
rect 13513 1110 13515 1162
rect 13515 1110 13567 1162
rect 13567 1110 13569 1162
rect 13513 1108 13569 1110
rect 13513 944 13569 946
rect 13513 892 13515 944
rect 13515 892 13567 944
rect 13567 892 13569 944
rect 13513 890 13569 892
rect 13513 726 13569 728
rect 13513 674 13515 726
rect 13515 674 13567 726
rect 13567 674 13569 726
rect 13513 672 13569 674
rect 13513 509 13569 511
rect 13513 457 13515 509
rect 13515 457 13567 509
rect 13567 457 13569 509
rect 13513 455 13569 457
rect 13513 291 13569 293
rect 13513 239 13515 291
rect 13515 239 13567 291
rect 13567 239 13569 291
rect 13513 237 13569 239
rect -347 -2102 -291 -2046
rect -135 -2102 -79 -2046
<< metal3 >>
rect 2733 16240 13946 16283
rect 2733 16184 6327 16240
rect 6383 16184 6775 16240
rect 6831 16184 7223 16240
rect 7279 16184 7671 16240
rect 7727 16184 8119 16240
rect 8175 16184 8567 16240
rect 8623 16184 8857 16240
rect 8913 16184 9305 16240
rect 9361 16184 9753 16240
rect 9809 16184 10201 16240
rect 10257 16184 10649 16240
rect 10705 16184 11097 16240
rect 11153 16184 11545 16240
rect 11601 16184 11993 16240
rect 12049 16184 12441 16240
rect 12497 16184 12889 16240
rect 12945 16184 13337 16240
rect 13393 16184 13946 16240
rect 2733 16022 13946 16184
rect 2733 15966 6327 16022
rect 6383 15966 6775 16022
rect 6831 15966 7223 16022
rect 7279 15966 7671 16022
rect 7727 15966 8119 16022
rect 8175 15966 8567 16022
rect 8623 15966 8857 16022
rect 8913 15966 9305 16022
rect 9361 15966 9753 16022
rect 9809 15966 10201 16022
rect 10257 15966 10649 16022
rect 10705 15966 11097 16022
rect 11153 15966 11545 16022
rect 11601 15966 11993 16022
rect 12049 15966 12441 16022
rect 12497 15966 12889 16022
rect 12945 15966 13337 16022
rect 13393 15966 13946 16022
rect 2733 15805 13946 15966
rect 2733 15749 6327 15805
rect 6383 15749 6775 15805
rect 6831 15749 7223 15805
rect 7279 15749 7671 15805
rect 7727 15749 8119 15805
rect 8175 15749 8567 15805
rect 8623 15749 8857 15805
rect 8913 15749 9305 15805
rect 9361 15749 9753 15805
rect 9809 15749 10201 15805
rect 10257 15749 10649 15805
rect 10705 15749 11097 15805
rect 11153 15749 11545 15805
rect 11601 15749 11993 15805
rect 12049 15749 12441 15805
rect 12497 15749 12889 15805
rect 12945 15749 13337 15805
rect 13393 15749 13946 15805
rect 2733 15587 13946 15749
rect 2733 15531 6327 15587
rect 6383 15531 6775 15587
rect 6831 15531 7223 15587
rect 7279 15531 7671 15587
rect 7727 15531 8119 15587
rect 8175 15531 8567 15587
rect 8623 15531 8857 15587
rect 8913 15531 9305 15587
rect 9361 15531 9753 15587
rect 9809 15531 10201 15587
rect 10257 15531 10649 15587
rect 10705 15531 11097 15587
rect 11153 15531 11545 15587
rect 11601 15531 11993 15587
rect 12049 15531 12441 15587
rect 12497 15531 12889 15587
rect 12945 15531 13337 15587
rect 13393 15531 13946 15587
rect 2733 15369 13946 15531
rect 2733 15313 6327 15369
rect 6383 15313 6775 15369
rect 6831 15313 7223 15369
rect 7279 15313 7671 15369
rect 7727 15313 8119 15369
rect 8175 15313 8567 15369
rect 8623 15313 8857 15369
rect 8913 15313 9305 15369
rect 9361 15313 9753 15369
rect 9809 15313 10201 15369
rect 10257 15313 10649 15369
rect 10705 15313 11097 15369
rect 11153 15313 11545 15369
rect 11601 15313 11993 15369
rect 12049 15313 12441 15369
rect 12497 15313 12889 15369
rect 12945 15313 13337 15369
rect 13393 15313 13946 15369
rect 2733 15151 13946 15313
rect 2733 15095 6327 15151
rect 6383 15095 6775 15151
rect 6831 15095 7223 15151
rect 7279 15095 7671 15151
rect 7727 15095 8119 15151
rect 8175 15095 8567 15151
rect 8623 15095 8857 15151
rect 8913 15095 9305 15151
rect 9361 15095 9753 15151
rect 9809 15095 10201 15151
rect 10257 15095 10649 15151
rect 10705 15095 11097 15151
rect 11153 15095 11545 15151
rect 11601 15095 11993 15151
rect 12049 15095 12441 15151
rect 12497 15095 12889 15151
rect 12945 15095 13337 15151
rect 13393 15095 13946 15151
rect 2733 14934 13946 15095
rect 2733 14878 6327 14934
rect 6383 14878 6775 14934
rect 6831 14878 7223 14934
rect 7279 14878 7671 14934
rect 7727 14878 8119 14934
rect 8175 14878 8567 14934
rect 8623 14878 8857 14934
rect 8913 14878 9305 14934
rect 9361 14878 9753 14934
rect 9809 14878 10201 14934
rect 10257 14878 10649 14934
rect 10705 14878 11097 14934
rect 11153 14878 11545 14934
rect 11601 14878 11993 14934
rect 12049 14878 12441 14934
rect 12497 14878 12889 14934
rect 12945 14878 13337 14934
rect 13393 14878 13946 14934
rect 2733 14716 13946 14878
rect 2733 14660 6327 14716
rect 6383 14660 6775 14716
rect 6831 14660 7223 14716
rect 7279 14660 7671 14716
rect 7727 14660 8119 14716
rect 8175 14660 8567 14716
rect 8623 14660 8857 14716
rect 8913 14660 9305 14716
rect 9361 14660 9753 14716
rect 9809 14660 10201 14716
rect 10257 14660 10649 14716
rect 10705 14660 11097 14716
rect 11153 14660 11545 14716
rect 11601 14660 11993 14716
rect 12049 14660 12441 14716
rect 12497 14660 12889 14716
rect 12945 14660 13337 14716
rect 13393 14660 13946 14716
rect 2733 14544 13946 14660
rect 5986 11295 13946 11359
rect 5986 11239 6312 11295
rect 6368 11239 13946 11295
rect 5986 11077 13946 11239
rect 5986 11021 6312 11077
rect 6368 11021 13946 11077
rect 5986 10860 13946 11021
rect 5986 10804 6312 10860
rect 6368 10804 13946 10860
rect 5986 10642 13946 10804
rect 5986 10586 6312 10642
rect 6368 10629 13946 10642
rect 6368 10595 13638 10629
rect 6368 10586 8859 10595
rect 5986 10539 8859 10586
rect 8915 10539 9307 10595
rect 9363 10539 9755 10595
rect 9811 10539 10203 10595
rect 10259 10539 10651 10595
rect 10707 10539 11099 10595
rect 11155 10539 11547 10595
rect 11603 10539 11995 10595
rect 12051 10539 12443 10595
rect 12499 10539 12891 10595
rect 12947 10539 13337 10595
rect 13393 10573 13638 10595
rect 13694 10573 13946 10629
rect 13393 10539 13946 10573
rect 5986 10476 13946 10539
rect 5986 10424 8015 10476
rect 5986 10368 6312 10424
rect 6368 10420 8015 10424
rect 8071 10420 8227 10476
rect 8283 10420 13946 10476
rect 6368 10411 13946 10420
rect 6368 10377 13638 10411
rect 6368 10368 8859 10377
rect 5986 10321 8859 10368
rect 8915 10321 9307 10377
rect 9363 10321 9755 10377
rect 9811 10321 10203 10377
rect 10259 10321 10651 10377
rect 10707 10321 11099 10377
rect 11155 10321 11547 10377
rect 11603 10321 11995 10377
rect 12051 10321 12443 10377
rect 12499 10321 12891 10377
rect 12947 10321 13337 10377
rect 13393 10355 13638 10377
rect 13694 10355 13946 10411
rect 13393 10321 13946 10355
rect 5986 10264 13946 10321
rect 5986 10208 7068 10264
rect 7124 10208 7515 10264
rect 7571 10259 13946 10264
rect 7571 10208 8015 10259
rect 5986 10207 8015 10208
rect 5986 10151 6312 10207
rect 6368 10203 8015 10207
rect 8071 10203 8227 10259
rect 8283 10203 13946 10259
rect 6368 10193 13946 10203
rect 6368 10159 13638 10193
rect 6368 10151 8859 10159
rect 5986 10103 8859 10151
rect 8915 10103 9307 10159
rect 9363 10103 9755 10159
rect 9811 10103 10203 10159
rect 10259 10103 10651 10159
rect 10707 10103 11099 10159
rect 11155 10103 11547 10159
rect 11603 10103 11995 10159
rect 12051 10103 12443 10159
rect 12499 10103 12891 10159
rect 12947 10103 13337 10159
rect 13393 10137 13638 10159
rect 13694 10137 13946 10193
rect 13393 10103 13946 10137
rect 5986 10046 13946 10103
rect 5986 9990 7068 10046
rect 7124 9990 7515 10046
rect 7571 10041 13946 10046
rect 7571 9990 8015 10041
rect 5986 9989 8015 9990
rect 5986 9933 6312 9989
rect 6368 9985 8015 9989
rect 8071 9985 8227 10041
rect 8283 9985 13946 10041
rect 6368 9975 13946 9985
rect 6368 9941 13638 9975
rect 6368 9933 8859 9941
rect 5986 9885 8859 9933
rect 8915 9885 9307 9941
rect 9363 9885 9755 9941
rect 9811 9885 10203 9941
rect 10259 9885 10651 9941
rect 10707 9885 11099 9941
rect 11155 9885 11547 9941
rect 11603 9885 11995 9941
rect 12051 9885 12443 9941
rect 12499 9885 12891 9941
rect 12947 9885 13337 9941
rect 13393 9919 13638 9941
rect 13694 9919 13946 9975
rect 13393 9885 13946 9919
rect 5986 9828 13946 9885
rect 5986 9772 7068 9828
rect 7124 9772 7515 9828
rect 7571 9823 13946 9828
rect 7571 9772 8015 9823
rect 5986 9767 8015 9772
rect 8071 9767 8227 9823
rect 8283 9767 13946 9823
rect 5986 9610 13946 9767
rect 5986 9554 7068 9610
rect 7124 9554 7515 9610
rect 7571 9606 13946 9610
rect 7571 9554 8015 9606
rect 5986 9550 8015 9554
rect 8071 9550 8227 9606
rect 8283 9550 13946 9606
rect 5986 9541 13946 9550
rect 5986 9511 10061 9541
rect 11812 9330 15246 9368
rect 11812 9274 11847 9330
rect 11903 9274 12058 9330
rect 12114 9274 12269 9330
rect 12325 9274 12480 9330
rect 12536 9274 12691 9330
rect 12747 9274 12902 9330
rect 12958 9274 13113 9330
rect 13169 9274 15246 9330
rect 6548 9257 6888 9258
rect 10607 9257 10733 9258
rect 11058 9257 11184 9258
rect 11506 9257 11632 9258
rect 6497 9219 11632 9257
rect 6497 9163 6584 9219
rect 6640 9163 6796 9219
rect 6852 9163 10642 9219
rect 10698 9163 11093 9219
rect 11149 9163 11541 9219
rect 11597 9163 11632 9219
rect 6497 9001 11632 9163
rect 6497 8945 6584 9001
rect 6640 8945 6796 9001
rect 6852 8945 10642 9001
rect 10698 8945 11093 9001
rect 11149 8945 11541 9001
rect 11597 8945 11632 9001
rect 6497 8906 11632 8945
rect 11812 9112 15246 9274
rect 11812 9056 11847 9112
rect 11903 9056 12058 9112
rect 12114 9056 12269 9112
rect 12325 9056 12480 9112
rect 12536 9056 12691 9112
rect 12747 9056 12902 9112
rect 12958 9056 13113 9112
rect 13169 9056 15246 9112
rect 11812 8894 15246 9056
rect 11812 8838 11847 8894
rect 11903 8838 12058 8894
rect 12114 8838 12269 8894
rect 12325 8838 12480 8894
rect 12536 8838 12691 8894
rect 12747 8838 12902 8894
rect 12958 8838 13113 8894
rect 13169 8838 15246 8894
rect 4611 8760 4951 8799
rect 4611 8704 4647 8760
rect 4703 8704 4859 8760
rect 4915 8704 4951 8760
rect 4611 8665 4951 8704
rect 11812 8676 15246 8838
rect 11812 8620 11847 8676
rect 11903 8620 12058 8676
rect 12114 8620 12269 8676
rect 12325 8620 12480 8676
rect 12536 8620 12691 8676
rect 12747 8620 12902 8676
rect 12958 8620 13113 8676
rect 13169 8620 15246 8676
rect 11812 8582 15246 8620
rect 5373 8527 8027 8566
rect 5373 8471 5409 8527
rect 5465 8471 5621 8527
rect 5677 8471 7723 8527
rect 7779 8471 7935 8527
rect 7991 8471 8027 8527
rect 5373 8428 8027 8471
rect 8529 8402 13873 8441
rect 8529 8397 12151 8402
rect 8529 8341 8975 8397
rect 9031 8341 9187 8397
rect 9243 8341 9446 8397
rect 9502 8341 9894 8397
rect 9950 8388 12151 8397
rect 9950 8341 10869 8388
rect -206 8260 8076 8335
rect -206 8204 455 8260
rect 511 8204 666 8260
rect 722 8204 876 8260
rect 932 8204 1087 8260
rect 1143 8204 1298 8260
rect 1354 8204 1509 8260
rect 1565 8204 1720 8260
rect 1776 8204 1930 8260
rect 1986 8204 2141 8260
rect 2197 8204 2353 8260
rect 2409 8204 2564 8260
rect 2620 8204 2774 8260
rect 2830 8204 2985 8260
rect 3041 8204 3196 8260
rect 3252 8204 3407 8260
rect 3463 8204 3618 8260
rect 3674 8204 3828 8260
rect 3884 8204 4039 8260
rect 4095 8204 8076 8260
rect -206 8155 8076 8204
rect -206 8099 7116 8155
rect 7172 8099 8076 8155
rect -206 8042 8076 8099
rect -206 7986 455 8042
rect 511 7986 666 8042
rect 722 7986 876 8042
rect 932 7986 1087 8042
rect 1143 7986 1298 8042
rect 1354 7986 1509 8042
rect 1565 7986 1720 8042
rect 1776 7986 1930 8042
rect 1986 7986 2141 8042
rect 2197 7986 2353 8042
rect 2409 7986 2564 8042
rect 2620 7986 2774 8042
rect 2830 7986 2985 8042
rect 3041 7986 3196 8042
rect 3252 7986 3407 8042
rect 3463 7986 3618 8042
rect 3674 7986 3828 8042
rect 3884 7986 4039 8042
rect 4095 7986 8076 8042
rect -206 7937 8076 7986
rect -206 7881 7116 7937
rect 7172 7881 8076 7937
rect -206 7824 8076 7881
rect -206 7768 455 7824
rect 511 7768 666 7824
rect 722 7768 876 7824
rect 932 7768 1087 7824
rect 1143 7768 1298 7824
rect 1354 7768 1509 7824
rect 1565 7768 1720 7824
rect 1776 7768 1930 7824
rect 1986 7768 2141 7824
rect 2197 7768 2353 7824
rect 2409 7768 2564 7824
rect 2620 7768 2774 7824
rect 2830 7768 2985 7824
rect 3041 7768 3196 7824
rect 3252 7768 3407 7824
rect 3463 7768 3618 7824
rect 3674 7768 3828 7824
rect 3884 7768 4039 7824
rect 4095 7768 8076 7824
rect -206 7653 8076 7768
rect 8529 8332 10869 8341
rect 10925 8332 11317 8388
rect 11373 8346 12151 8388
rect 12207 8346 12599 8402
rect 12655 8346 13398 8402
rect 13454 8346 13873 8402
rect 11373 8332 13873 8346
rect 8529 8185 13873 8332
rect 8529 8180 12151 8185
rect 8529 8124 8975 8180
rect 9031 8124 9187 8180
rect 9243 8124 9446 8180
rect 9502 8124 9894 8180
rect 9950 8171 12151 8180
rect 9950 8124 10869 8171
rect 8529 8115 10869 8124
rect 10925 8115 11317 8171
rect 11373 8129 12151 8171
rect 12207 8129 12599 8185
rect 12655 8129 13398 8185
rect 13454 8129 13873 8185
rect 11373 8115 13873 8129
rect 8529 7967 13873 8115
rect 8529 7962 12151 7967
rect 8529 7906 8975 7962
rect 9031 7906 9187 7962
rect 9243 7906 9446 7962
rect 9502 7906 9894 7962
rect 9950 7953 12151 7962
rect 9950 7906 10869 7953
rect 8529 7897 10869 7906
rect 10925 7897 11317 7953
rect 11373 7911 12151 7953
rect 12207 7911 12599 7967
rect 12655 7911 13398 7967
rect 13454 7911 13873 7967
rect 11373 7897 13873 7911
rect 8529 7750 13873 7897
rect 8529 7745 12151 7750
rect 8529 7689 8975 7745
rect 9031 7689 9187 7745
rect 9243 7689 9446 7745
rect 9502 7689 9894 7745
rect 9950 7736 12151 7745
rect 9950 7689 10869 7736
rect 8529 7680 10869 7689
rect 10925 7680 11317 7736
rect 11373 7694 12151 7736
rect 12207 7694 12599 7750
rect 12655 7694 13398 7750
rect 13454 7694 13873 7750
rect 11373 7680 13873 7694
rect 8529 7532 13873 7680
rect 8529 7527 12151 7532
rect 8529 7471 8975 7527
rect 9031 7471 9187 7527
rect 9243 7471 9446 7527
rect 9502 7471 9894 7527
rect 9950 7518 12151 7527
rect 9950 7471 10869 7518
rect 8529 7462 10869 7471
rect 10925 7462 11317 7518
rect 11373 7476 12151 7518
rect 12207 7476 12599 7532
rect 12655 7476 13398 7532
rect 13454 7476 13873 7532
rect 11373 7462 13873 7476
rect -319 7396 5981 7435
rect -319 7340 -283 7396
rect -227 7340 -71 7396
rect -15 7340 5677 7396
rect 5733 7340 5889 7396
rect 5945 7340 5981 7396
rect -319 7301 5981 7340
rect 8529 7314 13873 7462
rect 8529 7309 12151 7314
rect 8529 7253 8975 7309
rect 9031 7253 9187 7309
rect 9243 7253 9446 7309
rect 9502 7253 9894 7309
rect 9950 7300 12151 7309
rect 9950 7253 10869 7300
rect 8529 7244 10869 7253
rect 10925 7244 11317 7300
rect 11373 7258 12151 7300
rect 12207 7258 12599 7314
rect 12655 7258 13398 7314
rect 13454 7258 13873 7314
rect 11373 7244 13873 7258
rect 8529 7181 13873 7244
rect 24 7096 13873 7181
rect 24 7091 12151 7096
rect 24 7077 8975 7091
rect 24 7067 7116 7077
rect 24 7011 4974 7067
rect 5030 7021 7116 7067
rect 7172 7035 8975 7077
rect 9031 7035 9187 7091
rect 9243 7035 9446 7091
rect 9502 7035 9894 7091
rect 9950 7082 12151 7091
rect 9950 7035 10869 7082
rect 7172 7026 10869 7035
rect 10925 7026 11317 7082
rect 11373 7040 12151 7082
rect 12207 7040 12599 7096
rect 12655 7040 13398 7096
rect 13454 7040 13873 7096
rect 11373 7026 13873 7040
rect 7172 7021 13873 7026
rect 5030 7011 13873 7021
rect 24 6879 13873 7011
rect 24 6874 12151 6879
rect 24 6863 8975 6874
rect 24 6807 741 6863
rect 797 6807 952 6863
rect 1008 6807 1162 6863
rect 1218 6807 1373 6863
rect 1429 6807 1584 6863
rect 1640 6807 1795 6863
rect 1851 6807 2006 6863
rect 2062 6807 2216 6863
rect 2272 6807 2427 6863
rect 2483 6807 2639 6863
rect 2695 6807 2850 6863
rect 2906 6807 3060 6863
rect 3116 6807 3271 6863
rect 3327 6807 3482 6863
rect 3538 6807 3693 6863
rect 3749 6807 3904 6863
rect 3960 6807 4114 6863
rect 4170 6807 4325 6863
rect 4381 6859 8975 6863
rect 4381 6849 6384 6859
rect 4381 6807 4974 6849
rect 24 6793 4974 6807
rect 5030 6803 6384 6849
rect 6440 6803 7116 6859
rect 7172 6818 8975 6859
rect 9031 6818 9187 6874
rect 9243 6818 9446 6874
rect 9502 6818 9894 6874
rect 9950 6865 12151 6874
rect 9950 6818 10869 6865
rect 7172 6809 10869 6818
rect 10925 6809 11317 6865
rect 11373 6823 12151 6865
rect 12207 6823 12599 6879
rect 12655 6823 13398 6879
rect 13454 6823 13873 6879
rect 11373 6809 13873 6823
rect 7172 6803 13873 6809
rect 5030 6793 13873 6803
rect 24 6661 13873 6793
rect 24 6656 12151 6661
rect 24 6645 8975 6656
rect 24 6589 741 6645
rect 797 6589 952 6645
rect 1008 6589 1162 6645
rect 1218 6589 1373 6645
rect 1429 6589 1584 6645
rect 1640 6589 1795 6645
rect 1851 6589 2006 6645
rect 2062 6589 2216 6645
rect 2272 6589 2427 6645
rect 2483 6589 2639 6645
rect 2695 6589 2850 6645
rect 2906 6589 3060 6645
rect 3116 6589 3271 6645
rect 3327 6589 3482 6645
rect 3538 6589 3693 6645
rect 3749 6589 3904 6645
rect 3960 6589 4114 6645
rect 4170 6589 4325 6645
rect 4381 6641 8975 6645
rect 4381 6631 6384 6641
rect 4381 6589 4974 6631
rect 24 6575 4974 6589
rect 5030 6585 6384 6631
rect 6440 6585 7116 6641
rect 7172 6600 8975 6641
rect 9031 6600 9187 6656
rect 9243 6600 9446 6656
rect 9502 6600 9894 6656
rect 9950 6647 12151 6656
rect 9950 6600 10869 6647
rect 7172 6591 10869 6600
rect 10925 6591 11317 6647
rect 11373 6605 12151 6647
rect 12207 6605 12599 6661
rect 12655 6605 13398 6661
rect 13454 6605 13873 6661
rect 11373 6591 13873 6605
rect 7172 6585 13873 6591
rect 5030 6575 13873 6585
rect 24 6444 13873 6575
rect 24 6439 12151 6444
rect 24 6423 8975 6439
rect 24 6367 6384 6423
rect 6440 6367 7116 6423
rect 7172 6383 8975 6423
rect 9031 6383 9187 6439
rect 9243 6383 9446 6439
rect 9502 6383 9894 6439
rect 9950 6430 12151 6439
rect 9950 6383 10869 6430
rect 7172 6374 10869 6383
rect 10925 6374 11317 6430
rect 11373 6388 12151 6430
rect 12207 6388 12599 6444
rect 12655 6388 13398 6444
rect 13454 6388 13873 6444
rect 11373 6374 13873 6388
rect 7172 6367 13873 6374
rect 24 6272 13873 6367
rect 562 5972 13878 6102
rect 562 5916 6384 5972
rect 6440 5916 13878 5972
rect 562 5879 13878 5916
rect 562 5823 741 5879
rect 797 5823 952 5879
rect 1008 5823 1162 5879
rect 1218 5823 1373 5879
rect 1429 5823 1584 5879
rect 1640 5823 1795 5879
rect 1851 5823 2006 5879
rect 2062 5823 2216 5879
rect 2272 5823 2427 5879
rect 2483 5823 2639 5879
rect 2695 5823 2850 5879
rect 2906 5823 3060 5879
rect 3116 5823 3271 5879
rect 3327 5823 3482 5879
rect 3538 5823 3693 5879
rect 3749 5823 3904 5879
rect 3960 5823 4114 5879
rect 4170 5823 4325 5879
rect 4381 5823 13878 5879
rect 562 5754 13878 5823
rect 562 5698 6384 5754
rect 6440 5698 13878 5754
rect 562 5661 13878 5698
rect 562 5605 741 5661
rect 797 5605 952 5661
rect 1008 5605 1162 5661
rect 1218 5605 1373 5661
rect 1429 5605 1584 5661
rect 1640 5605 1795 5661
rect 1851 5605 2006 5661
rect 2062 5605 2216 5661
rect 2272 5605 2427 5661
rect 2483 5605 2639 5661
rect 2695 5605 2850 5661
rect 2906 5605 3060 5661
rect 3116 5605 3271 5661
rect 3327 5605 3482 5661
rect 3538 5605 3693 5661
rect 3749 5605 3904 5661
rect 3960 5605 4114 5661
rect 4170 5605 4325 5661
rect 4381 5628 13878 5661
rect 4381 5605 5198 5628
rect 562 5572 5198 5605
rect 5254 5572 13878 5628
rect 562 5410 13878 5572
rect 562 5354 5198 5410
rect 5254 5354 13878 5410
rect 562 5315 13878 5354
rect 158 4939 9731 4995
rect 158 4883 253 4939
rect 309 4883 464 4939
rect 520 4883 675 4939
rect 731 4883 885 4939
rect 941 4883 1096 4939
rect 1152 4883 1307 4939
rect 1363 4883 1518 4939
rect 1574 4883 1729 4939
rect 1785 4883 1939 4939
rect 1995 4883 2150 4939
rect 2206 4883 2361 4939
rect 2417 4883 2572 4939
rect 2628 4883 2783 4939
rect 2839 4883 2994 4939
rect 3050 4883 3205 4939
rect 3261 4883 3416 4939
rect 3472 4883 3627 4939
rect 3683 4883 3837 4939
rect 3893 4883 4048 4939
rect 4104 4883 4259 4939
rect 4315 4883 4470 4939
rect 4526 4883 4681 4939
rect 4737 4883 4891 4939
rect 4947 4883 5102 4939
rect 5158 4883 5313 4939
rect 5369 4883 9731 4939
rect 158 4736 9731 4883
rect 158 4721 9452 4736
rect 158 4665 253 4721
rect 309 4665 464 4721
rect 520 4665 675 4721
rect 731 4665 885 4721
rect 941 4665 1096 4721
rect 1152 4665 1307 4721
rect 1363 4665 1518 4721
rect 1574 4665 1729 4721
rect 1785 4665 1939 4721
rect 1995 4665 2150 4721
rect 2206 4665 2361 4721
rect 2417 4665 2572 4721
rect 2628 4665 2783 4721
rect 2839 4665 2994 4721
rect 3050 4665 3205 4721
rect 3261 4665 3416 4721
rect 3472 4665 3627 4721
rect 3683 4665 3837 4721
rect 3893 4665 4048 4721
rect 4104 4665 4259 4721
rect 4315 4665 4470 4721
rect 4526 4665 4681 4721
rect 4737 4665 4891 4721
rect 4947 4665 5102 4721
rect 5158 4665 5313 4721
rect 5369 4703 9452 4721
rect 5369 4665 8979 4703
rect 158 4647 8979 4665
rect 9035 4647 9191 4703
rect 9247 4680 9452 4703
rect 9508 4680 9731 4736
rect 9247 4647 9731 4680
rect 158 4519 9731 4647
rect 158 4503 9452 4519
rect 158 4447 253 4503
rect 309 4447 464 4503
rect 520 4447 675 4503
rect 731 4447 885 4503
rect 941 4447 1096 4503
rect 1152 4447 1307 4503
rect 1363 4447 1518 4503
rect 1574 4447 1729 4503
rect 1785 4447 1939 4503
rect 1995 4447 2150 4503
rect 2206 4447 2361 4503
rect 2417 4447 2572 4503
rect 2628 4447 2783 4503
rect 2839 4447 2994 4503
rect 3050 4447 3205 4503
rect 3261 4447 3416 4503
rect 3472 4447 3627 4503
rect 3683 4447 3837 4503
rect 3893 4447 4048 4503
rect 4104 4447 4259 4503
rect 4315 4447 4470 4503
rect 4526 4447 4681 4503
rect 4737 4447 4891 4503
rect 4947 4447 5102 4503
rect 5158 4447 5313 4503
rect 5369 4485 9452 4503
rect 5369 4447 8979 4485
rect 158 4429 8979 4447
rect 9035 4429 9191 4485
rect 9247 4463 9452 4485
rect 9508 4463 9731 4519
rect 9247 4429 9731 4463
rect 158 4301 9731 4429
rect 12595 4514 12935 4553
rect 12595 4458 12631 4514
rect 12687 4458 12843 4514
rect 12899 4458 12935 4514
rect 12595 4419 12935 4458
rect 158 4285 9452 4301
rect 158 4229 253 4285
rect 309 4229 464 4285
rect 520 4229 675 4285
rect 731 4229 885 4285
rect 941 4229 1096 4285
rect 1152 4229 1307 4285
rect 1363 4229 1518 4285
rect 1574 4229 1729 4285
rect 1785 4229 1939 4285
rect 1995 4229 2150 4285
rect 2206 4229 2361 4285
rect 2417 4229 2572 4285
rect 2628 4229 2783 4285
rect 2839 4229 2994 4285
rect 3050 4229 3205 4285
rect 3261 4229 3416 4285
rect 3472 4229 3627 4285
rect 3683 4229 3837 4285
rect 3893 4229 4048 4285
rect 4104 4229 4259 4285
rect 4315 4229 4470 4285
rect 4526 4229 4681 4285
rect 4737 4229 4891 4285
rect 4947 4229 5102 4285
rect 5158 4229 5313 4285
rect 5369 4267 9452 4285
rect 5369 4229 8979 4267
rect 158 4211 8979 4229
rect 9035 4211 9191 4267
rect 9247 4245 9452 4267
rect 9508 4245 9731 4301
rect 12596 4352 12935 4419
rect 12596 4256 17136 4352
rect 9247 4211 9731 4245
rect 158 4083 9731 4211
rect 158 4049 9452 4083
rect 158 3993 8979 4049
rect 9035 3993 9191 4049
rect 9247 4027 9452 4049
rect 9508 4077 9731 4083
rect 9508 4027 13783 4077
rect 9247 3993 13783 4027
rect 158 3937 10645 3993
rect 10701 3937 11541 3993
rect 11597 3937 11929 3993
rect 11985 3937 12825 3993
rect 12881 3937 13513 3993
rect 13569 3937 13783 3993
rect 158 3866 13783 3937
rect 158 3810 9452 3866
rect 9508 3810 13783 3866
rect 158 3775 13783 3810
rect 158 3740 10645 3775
rect 9223 3719 10645 3740
rect 10701 3719 11541 3775
rect 11597 3719 11929 3775
rect 11985 3719 12825 3775
rect 12881 3719 13513 3775
rect 13569 3719 13783 3775
rect 9223 3648 13783 3719
rect 9223 3592 9452 3648
rect 9508 3592 13783 3648
rect 9223 3558 13783 3592
rect 9223 3502 10645 3558
rect 10701 3502 11541 3558
rect 11597 3502 11929 3558
rect 11985 3502 12825 3558
rect 12881 3502 13513 3558
rect 13569 3502 13783 3558
rect 9223 3431 13783 3502
rect 9223 3375 9452 3431
rect 9508 3375 13783 3431
rect 9223 3340 13783 3375
rect 71 3065 8829 3327
rect 71 2732 8034 3065
rect 71 2676 2524 2732
rect 2580 2676 2656 2732
rect 2712 2676 2788 2732
rect 2844 2676 2920 2732
rect 2976 2676 3052 2732
rect 3108 2676 3184 2732
rect 3240 2676 3316 2732
rect 3372 2676 3448 2732
rect 3504 2676 3580 2732
rect 3636 2676 3712 2732
rect 3768 2676 3844 2732
rect 3900 2676 3976 2732
rect 4032 2676 4108 2732
rect 4164 2676 4240 2732
rect 4296 2676 4372 2732
rect 4428 2676 4504 2732
rect 4560 2676 4636 2732
rect 4692 2676 4768 2732
rect 4824 2676 4900 2732
rect 4956 2676 5032 2732
rect 5088 2676 5164 2732
rect 5220 2676 5296 2732
rect 5352 2676 5428 2732
rect 5484 2676 5560 2732
rect 5616 2676 5692 2732
rect 5748 2676 5824 2732
rect 5880 2676 5956 2732
rect 6012 2676 6088 2732
rect 6144 2676 6220 2732
rect 6276 2676 6352 2732
rect 6408 2676 6484 2732
rect 6540 2676 6616 2732
rect 6672 2676 6748 2732
rect 6804 2676 6880 2732
rect 6936 2676 7012 2732
rect 7068 2676 7144 2732
rect 7200 2676 7276 2732
rect 7332 2676 7408 2732
rect 7464 2676 7540 2732
rect 7596 2697 8034 2732
rect 8090 2697 8482 3065
rect 8538 2697 8829 3065
rect 7596 2676 8829 2697
rect 71 2600 8829 2676
rect 71 2544 2524 2600
rect 2580 2544 2656 2600
rect 2712 2544 2788 2600
rect 2844 2544 2920 2600
rect 2976 2544 3052 2600
rect 3108 2544 3184 2600
rect 3240 2544 3316 2600
rect 3372 2544 3448 2600
rect 3504 2544 3580 2600
rect 3636 2544 3712 2600
rect 3768 2544 3844 2600
rect 3900 2544 3976 2600
rect 4032 2544 4108 2600
rect 4164 2544 4240 2600
rect 4296 2544 4372 2600
rect 4428 2544 4504 2600
rect 4560 2544 4636 2600
rect 4692 2544 4768 2600
rect 4824 2544 4900 2600
rect 4956 2544 5032 2600
rect 5088 2544 5164 2600
rect 5220 2544 5296 2600
rect 5352 2544 5428 2600
rect 5484 2544 5560 2600
rect 5616 2544 5692 2600
rect 5748 2544 5824 2600
rect 5880 2544 5956 2600
rect 6012 2544 6088 2600
rect 6144 2544 6220 2600
rect 6276 2544 6352 2600
rect 6408 2544 6484 2600
rect 6540 2544 6616 2600
rect 6672 2544 6748 2600
rect 6804 2544 6880 2600
rect 6936 2544 7012 2600
rect 7068 2544 7144 2600
rect 7200 2544 7276 2600
rect 7332 2544 7408 2600
rect 7464 2544 7540 2600
rect 7596 2544 8829 2600
rect 71 2468 8829 2544
rect 71 2412 2524 2468
rect 2580 2412 2656 2468
rect 2712 2412 2788 2468
rect 2844 2412 2920 2468
rect 2976 2412 3052 2468
rect 3108 2412 3184 2468
rect 3240 2412 3316 2468
rect 3372 2412 3448 2468
rect 3504 2412 3580 2468
rect 3636 2412 3712 2468
rect 3768 2412 3844 2468
rect 3900 2412 3976 2468
rect 4032 2412 4108 2468
rect 4164 2412 4240 2468
rect 4296 2412 4372 2468
rect 4428 2412 4504 2468
rect 4560 2412 4636 2468
rect 4692 2412 4768 2468
rect 4824 2412 4900 2468
rect 4956 2412 5032 2468
rect 5088 2412 5164 2468
rect 5220 2412 5296 2468
rect 5352 2412 5428 2468
rect 5484 2412 5560 2468
rect 5616 2412 5692 2468
rect 5748 2412 5824 2468
rect 5880 2412 5956 2468
rect 6012 2412 6088 2468
rect 6144 2412 6220 2468
rect 6276 2412 6352 2468
rect 6408 2412 6484 2468
rect 6540 2412 6616 2468
rect 6672 2412 6748 2468
rect 6804 2412 6880 2468
rect 6936 2412 7012 2468
rect 7068 2412 7144 2468
rect 7200 2412 7276 2468
rect 7332 2412 7408 2468
rect 7464 2412 7540 2468
rect 7596 2412 8829 2468
rect 71 2336 8829 2412
rect 71 2280 2524 2336
rect 2580 2280 2656 2336
rect 2712 2280 2788 2336
rect 2844 2280 2920 2336
rect 2976 2280 3052 2336
rect 3108 2280 3184 2336
rect 3240 2280 3316 2336
rect 3372 2280 3448 2336
rect 3504 2280 3580 2336
rect 3636 2280 3712 2336
rect 3768 2280 3844 2336
rect 3900 2280 3976 2336
rect 4032 2280 4108 2336
rect 4164 2280 4240 2336
rect 4296 2280 4372 2336
rect 4428 2280 4504 2336
rect 4560 2280 4636 2336
rect 4692 2280 4768 2336
rect 4824 2280 4900 2336
rect 4956 2280 5032 2336
rect 5088 2280 5164 2336
rect 5220 2280 5296 2336
rect 5352 2280 5428 2336
rect 5484 2280 5560 2336
rect 5616 2280 5692 2336
rect 5748 2280 5824 2336
rect 5880 2280 5956 2336
rect 6012 2280 6088 2336
rect 6144 2280 6220 2336
rect 6276 2280 6352 2336
rect 6408 2280 6484 2336
rect 6540 2280 6616 2336
rect 6672 2280 6748 2336
rect 6804 2280 6880 2336
rect 6936 2280 7012 2336
rect 7068 2280 7144 2336
rect 7200 2280 7276 2336
rect 7332 2280 7408 2336
rect 7464 2280 7540 2336
rect 7596 2280 8829 2336
rect 71 2265 8829 2280
rect 9223 3284 10645 3340
rect 10701 3284 11541 3340
rect 11597 3284 11929 3340
rect 11985 3284 12825 3340
rect 12881 3284 13513 3340
rect 13569 3284 13783 3340
rect 9223 3213 13783 3284
rect 9223 3157 9452 3213
rect 9508 3157 13783 3213
rect 9223 3122 13783 3157
rect 9223 3066 10645 3122
rect 10701 3066 11541 3122
rect 11597 3066 11929 3122
rect 11985 3066 12825 3122
rect 12881 3066 13513 3122
rect 13569 3066 13783 3122
rect 9223 2995 13783 3066
rect 9223 2939 9452 2995
rect 9508 2939 13783 2995
rect 9223 2905 13783 2939
rect 9223 2849 10645 2905
rect 10701 2849 11541 2905
rect 11597 2849 11929 2905
rect 11985 2849 12825 2905
rect 12881 2849 13513 2905
rect 13569 2849 13783 2905
rect 9223 2778 13783 2849
rect 9223 2722 9452 2778
rect 9508 2722 13783 2778
rect 9223 2687 13783 2722
rect 9223 2631 10645 2687
rect 10701 2631 11541 2687
rect 11597 2631 11929 2687
rect 11985 2631 12825 2687
rect 12881 2631 13513 2687
rect 13569 2631 13783 2687
rect 9223 2560 13783 2631
rect 9223 2504 9452 2560
rect 9508 2504 13783 2560
rect 9223 2470 13783 2504
rect 9223 2414 10645 2470
rect 10701 2414 11541 2470
rect 11597 2414 11929 2470
rect 11985 2414 12825 2470
rect 12881 2414 13513 2470
rect 13569 2414 13783 2470
rect 9223 2342 13783 2414
rect 9223 2286 9452 2342
rect 9508 2286 13783 2342
rect 9223 2252 13783 2286
rect 9223 2196 10645 2252
rect 10701 2196 11541 2252
rect 11597 2196 11929 2252
rect 11985 2196 12825 2252
rect 12881 2196 13513 2252
rect 13569 2196 13783 2252
rect 9223 2125 13783 2196
rect 9223 2069 9452 2125
rect 9508 2069 13783 2125
rect 9223 2034 13783 2069
rect 9223 1978 10645 2034
rect 10701 1978 11541 2034
rect 11597 1978 11929 2034
rect 11985 1978 12825 2034
rect 12881 1978 13513 2034
rect 13569 1978 13783 2034
rect 9223 1907 13783 1978
rect 9223 1851 9452 1907
rect 9508 1851 13783 1907
rect 9223 1816 13783 1851
rect 9223 1760 10645 1816
rect 10701 1760 11541 1816
rect 11597 1760 11929 1816
rect 11985 1760 12825 1816
rect 12881 1760 13513 1816
rect 13569 1760 13783 1816
rect 9223 1689 13783 1760
rect 9223 1633 9452 1689
rect 9508 1633 13783 1689
rect 9223 1599 13783 1633
rect 9223 1543 10645 1599
rect 10701 1543 11541 1599
rect 11597 1543 11929 1599
rect 11985 1543 12825 1599
rect 12881 1543 13513 1599
rect 13569 1543 13783 1599
rect 9223 1472 13783 1543
rect 9223 1450 9452 1472
rect -930 1416 9452 1450
rect 9508 1416 13783 1472
rect -930 1381 13783 1416
rect -930 1325 10645 1381
rect 10701 1325 11541 1381
rect 11597 1325 11929 1381
rect 11985 1325 12825 1381
rect 12881 1325 13513 1381
rect 13569 1325 13783 1381
rect -930 1254 13783 1325
rect -930 1198 9452 1254
rect 9508 1198 13783 1254
rect -930 1167 13783 1198
rect 9223 1164 13783 1167
rect 9223 1108 10645 1164
rect 10701 1108 11541 1164
rect 11597 1108 11929 1164
rect 11985 1108 12825 1164
rect 12881 1108 13513 1164
rect 13569 1108 13783 1164
rect 9223 1037 13783 1108
rect 9223 981 9452 1037
rect 9508 981 13783 1037
rect 9223 946 13783 981
rect 9223 890 10645 946
rect 10701 890 11541 946
rect 11597 890 11929 946
rect 11985 890 12825 946
rect 12881 890 13513 946
rect 13569 890 13783 946
rect 9223 819 13783 890
rect 9223 763 9452 819
rect 9508 763 13783 819
rect 9223 728 13783 763
rect 9223 672 10645 728
rect 10701 672 11541 728
rect 11597 672 11929 728
rect 11985 672 12825 728
rect 12881 672 13513 728
rect 13569 672 13783 728
rect 9223 601 13783 672
rect 9223 545 9452 601
rect 9508 545 13783 601
rect 9223 511 13783 545
rect 9223 455 10645 511
rect 10701 455 11541 511
rect 11597 455 11929 511
rect 11985 455 12825 511
rect 12881 455 13513 511
rect 13569 455 13783 511
rect 9223 384 13783 455
rect 9223 328 9452 384
rect 9508 328 13783 384
rect 9223 293 13783 328
rect 9223 237 10645 293
rect 10701 237 11541 293
rect 11597 237 11929 293
rect 11985 237 12825 293
rect 12881 237 13513 293
rect 13569 237 13783 293
rect 9223 180 13783 237
rect -930 -109 8587 175
rect -17790 -1261 17624 -806
rect -17790 -1901 15799 -1550
rect -383 -2008 -43 -2007
rect -14200 -2046 15799 -2008
rect -14200 -2102 -347 -2046
rect -291 -2102 -135 -2046
rect -79 -2102 15799 -2046
rect -14200 -2141 15799 -2102
use CON_64x8m81  CON_64x8m81_0
timestamp 1755005639
transform 1 0 6373 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_1
timestamp 1755005639
transform 1 0 6531 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_2
timestamp 1755005639
transform 1 0 6689 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_3
timestamp 1755005639
transform 1 0 6689 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_4
timestamp 1755005639
transform 1 0 6215 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_5
timestamp 1755005639
transform 1 0 6373 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_6
timestamp 1755005639
transform 1 0 6531 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_7
timestamp 1755005639
transform 1 0 6061 0 1 11988
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_8
timestamp 1755005639
transform 1 0 6061 0 1 12151
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_9
timestamp 1755005639
transform 1 0 6061 0 1 12314
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_10
timestamp 1755005639
transform 1 0 6061 0 1 12478
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_11
timestamp 1755005639
transform 1 0 6061 0 1 12641
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_12
timestamp 1755005639
transform 1 0 6061 0 1 12804
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_13
timestamp 1755005639
transform 1 0 6061 0 1 12967
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_14
timestamp 1755005639
transform 1 0 6061 0 1 13130
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_15
timestamp 1755005639
transform 1 0 6061 0 1 13294
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_16
timestamp 1755005639
transform 1 0 6061 0 1 13457
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_17
timestamp 1755005639
transform 1 0 6061 0 1 13620
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_18
timestamp 1755005639
transform 1 0 6061 0 1 13783
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_19
timestamp 1755005639
transform 1 0 6061 0 1 13947
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_20
timestamp 1755005639
transform 1 0 6061 0 1 14110
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_21
timestamp 1755005639
transform 1 0 6061 0 1 14273
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_22
timestamp 1755005639
transform 1 0 6061 0 1 14436
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_23
timestamp 1755005639
transform 1 0 6061 0 1 14599
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_24
timestamp 1755005639
transform 1 0 6061 0 1 14763
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_25
timestamp 1755005639
transform 1 0 6061 0 1 14926
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_26
timestamp 1755005639
transform 1 0 6061 0 1 15089
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_27
timestamp 1755005639
transform 1 0 6061 0 1 15252
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_28
timestamp 1755005639
transform 1 0 6061 0 1 15416
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_29
timestamp 1755005639
transform 1 0 6061 0 1 15579
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_30
timestamp 1755005639
transform 1 0 6061 0 1 15742
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_31
timestamp 1755005639
transform 1 0 6061 0 1 15905
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_32
timestamp 1755005639
transform 1 0 6061 0 1 16069
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_33
timestamp 1755005639
transform 1 0 6215 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_34
timestamp 1755005639
transform 1 0 6847 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_35
timestamp 1755005639
transform 1 0 7005 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_36
timestamp 1755005639
transform 1 0 7163 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_37
timestamp 1755005639
transform 1 0 7321 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_38
timestamp 1755005639
transform 1 0 7480 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_39
timestamp 1755005639
transform 1 0 7638 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_40
timestamp 1755005639
transform 1 0 7796 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_41
timestamp 1755005639
transform 1 0 7954 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_42
timestamp 1755005639
transform 1 0 8112 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_43
timestamp 1755005639
transform 1 0 8270 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_44
timestamp 1755005639
transform 1 0 8428 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_45
timestamp 1755005639
transform 1 0 8586 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_46
timestamp 1755005639
transform 1 0 8744 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_47
timestamp 1755005639
transform 1 0 8903 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_48
timestamp 1755005639
transform 1 0 9061 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_49
timestamp 1755005639
transform 1 0 9219 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_50
timestamp 1755005639
transform 1 0 9377 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_51
timestamp 1755005639
transform 1 0 9535 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_52
timestamp 1755005639
transform 1 0 9693 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_53
timestamp 1755005639
transform 1 0 9851 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_54
timestamp 1755005639
transform 1 0 10009 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_55
timestamp 1755005639
transform 1 0 10167 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_56
timestamp 1755005639
transform 1 0 6847 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_57
timestamp 1755005639
transform 1 0 7005 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_58
timestamp 1755005639
transform 1 0 7163 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_59
timestamp 1755005639
transform 1 0 7321 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_60
timestamp 1755005639
transform 1 0 7480 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_61
timestamp 1755005639
transform 1 0 7638 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_62
timestamp 1755005639
transform 1 0 7796 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_63
timestamp 1755005639
transform 1 0 7954 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_64
timestamp 1755005639
transform 1 0 8112 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_65
timestamp 1755005639
transform 1 0 8270 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_66
timestamp 1755005639
transform 1 0 8428 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_67
timestamp 1755005639
transform 1 0 8586 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_68
timestamp 1755005639
transform 1 0 8744 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_69
timestamp 1755005639
transform 1 0 8903 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_70
timestamp 1755005639
transform 1 0 9061 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_71
timestamp 1755005639
transform 1 0 9219 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_72
timestamp 1755005639
transform 1 0 9377 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_73
timestamp 1755005639
transform 1 0 9535 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_74
timestamp 1755005639
transform 1 0 9693 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_75
timestamp 1755005639
transform 1 0 9851 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_76
timestamp 1755005639
transform 1 0 10009 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_77
timestamp 1755005639
transform 1 0 10167 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_78
timestamp 1755005639
transform 1 0 13655 0 1 11988
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_79
timestamp 1755005639
transform 1 0 13655 0 1 12151
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_80
timestamp 1755005639
transform 1 0 13655 0 1 12314
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_81
timestamp 1755005639
transform 1 0 13655 0 1 12478
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_82
timestamp 1755005639
transform 1 0 13655 0 1 12641
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_83
timestamp 1755005639
transform 1 0 13655 0 1 12804
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_84
timestamp 1755005639
transform 1 0 13655 0 1 12967
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_85
timestamp 1755005639
transform 1 0 13655 0 1 13130
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_86
timestamp 1755005639
transform 1 0 13655 0 1 13294
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_87
timestamp 1755005639
transform 1 0 13655 0 1 13457
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_88
timestamp 1755005639
transform 1 0 13655 0 1 13620
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_89
timestamp 1755005639
transform 1 0 13655 0 1 13783
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_90
timestamp 1755005639
transform 1 0 13655 0 1 13947
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_91
timestamp 1755005639
transform 1 0 13655 0 1 14110
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_92
timestamp 1755005639
transform 1 0 13655 0 1 14273
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_93
timestamp 1755005639
transform 1 0 13655 0 1 14436
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_94
timestamp 1755005639
transform 1 0 13655 0 1 14599
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_95
timestamp 1755005639
transform 1 0 13655 0 1 14763
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_96
timestamp 1755005639
transform 1 0 13655 0 1 14926
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_97
timestamp 1755005639
transform 1 0 13655 0 1 15089
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_98
timestamp 1755005639
transform 1 0 13655 0 1 15252
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_99
timestamp 1755005639
transform 1 0 13655 0 1 15416
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_100
timestamp 1755005639
transform 1 0 13655 0 1 15579
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_101
timestamp 1755005639
transform 1 0 13655 0 1 15742
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_102
timestamp 1755005639
transform 1 0 13655 0 1 15905
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_103
timestamp 1755005639
transform 1 0 13655 0 1 16069
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_104
timestamp 1755005639
transform 1 0 10326 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_105
timestamp 1755005639
transform 1 0 10484 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_106
timestamp 1755005639
transform 1 0 10642 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_107
timestamp 1755005639
transform 1 0 10800 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_108
timestamp 1755005639
transform 1 0 10958 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_109
timestamp 1755005639
transform 1 0 11116 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_110
timestamp 1755005639
transform 1 0 11274 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_111
timestamp 1755005639
transform 1 0 11432 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_112
timestamp 1755005639
transform 1 0 11590 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_113
timestamp 1755005639
transform 1 0 11749 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_114
timestamp 1755005639
transform 1 0 11907 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_115
timestamp 1755005639
transform 1 0 12065 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_116
timestamp 1755005639
transform 1 0 12223 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_117
timestamp 1755005639
transform 1 0 12381 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_118
timestamp 1755005639
transform 1 0 12539 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_119
timestamp 1755005639
transform 1 0 12697 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_120
timestamp 1755005639
transform 1 0 12855 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_121
timestamp 1755005639
transform 1 0 13013 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_122
timestamp 1755005639
transform 1 0 13172 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_123
timestamp 1755005639
transform 1 0 13330 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_124
timestamp 1755005639
transform 1 0 13488 0 1 11938
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_125
timestamp 1755005639
transform 1 0 10326 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_126
timestamp 1755005639
transform 1 0 10484 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_127
timestamp 1755005639
transform 1 0 10642 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_128
timestamp 1755005639
transform 1 0 10800 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_129
timestamp 1755005639
transform 1 0 10958 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_130
timestamp 1755005639
transform 1 0 11116 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_131
timestamp 1755005639
transform 1 0 11274 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_132
timestamp 1755005639
transform 1 0 11432 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_133
timestamp 1755005639
transform 1 0 11590 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_134
timestamp 1755005639
transform 1 0 11749 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_135
timestamp 1755005639
transform 1 0 11907 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_136
timestamp 1755005639
transform 1 0 12065 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_137
timestamp 1755005639
transform 1 0 12223 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_138
timestamp 1755005639
transform 1 0 12381 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_139
timestamp 1755005639
transform 1 0 12539 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_140
timestamp 1755005639
transform 1 0 12697 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_141
timestamp 1755005639
transform 1 0 12855 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_142
timestamp 1755005639
transform 1 0 13013 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_143
timestamp 1755005639
transform 1 0 13172 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_144
timestamp 1755005639
transform 1 0 13330 0 1 16250
box 0 0 1 1
use CON_64x8m81  CON_64x8m81_145
timestamp 1755005639
transform 1 0 13488 0 1 16250
box 0 0 1 1
use M1_NACTIVE4310589983264_64x8m81  M1_NACTIVE4310589983264_64x8m81_0
timestamp 1755005639
transform 1 0 5593 0 1 2510
box 0 0 1 1
use M1_NWELL$$47635500_R90_64x8m81  M1_NWELL$$47635500_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 9084 1 0 7595
box 0 0 1 1
use M1_NWELL$$48078892_64x8m81  M1_NWELL$$48078892_64x8m81_0
timestamp 1755005639
transform -1 0 11140 0 -1 9472
box 0 0 1 1
use M1_NWELL$$48079916_R90_64x8m81  M1_NWELL$$48079916_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 13354 1 0 7187
box 0 0 1 1
use M1_NWELL$$48080940_64x8m81  M1_NWELL$$48080940_64x8m81_0
timestamp 1755005639
transform 1 0 7479 0 1 12591
box 0 0 1 1
use M1_NWELL$$169758764_64x8m81  M1_NWELL$$169758764_64x8m81_0
timestamp 1755005639
transform 1 0 2580 0 1 6728
box 0 0 1 1
use M1_PACTIVE$$48_R90_64x8m81  M1_PACTIVE$$48_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 6346 1 0 10149
box 0 0 1 1
use M1_PACTIVE$$480_R90_64x8m81  M1_PACTIVE$$480_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 13666 1 0 10757
box 0 0 1 1
use M1_PACTIVE$$4807_R90_64x8m81  M1_PACTIVE$$4807_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 8147 1 0 9914
box 0 0 1 1
use M1_PACTIVE$$48067628_64x8m81  M1_PACTIVE$$48067628_64x8m81_0
timestamp 1755005639
transform 1 0 4139 0 1 8608
box 0 0 1 1
use M1_PACTIVE$$48072748_64x8m81  M1_PACTIVE$$48072748_64x8m81_0
timestamp 1755005639
transform -1 0 7216 0 -1 11455
box 0 0 1 1
use M1_PACTIVE$$169762860_64x8m81  M1_PACTIVE$$169762860_64x8m81_0
timestamp 1755005639
transform 1 0 2580 0 1 5745
box 0 0 1 1
use M1_PACTIVE4310589983270_64x8m81  M1_PACTIVE4310589983270_64x8m81_0
timestamp 1755005639
transform 1 0 4037 0 1 4674
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_0
timestamp 1755005639
transform 1 0 7157 0 1 5994
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_1
timestamp 1755005639
transform 1 0 7816 0 1 6010
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_2
timestamp 1755005639
transform 1 0 8088 0 1 3534
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_3
timestamp 1755005639
transform 1 0 7570 0 1 3534
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_4
timestamp 1755005639
transform 1 0 6930 0 1 3534
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_5
timestamp 1755005639
transform -1 0 5077 0 1 6001
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_6
timestamp 1755005639
transform 1 0 6206 0 1 3534
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_7
timestamp 1755005639
transform 1 0 5279 0 1 7055
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_8
timestamp 1755005639
transform 1 0 7627 0 1 7409
box 0 0 1 1
use M1_POLY2$$44754988_64x8m81  M1_POLY2$$44754988_64x8m81_0
timestamp 1755005639
transform 1 0 7851 0 1 7880
box 0 0 1 1
use M1_POLY2$$46559276_64x8m81_0  M1_POLY2$$46559276_64x8m81_0_0
timestamp 1755005639
transform 1 0 5447 0 1 3534
box 0 0 1 1
use M1_POLY2$$46559276_64x8m81_0  M1_POLY2$$46559276_64x8m81_0_1
timestamp 1755005639
transform 1 0 6342 0 1 7368
box 0 0 1 1
use M1_POLY24310589983234_64x8m81  M1_POLY24310589983234_64x8m81_0
timestamp 1755005639
transform 1 0 12411 0 1 4483
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_0
timestamp 1755005639
transform 1 0 12741 0 1 4265
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_1
timestamp 1755005639
transform 1 0 12069 0 1 4265
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_2
timestamp 1755005639
transform 1 0 11457 0 1 4514
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_3
timestamp 1755005639
transform 1 0 10786 0 1 4514
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_4
timestamp 1755005639
transform 1 0 5811 0 1 5788
box 0 0 1 1
use M1_POLY24310589983237_64x8m81  M1_POLY24310589983237_64x8m81_0
timestamp 1755005639
transform 1 0 11119 0 1 4296
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_0
timestamp 1755005639
transform 1 0 9814 0 1 5025
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_1
timestamp 1755005639
transform 1 0 9591 0 1 5025
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_2
timestamp 1755005639
transform 1 0 10038 0 1 5025
box 0 0 1 1
use M1_POLY24310589983262_64x8m81  M1_POLY24310589983262_64x8m81_0
timestamp 1755005639
transform 1 0 11141 0 1 12181
box 0 0 1 1
use M1_POLY24310589983263_64x8m81  M1_POLY24310589983263_64x8m81_0
timestamp 1755005639
transform 1 0 11109 0 1 11415
box 0 0 1 1
use M1_POLY24310589983268_64x8m81  M1_POLY24310589983268_64x8m81_0
timestamp 1755005639
transform 1 0 7484 0 1 13359
box 0 0 1 1
use M1_POLY24310589983269_64x8m81  M1_POLY24310589983269_64x8m81_0
timestamp 1755005639
transform 1 0 7212 0 1 11137
box 0 0 1 1
use M1_PSUB$$48310316_R90_64x8m81  M1_PSUB$$48310316_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 13455 1 0 2086
box 0 0 1 1
use M1_PSUB$$48311340_R90_64x8m81  M1_PSUB$$48311340_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 9028 1 0 2330
box 0 0 1 1
use M1_PSUB$$48312364_64x8m81  M1_PSUB$$48312364_64x8m81_0
timestamp 1755005639
transform 1 0 11321 0 1 -37
box 0 0 1 1
use M1_PSUB$$169764908_64x8m81  M1_PSUB$$169764908_64x8m81_0
timestamp 1755005639
transform -1 0 2323 0 1 8120
box 0 0 1 1
use M2_M1$$34864172_64x8m81  M2_M1$$34864172_64x8m81_0
timestamp 1755005639
transform 1 0 11727 0 1 4264
box 0 0 1 1
use M2_M1$$34864172_64x8m81  M2_M1$$34864172_64x8m81_1
timestamp 1755005639
transform 1 0 12765 0 1 4486
box 0 0 1 1
use M2_M1$$34864172_64x8m81  M2_M1$$34864172_64x8m81_2
timestamp 1755005639
transform 1 0 4972 0 1 5994
box 0 0 1 1
use M2_M1$$34864172_64x8m81  M2_M1$$34864172_64x8m81_3
timestamp 1755005639
transform 1 0 5494 0 1 3532
box 0 0 1 1
use M2_M1$$34864172_R90_64x8m81  M2_M1$$34864172_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 10036 1 0 5026
box 0 0 1 1
use M2_M1$$34864172_R90_64x8m81  M2_M1$$34864172_R90_64x8m81_1
timestamp 1755005639
transform 0 -1 9810 1 0 5026
box 0 0 1 1
use M2_M1$$34864172_R90_64x8m81  M2_M1$$34864172_R90_64x8m81_2
timestamp 1755005639
transform 0 -1 6920 1 0 5983
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_0
timestamp 1755005639
transform -1 0 5226 0 1 5491
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_1
timestamp 1755005639
transform 1 0 6412 0 1 5835
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_2
timestamp 1755005639
transform -1 0 5457 0 1 6595
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_3
timestamp 1755005639
transform 1 0 7857 0 1 7948
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_4
timestamp 1755005639
transform 1 0 9698 0 1 8855
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_5
timestamp 1755005639
transform 1 0 10148 0 1 8855
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_6
timestamp 1755005639
transform 1 0 7144 0 1 8018
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_7
timestamp 1755005639
transform 1 0 7857 0 1 7293
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_8
timestamp 1755005639
transform 1 0 6920 0 1 7087
box 0 0 1 1
use M2_M1$$43375660_R90_64x8m81  M2_M1$$43375660_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 8755 1 0 5182
box 0 0 1 1
use M2_M1$$43375660_R90_64x8m81  M2_M1$$43375660_R90_64x8m81_1
timestamp 1755005639
transform 0 -1 6324 1 0 7365
box 0 0 1 1
use M2_M1$$43375660_R270_64x8m81  M2_M1$$43375660_R270_64x8m81_0
timestamp 1755005639
transform 0 -1 5543 -1 0 7887
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_0
timestamp 1755005639
transform 1 0 6355 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_1
timestamp 1755005639
transform 1 0 7699 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_2
timestamp 1755005639
transform 1 0 8147 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_3
timestamp 1755005639
transform 1 0 9781 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_4
timestamp 1755005639
transform 1 0 9333 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_5
timestamp 1755005639
transform 1 0 8885 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_6
timestamp 1755005639
transform 1 0 8595 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_7
timestamp 1755005639
transform 1 0 6803 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_8
timestamp 1755005639
transform 1 0 7251 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_9
timestamp 1755005639
transform 1 0 11573 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_10
timestamp 1755005639
transform 1 0 11125 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_11
timestamp 1755005639
transform 1 0 10677 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_12
timestamp 1755005639
transform 1 0 13365 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_13
timestamp 1755005639
transform 1 0 12917 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_14
timestamp 1755005639
transform 1 0 12469 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_15
timestamp 1755005639
transform 1 0 12021 0 1 15450
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_16
timestamp 1755005639
transform 1 0 10229 0 1 15450
box 0 0 1 1
use M2_M1$$43377708_64x8m81  M2_M1$$43377708_64x8m81_0
timestamp 1755005639
transform 1 0 12693 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_64x8m81  M2_M1$$43377708_64x8m81_1
timestamp 1755005639
transform 1 0 12245 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_64x8m81  M2_M1$$43377708_64x8m81_2
timestamp 1755005639
transform 1 0 11797 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_64x8m81  M2_M1$$43377708_64x8m81_3
timestamp 1755005639
transform 1 0 13141 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_64x8m81  M2_M1$$43377708_64x8m81_4
timestamp 1755005639
transform 1 0 11349 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_64x8m81  M2_M1$$43377708_64x8m81_5
timestamp 1755005639
transform 1 0 10901 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_64x8m81  M2_M1$$43377708_64x8m81_6
timestamp 1755005639
transform 1 0 10453 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_64x8m81  M2_M1$$43377708_64x8m81_7
timestamp 1755005639
transform 1 0 9109 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_64x8m81  M2_M1$$43377708_64x8m81_8
timestamp 1755005639
transform 1 0 9557 0 1 10625
box 0 0 1 1
use M2_M1$$43377708_64x8m81  M2_M1$$43377708_64x8m81_9
timestamp 1755005639
transform 1 0 10005 0 1 10625
box 0 0 1 1
use M2_M1$$43378732_64x8m81  M2_M1$$43378732_64x8m81_0
timestamp 1755005639
transform 1 0 6577 0 1 13972
box 0 0 1 1
use M2_M1$$43378732_64x8m81  M2_M1$$43378732_64x8m81_1
timestamp 1755005639
transform 1 0 7025 0 1 13972
box 0 0 1 1
use M2_M1$$43378732_64x8m81  M2_M1$$43378732_64x8m81_2
timestamp 1755005639
transform 1 0 7921 0 1 13972
box 0 0 1 1
use M2_M1$$43378732_64x8m81  M2_M1$$43378732_64x8m81_3
timestamp 1755005639
transform 1 0 8369 0 1 13972
box 0 0 1 1
use M2_M1$$43378732_64x8m81  M2_M1$$43378732_64x8m81_4
timestamp 1755005639
transform 1 0 7473 0 1 13972
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_0
timestamp 1755005639
transform 1 0 12405 0 1 5060
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_1
timestamp 1755005639
transform 1 0 12853 0 1 5060
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_2
timestamp 1755005639
transform 1 0 11957 0 1 5060
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_3
timestamp 1755005639
transform 1 0 13365 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_4
timestamp 1755005639
transform 1 0 12919 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_5
timestamp 1755005639
transform 1 0 11575 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_6
timestamp 1755005639
transform 1 0 12023 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_7
timestamp 1755005639
transform 1 0 12471 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_8
timestamp 1755005639
transform 1 0 10679 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_9
timestamp 1755005639
transform 1 0 11127 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_10
timestamp 1755005639
transform 1 0 13666 0 1 10274
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_11
timestamp 1755005639
transform 1 0 7543 0 1 9909
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_12
timestamp 1755005639
transform 1 0 9783 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_13
timestamp 1755005639
transform 1 0 9335 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_14
timestamp 1755005639
transform 1 0 8887 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_15
timestamp 1755005639
transform 1 0 7096 0 1 9909
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_16
timestamp 1755005639
transform 1 0 10231 0 1 10240
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_17
timestamp 1755005639
transform 1 0 7144 0 1 6722
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_0
timestamp 1755005639
transform 1 0 6412 0 1 6613
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_1
timestamp 1755005639
transform -1 0 5002 0 1 6821
box 0 0 1 1
use M2_M1$$45013036_64x8m81  M2_M1$$45013036_64x8m81_0
timestamp 1755005639
transform 1 0 6920 0 1 13310
box 0 0 1 1
use M2_M1$$45013036_64x8m81  M2_M1$$45013036_64x8m81_1
timestamp 1755005639
transform 1 0 6950 0 1 11174
box 0 0 1 1
use M2_M1$$47500332_64x8m81  M2_M1$$47500332_64x8m81_0
timestamp 1755005639
transform 1 0 13426 0 1 7395
box 0 0 1 1
use M2_M1$$47500332_64x8m81  M2_M1$$47500332_64x8m81_1
timestamp 1755005639
transform 1 0 12179 0 1 7395
box 0 0 1 1
use M2_M1$$47500332_64x8m81  M2_M1$$47500332_64x8m81_2
timestamp 1755005639
transform 1 0 12627 0 1 7395
box 0 0 1 1
use M2_M1$$47500332_64x8m81  M2_M1$$47500332_64x8m81_3
timestamp 1755005639
transform 1 0 9922 0 1 7390
box 0 0 1 1
use M2_M1$$47500332_64x8m81  M2_M1$$47500332_64x8m81_4
timestamp 1755005639
transform 1 0 9474 0 1 7390
box 0 0 1 1
use M2_M1$$47500332_64x8m81  M2_M1$$47500332_64x8m81_5
timestamp 1755005639
transform 1 0 11345 0 1 7381
box 0 0 1 1
use M2_M1$$47500332_64x8m81  M2_M1$$47500332_64x8m81_6
timestamp 1755005639
transform 1 0 10897 0 1 7381
box 0 0 1 1
use M2_M1$$47515692_64x8m81  M2_M1$$47515692_64x8m81_0
timestamp 1755005639
transform 1 0 6340 0 1 10614
box 0 0 1 1
use M2_M1$$47515692_64x8m81  M2_M1$$47515692_64x8m81_1
timestamp 1755005639
transform 1 0 7767 0 1 10236
box 0 0 1 1
use M2_M1$$47515692_64x8m81  M2_M1$$47515692_64x8m81_2
timestamp 1755005639
transform 1 0 7319 0 1 10236
box 0 0 1 1
use M2_M1$$47515692_64x8m81  M2_M1$$47515692_64x8m81_3
timestamp 1755005639
transform 1 0 6872 0 1 10236
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_0
timestamp 1755005639
transform 1 0 11121 0 1 3167
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_1
timestamp 1755005639
transform 1 0 12405 0 1 3167
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_2
timestamp 1755005639
transform 1 0 10005 0 1 13439
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_3
timestamp 1755005639
transform 1 0 9557 0 1 13439
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_4
timestamp 1755005639
transform 1 0 9109 0 1 13439
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_5
timestamp 1755005639
transform 1 0 13141 0 1 13439
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_6
timestamp 1755005639
transform 1 0 11797 0 1 13439
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_7
timestamp 1755005639
transform 1 0 12245 0 1 13439
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_8
timestamp 1755005639
transform 1 0 12693 0 1 13439
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_9
timestamp 1755005639
transform 1 0 10453 0 1 13439
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_10
timestamp 1755005639
transform 1 0 10901 0 1 13439
box 0 0 1 1
use M2_M1$$48217132_64x8m81  M2_M1$$48217132_64x8m81_11
timestamp 1755005639
transform 1 0 11349 0 1 13439
box 0 0 1 1
use M2_M1$$48218156_64x8m81  M2_M1$$48218156_64x8m81_0
timestamp 1755005639
transform 1 0 10117 0 1 12144
box 0 0 1 1
use M2_M1$$48218156_64x8m81  M2_M1$$48218156_64x8m81_1
timestamp 1755005639
transform 1 0 10117 0 1 11451
box 0 0 1 1
use M2_M1$$48219180_64x8m81  M2_M1$$48219180_64x8m81_0
timestamp 1755005639
transform 1 0 9113 0 1 4348
box 0 0 1 1
use M2_M1$$48220204_64x8m81  M2_M1$$48220204_64x8m81_0
timestamp 1755005639
transform 1 0 9109 0 1 7390
box 0 0 1 1
use M2_M1$$48221228_64x8m81  M2_M1$$48221228_64x8m81_0
timestamp 1755005639
transform 1 0 13541 0 1 2115
box 0 0 1 1
use M2_M1$$48221228_64x8m81  M2_M1$$48221228_64x8m81_1
timestamp 1755005639
transform 1 0 11569 0 1 2115
box 0 0 1 1
use M2_M1$$48221228_64x8m81  M2_M1$$48221228_64x8m81_2
timestamp 1755005639
transform 1 0 11957 0 1 2115
box 0 0 1 1
use M2_M1$$48221228_64x8m81  M2_M1$$48221228_64x8m81_3
timestamp 1755005639
transform 1 0 12853 0 1 2115
box 0 0 1 1
use M2_M1$$48221228_64x8m81  M2_M1$$48221228_64x8m81_4
timestamp 1755005639
transform 1 0 10673 0 1 2115
box 0 0 1 1
use M2_M1$$48222252_64x8m81  M2_M1$$48222252_64x8m81_0
timestamp 1755005639
transform 1 0 11569 0 1 7003
box 0 0 1 1
use M2_M1$$48222252_64x8m81  M2_M1$$48222252_64x8m81_1
timestamp 1755005639
transform 1 0 10673 0 1 7003
box 0 0 1 1
use M2_M1$$48222252_64x8m81  M2_M1$$48222252_64x8m81_2
timestamp 1755005639
transform 1 0 11121 0 1 7003
box 0 0 1 1
use M2_M1$$48224300_64x8m81  M2_M1$$48224300_64x8m81_0
timestamp 1755005639
transform 1 0 8149 0 1 10013
box 0 0 1 1
use M2_M1$$48316460_64x8m81  M2_M1$$48316460_64x8m81_0
timestamp 1755005639
transform 1 0 9480 0 1 2532
box 0 0 1 1
use M2_M1$$168351788_64x8m81  M2_M1$$168351788_64x8m81_0
timestamp 1755005639
transform 1 0 5815 0 1 5672
box 0 0 1 1
use M2_M1$$170061868_64x8m81  M2_M1$$170061868_64x8m81_0
timestamp 1755005639
transform 1 0 2811 0 1 4584
box 0 0 1 1
use M2_M1$$170063916_64x8m81  M2_M1$$170063916_64x8m81_0
timestamp 1755005639
transform -1 0 2275 0 1 8014
box 0 0 1 1
use M2_M1$$170064940_64x8m81  M2_M1$$170064940_64x8m81_0
timestamp 1755005639
transform -1 0 2561 0 1 5742
box 0 0 1 1
use M2_M1$$170064940_64x8m81  M2_M1$$170064940_64x8m81_1
timestamp 1755005639
transform -1 0 2561 0 1 6726
box 0 0 1 1
use M2_M1$$199746604_64x8m81  M2_M1$$199746604_64x8m81_0
timestamp 1755005639
transform 1 0 13108 0 1 -612
box 0 0 1 1
use M2_M1$$199746604_64x8m81  M2_M1$$199746604_64x8m81_1
timestamp 1755005639
transform 1 0 10385 0 1 -612
box 0 0 1 1
use M2_M14310589983218_64x8m81  M2_M14310589983218_64x8m81_0
timestamp 1755005639
transform 1 0 8062 0 1 2881
box 0 0 1 1
use M2_M14310589983218_64x8m81  M2_M14310589983218_64x8m81_1
timestamp 1755005639
transform 1 0 8510 0 1 2881
box 0 0 1 1
use M2_M14310589983266_64x8m81  M2_M14310589983266_64x8m81_0
timestamp 1755005639
transform 1 0 5060 0 1 2506
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_0
timestamp 1755005639
transform -1 0 5226 0 1 5491
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_1
timestamp 1755005639
transform 1 0 6412 0 1 5835
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_2
timestamp 1755005639
transform 1 0 11569 0 1 9082
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_3
timestamp 1755005639
transform 1 0 11121 0 1 9082
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_4
timestamp 1755005639
transform 1 0 10670 0 1 9082
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_5
timestamp 1755005639
transform 1 0 7144 0 1 8018
box 0 0 1 1
use M3_M2$$43368492_R270_64x8m81  M3_M2$$43368492_R270_64x8m81_0
timestamp 1755005639
transform 0 -1 5543 -1 0 8499
box 0 0 1 1
use M3_M2$$43368492_R270_64x8m81  M3_M2$$43368492_R270_64x8m81_1
timestamp 1755005639
transform 0 -1 7857 -1 0 8499
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_0
timestamp 1755005639
transform 1 0 12765 0 1 4486
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_1
timestamp 1755005639
transform 1 0 5811 0 1 7368
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_2
timestamp 1755005639
transform 1 0 -149 0 1 7368
box 0 0 1 1
use M3_M2$$43371564_64x8m81  M3_M2$$43371564_64x8m81_3
timestamp 1755005639
transform 1 0 4781 0 1 8732
box 0 0 1 1
use M3_M2$$45008940_64x8m81  M3_M2$$45008940_64x8m81_0
timestamp 1755005639
transform 1 0 6718 0 1 9082
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_0
timestamp 1755005639
transform 1 0 6412 0 1 6613
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_1
timestamp 1755005639
transform -1 0 5002 0 1 6821
box 0 0 1 1
use M3_M2$$47115308_64x8m81  M3_M2$$47115308_64x8m81_0
timestamp 1755005639
transform 1 0 9113 0 1 4348
box 0 0 1 1
use M3_M2$$47332396_64x8m81  M3_M2$$47332396_64x8m81_0
timestamp 1755005639
transform 1 0 6340 0 1 10614
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_0
timestamp 1755005639
transform 1 0 12471 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_1
timestamp 1755005639
transform 1 0 12023 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_2
timestamp 1755005639
transform 1 0 11575 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_3
timestamp 1755005639
transform 1 0 12919 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_4
timestamp 1755005639
transform 1 0 13365 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_5
timestamp 1755005639
transform 1 0 13666 0 1 10274
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_6
timestamp 1755005639
transform 1 0 11127 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_7
timestamp 1755005639
transform 1 0 10679 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_8
timestamp 1755005639
transform 1 0 7543 0 1 9909
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_9
timestamp 1755005639
transform 1 0 8887 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_10
timestamp 1755005639
transform 1 0 9335 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_11
timestamp 1755005639
transform 1 0 9783 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_12
timestamp 1755005639
transform 1 0 7096 0 1 9909
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_13
timestamp 1755005639
transform 1 0 10231 0 1 10240
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_14
timestamp 1755005639
transform 1 0 7144 0 1 6722
box 0 0 1 1
use M3_M2$$47644716_64x8m81  M3_M2$$47644716_64x8m81_0
timestamp 1755005639
transform 1 0 12179 0 1 7395
box 0 0 1 1
use M3_M2$$47644716_64x8m81  M3_M2$$47644716_64x8m81_1
timestamp 1755005639
transform 1 0 12627 0 1 7395
box 0 0 1 1
use M3_M2$$47644716_64x8m81  M3_M2$$47644716_64x8m81_2
timestamp 1755005639
transform 1 0 9922 0 1 7390
box 0 0 1 1
use M3_M2$$47644716_64x8m81  M3_M2$$47644716_64x8m81_3
timestamp 1755005639
transform 1 0 9474 0 1 7390
box 0 0 1 1
use M3_M2$$47644716_64x8m81  M3_M2$$47644716_64x8m81_4
timestamp 1755005639
transform 1 0 11345 0 1 7381
box 0 0 1 1
use M3_M2$$47644716_64x8m81  M3_M2$$47644716_64x8m81_5
timestamp 1755005639
transform 1 0 10897 0 1 7381
box 0 0 1 1
use M3_M2$$47644716_64x8m81  M3_M2$$47644716_64x8m81_6
timestamp 1755005639
transform 1 0 13426 0 1 7395
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_0
timestamp 1755005639
transform 1 0 6355 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_1
timestamp 1755005639
transform 1 0 8147 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_2
timestamp 1755005639
transform 1 0 9781 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_3
timestamp 1755005639
transform 1 0 9333 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_4
timestamp 1755005639
transform 1 0 8885 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_5
timestamp 1755005639
transform 1 0 8595 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_6
timestamp 1755005639
transform 1 0 6803 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_7
timestamp 1755005639
transform 1 0 7251 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_8
timestamp 1755005639
transform 1 0 7699 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_9
timestamp 1755005639
transform 1 0 10677 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_10
timestamp 1755005639
transform 1 0 13365 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_11
timestamp 1755005639
transform 1 0 12917 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_12
timestamp 1755005639
transform 1 0 12469 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_13
timestamp 1755005639
transform 1 0 12021 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_14
timestamp 1755005639
transform 1 0 11573 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_15
timestamp 1755005639
transform 1 0 11125 0 1 15450
box 0 0 1 1
use M3_M2$$47645740_64x8m81  M3_M2$$47645740_64x8m81_16
timestamp 1755005639
transform 1 0 10229 0 1 15450
box 0 0 1 1
use M3_M2$$48066604_64x8m81  M3_M2$$48066604_64x8m81_0
timestamp 1755005639
transform 1 0 12508 0 1 8975
box 0 0 1 1
use M3_M2$$48227372_64x8m81  M3_M2$$48227372_64x8m81_0
timestamp 1755005639
transform 1 0 9480 0 1 2532
box 0 0 1 1
use M3_M2$$48228396_64x8m81  M3_M2$$48228396_64x8m81_0
timestamp 1755005639
transform 1 0 9109 0 1 7390
box 0 0 1 1
use M3_M2$$48229420_64x8m81  M3_M2$$48229420_64x8m81_0
timestamp 1755005639
transform 1 0 11569 0 1 2115
box 0 0 1 1
use M3_M2$$48229420_64x8m81  M3_M2$$48229420_64x8m81_1
timestamp 1755005639
transform 1 0 11957 0 1 2115
box 0 0 1 1
use M3_M2$$48229420_64x8m81  M3_M2$$48229420_64x8m81_2
timestamp 1755005639
transform 1 0 12853 0 1 2115
box 0 0 1 1
use M3_M2$$48229420_64x8m81  M3_M2$$48229420_64x8m81_3
timestamp 1755005639
transform 1 0 10673 0 1 2115
box 0 0 1 1
use M3_M2$$48229420_64x8m81  M3_M2$$48229420_64x8m81_4
timestamp 1755005639
transform 1 0 13541 0 1 2115
box 0 0 1 1
use M3_M2$$48231468_64x8m81  M3_M2$$48231468_64x8m81_0
timestamp 1755005639
transform 1 0 8149 0 1 10013
box 0 0 1 1
use M3_M2$$169753644_64x8m81  M3_M2$$169753644_64x8m81_0
timestamp 1755005639
transform 1 0 2811 0 1 4584
box 0 0 1 1
use M3_M2$$169755692_64x8m81  M3_M2$$169755692_64x8m81_0
timestamp 1755005639
transform -1 0 2275 0 1 8014
box 0 0 1 1
use M3_M2$$169756716_64x8m81  M3_M2$$169756716_64x8m81_0
timestamp 1755005639
transform -1 0 2561 0 1 6726
box 0 0 1 1
use M3_M2$$169756716_64x8m81  M3_M2$$169756716_64x8m81_1
timestamp 1755005639
transform -1 0 2561 0 1 5742
box 0 0 1 1
use M3_M2$$201255980_64x8m81  M3_M2$$201255980_64x8m81_0
timestamp 1755005639
transform 1 0 -213 0 1 -2074
box 0 0 1 1
use M3_M24310589983265_64x8m81  M3_M24310589983265_64x8m81_0
timestamp 1755005639
transform 1 0 5060 0 1 2506
box 0 0 1 1
use M3_M24310589983267_64x8m81  M3_M24310589983267_64x8m81_0
timestamp 1755005639
transform 1 0 8062 0 1 2881
box 0 0 1 1
use M3_M24310589983267_64x8m81  M3_M24310589983267_64x8m81_1
timestamp 1755005639
transform 1 0 8510 0 1 2881
box 0 0 1 1
use nmos_1p2$$46551084_64x8m81  nmos_1p2$$46551084_64x8m81_0
timestamp 1755005639
transform 1 0 7517 0 1 5402
box -31 0 -30 1
use nmos_1p2$$46563372_64x8m81  nmos_1p2$$46563372_64x8m81_0
timestamp 1755005639
transform 1 0 5086 0 1 7941
box -31 0 -30 1
use nmos_1p2$$46563372_64x8m81  nmos_1p2$$46563372_64x8m81_1
timestamp 1755005639
transform 1 0 7003 0 -1 8213
box -31 0 -30 1
use nmos_1p2$$46563372_64x8m81  nmos_1p2$$46563372_64x8m81_2
timestamp 1755005639
transform 1 0 7517 0 -1 8213
box -31 0 -30 1
use nmos_1p2$$47342636_64x8m81  nmos_1p2$$47342636_64x8m81_0
timestamp 1755005639
transform 1 0 5310 0 1 5402
box -31 0 -30 1
use nmos_1p2$$47342636_64x8m81  nmos_1p2$$47342636_64x8m81_1
timestamp 1755005639
transform 1 0 5086 0 1 5402
box -31 0 -30 1
use nmos_1p2$$48302124_64x8m81  nmos_1p2$$48302124_64x8m81_0
timestamp 1755005639
transform 1 0 8145 0 -1 4393
box -31 0 -30 1
use nmos_1p2$$48306220_64x8m81  nmos_1p2$$48306220_64x8m81_0
timestamp 1755005639
transform 1 0 6731 0 1 9039
box -31 0 -30 1
use nmos_1p2$$48308268_64x8m81  nmos_1p2$$48308268_64x8m81_0
timestamp 1755005639
transform 1 0 8968 0 1 9839
box -31 0 -30 1
use nmos_1p2$$48629804_64x8m81  nmos_1p2$$48629804_64x8m81_0
timestamp 1755005639
transform 1 0 6779 0 1 5402
box -31 0 -30 1
use nmos_5p04310589983293_64x8m81  nmos_5p04310589983293_64x8m81_0
timestamp 1755005639
transform 1 0 5157 0 -1 3892
box 0 0 1 1
use nmos_5p04310589983293_64x8m81  nmos_5p04310589983293_64x8m81_1
timestamp 1755005639
transform 1 0 6235 0 -1 3892
box 0 0 1 1
use nmos_5p04310589983297_64x8m81  nmos_5p04310589983297_64x8m81_0
timestamp 1755005639
transform 1 0 7600 0 -1 3940
box 0 0 1 1
use nmos_5p04310589983298_64x8m81  nmos_5p04310589983298_64x8m81_0
timestamp 1755005639
transform 1 0 6954 0 -1 3897
box 0 0 1 1
use pmos_1p2$$46273580_64x8m81  pmos_1p2$$46273580_64x8m81_0
timestamp 1755005639
transform 1 0 6779 0 -1 7742
box -31 0 -30 1
use pmos_1p2$$46285868_64x8m81  pmos_1p2$$46285868_64x8m81_0
timestamp 1755005639
transform 1 0 5086 0 1 7195
box -31 0 -30 1
use pmos_1p2$$46285868_64x8m81  pmos_1p2$$46285868_64x8m81_1
timestamp 1755005639
transform 1 0 7517 0 1 6377
box -31 0 -30 1
use pmos_1p2$$47330348_64x8m81  pmos_1p2$$47330348_64x8m81_0
timestamp 1755005639
transform 1 0 7517 0 -1 7742
box -31 0 -30 1
use pmos_1p2$$47815724_64x8m81  pmos_1p2$$47815724_64x8m81_0
timestamp 1755005639
transform 1 0 12489 0 1 4659
box -31 0 -30 1
use pmos_1p2$$47815724_64x8m81  pmos_1p2$$47815724_64x8m81_1
timestamp 1755005639
transform 1 0 12713 0 1 4659
box -31 0 -30 1
use pmos_1p2$$47815724_64x8m81  pmos_1p2$$47815724_64x8m81_2
timestamp 1755005639
transform 1 0 12265 0 1 4659
box -31 0 -30 1
use pmos_1p2$$47815724_64x8m81  pmos_1p2$$47815724_64x8m81_3
timestamp 1755005639
transform 1 0 12041 0 1 4659
box -31 0 -30 1
use pmos_1p2$$47815724_64x8m81  pmos_1p2$$47815724_64x8m81_4
timestamp 1755005639
transform 1 0 11428 0 1 4659
box -31 0 -30 1
use pmos_1p2$$47815724_64x8m81  pmos_1p2$$47815724_64x8m81_5
timestamp 1755005639
transform 1 0 10980 0 1 4659
box -31 0 -30 1
use pmos_1p2$$47815724_64x8m81  pmos_1p2$$47815724_64x8m81_6
timestamp 1755005639
transform 1 0 10756 0 1 4659
box -31 0 -30 1
use pmos_1p2$$47815724_64x8m81  pmos_1p2$$47815724_64x8m81_7
timestamp 1755005639
transform 1 0 11204 0 1 4659
box -31 0 -30 1
use pmos_1p2$$48623660_64x8m81  pmos_1p2$$48623660_64x8m81_0
timestamp 1755005639
transform 1 0 8145 0 -1 3260
box -31 0 -30 1
use pmos_1p2$$48624684_64x8m81  pmos_1p2$$48624684_64x8m81_0
timestamp 1755005639
transform 1 0 10005 0 1 5293
box -31 0 -30 1
use pmos_1p2$$48624684_64x8m81  pmos_1p2$$48624684_64x8m81_1
timestamp 1755005639
transform 1 0 9557 0 1 5293
box -31 0 -30 1
use pmos_1p2$$48624684_64x8m81  pmos_1p2$$48624684_64x8m81_2
timestamp 1755005639
transform 1 0 9781 0 1 5293
box -31 0 -30 1
use pmos_5p04310589983251_64x8m81  pmos_5p04310589983251_64x8m81_0
timestamp 1755005639
transform 1 0 6748 0 1 6137
box 0 0 1 1
use pmos_5p04310589983278_64x8m81  pmos_5p04310589983278_64x8m81_0
timestamp 1755005639
transform 1 0 5157 0 -1 3260
box 0 0 1 1
use pmos_5p04310589983278_64x8m81  pmos_5p04310589983278_64x8m81_1
timestamp 1755005639
transform 1 0 6235 0 -1 3260
box 0 0 1 1
use pmos_5p04310589983287_64x8m81  pmos_5p04310589983287_64x8m81_0
timestamp 1755005639
transform 1 0 7600 0 -1 3260
box 0 0 1 1
use pmos_5p04310589983292_64x8m81  pmos_5p04310589983292_64x8m81_0
timestamp 1755005639
transform 1 0 6408 0 1 13461
box 0 0 1 1
use pmos_5p04310589983295_64x8m81  pmos_5p04310589983295_64x8m81_0
timestamp 1755005639
transform 1 0 6954 0 -1 3260
box 0 0 1 1
use pmos_5p04310589983296_64x8m81  pmos_5p04310589983296_64x8m81_0
timestamp 1755005639
transform 1 0 8937 0 1 12283
box 0 0 1 1
use wen_v2_64x8m81  wen_v2_64x8m81_0
timestamp 1755005639
transform 1 0 -16 0 1 -2104
box -27 -266 7407 3658
<< labels >>
flabel metal1 s 529 -493 529 -493 0 FreeSans 1000 0 0 0 WEN
port 1 nsew
flabel metal1 s 6616 1004 6616 1004 0 FreeSans 1000 0 0 0 GWE
port 2 nsew
flabel metal3 s 847 5774 847 5774 0 FreeSans 1000 0 0 0 VSS
port 3 nsew
flabel metal3 s 320 4011 320 4011 0 FreeSans 1000 0 0 0 VSS
port 3 nsew
flabel metal3 s 429 6678 429 6678 0 FreeSans 1000 0 0 0 VDD
port 4 nsew
flabel metal3 s 847 8050 847 8050 0 FreeSans 1000 0 0 0 VSS
port 3 nsew
flabel metal3 s -445 -1708 -445 -1708 0 FreeSans 1000 0 0 0 VSS
port 3 nsew
rlabel metal3 s 12652 4305 12652 4305 4 tblhl
port 5 nsew
flabel metal3 s 6414 10067 6414 10067 0 FreeSans 1000 0 0 0 VSS
port 3 nsew
flabel metal3 s -445 -1060 -445 -1060 0 FreeSans 1000 0 0 0 VDD
port 4 nsew
flabel metal3 s -445 -26 -445 -26 0 FreeSans 1000 0 0 0 VDD
port 4 nsew
flabel metal3 s 344 2456 344 2456 0 FreeSans 1000 0 0 0 VDD
port 4 nsew
flabel metal3 s 6414 15414 6414 15414 0 FreeSans 1000 0 0 0 VDD
port 4 nsew
flabel metal3 s -445 1250 -445 1250 0 FreeSans 1000 0 0 0 VSS
port 3 nsew
rlabel metal2 s 8753 -181 8753 -181 4 cen
port 6 nsew
rlabel metal2 s -215 7409 -215 7409 4 clk
port 7 nsew
rlabel metal2 s 12456 13280 12456 13280 4 men
port 8 nsew
<< properties >>
string GDS_END 1305342
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1258880
string path 25.525 19.160 25.525 21.230 
<< end >>
