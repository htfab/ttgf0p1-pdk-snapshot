magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
use nmos_5p04310589983269_64x8m81  nmos_5p04310589983269_64x8m81_0
timestamp 1755005639
transform 1 0 -31 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 78474
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 78224
<< end >>
