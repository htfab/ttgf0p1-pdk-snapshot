magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 770 1486
<< nmos >>
rect 120 209 176 385
rect 280 209 336 385
rect 440 209 496 385
<< pmos >>
rect 120 1015 176 1191
rect 280 1015 336 1191
rect 440 1015 496 1191
<< ndiff >>
rect 32 268 120 385
rect 32 222 45 268
rect 91 222 120 268
rect 32 209 120 222
rect 176 209 280 385
rect 336 209 440 385
rect 496 371 584 385
rect 496 325 525 371
rect 571 325 584 371
rect 496 209 584 325
<< pdiff >>
rect 32 1178 120 1191
rect 32 1132 45 1178
rect 91 1132 120 1178
rect 32 1015 120 1132
rect 176 1075 280 1191
rect 176 1029 205 1075
rect 251 1029 280 1075
rect 176 1015 280 1029
rect 336 1178 440 1191
rect 336 1132 365 1178
rect 411 1132 440 1178
rect 336 1015 440 1132
rect 496 1075 584 1191
rect 496 1029 525 1075
rect 571 1029 584 1075
rect 496 1015 584 1029
<< ndiffc >>
rect 45 222 91 268
rect 525 325 571 371
<< pdiffc >>
rect 45 1132 91 1178
rect 205 1029 251 1075
rect 365 1132 411 1178
rect 525 1029 571 1075
<< psubdiff >>
rect 28 87 656 100
rect 28 41 69 87
rect 615 41 656 87
rect 28 28 656 41
<< nsubdiff >>
rect 28 1359 656 1372
rect 28 1313 69 1359
rect 615 1313 656 1359
rect 28 1300 656 1313
<< psubdiffcont >>
rect 69 41 615 87
<< nsubdiffcont >>
rect 69 1313 615 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 120 716 176 1015
rect 280 716 336 1015
rect 440 716 496 1015
rect 32 703 176 716
rect 32 657 45 703
rect 91 657 176 703
rect 32 644 176 657
rect 224 703 336 716
rect 224 657 237 703
rect 283 657 336 703
rect 224 644 336 657
rect 384 703 496 716
rect 384 657 397 703
rect 443 657 496 703
rect 384 644 496 657
rect 120 385 176 644
rect 280 385 336 644
rect 440 385 496 644
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
<< polycontact >>
rect 45 657 91 703
rect 237 657 283 703
rect 397 657 443 703
<< metal1 >>
rect 0 1359 684 1400
rect 0 1313 69 1359
rect 615 1313 684 1359
rect 0 1178 684 1313
rect 0 1132 45 1178
rect 91 1132 365 1178
rect 411 1132 684 1178
rect 42 703 94 1086
rect 205 1075 574 1086
rect 251 1029 525 1075
rect 571 1029 574 1075
rect 205 1018 574 1029
rect 42 657 45 703
rect 91 657 94 703
rect 42 314 94 657
rect 234 703 286 972
rect 234 657 237 703
rect 283 657 286 703
rect 234 314 286 657
rect 394 703 446 972
rect 394 657 397 703
rect 443 657 446 703
rect 394 314 446 657
rect 522 371 574 1018
rect 522 325 525 371
rect 571 325 574 371
rect 522 314 574 325
rect 0 222 45 268
rect 91 222 684 268
rect 0 87 684 222
rect 0 41 69 87
rect 615 41 684 87
rect 0 0 684 41
<< labels >>
rlabel metal1 s 0 0 684 268 4 vss
port 3 nsew
rlabel metal1 s 0 1132 684 1400 4 vdd
port 5 nsew
rlabel metal1 s 42 314 94 1086 4 i0
port 7 nsew
rlabel metal1 s 522 314 574 1086 4 nq
port 9 nsew
rlabel metal1 s 234 314 286 972 4 i1
port 11 nsew
rlabel metal1 s 394 314 446 972 4 i2
port 13 nsew
<< end >>
