magic
tech gf180mcuD
magscale 1 10
timestamp 1751889808
<< nwell >>
rect -86 354 870 870
<< pwell >>
rect -86 -86 870 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
<< ndiff >>
rect 28 127 116 268
rect 28 81 41 127
rect 87 81 116 127
rect 28 68 116 81
rect 172 230 276 268
rect 172 184 201 230
rect 247 184 276 230
rect 172 68 276 184
rect 332 127 436 268
rect 332 81 361 127
rect 407 81 436 127
rect 332 68 436 81
rect 492 251 596 268
rect 492 205 521 251
rect 567 205 596 251
rect 492 68 596 205
rect 652 255 756 268
rect 652 81 681 255
rect 727 81 756 255
rect 652 68 756 81
<< pdiff >>
rect 28 585 116 716
rect 28 539 41 585
rect 87 539 116 585
rect 28 440 116 539
rect 172 440 276 716
rect 332 703 436 716
rect 332 657 361 703
rect 407 657 436 703
rect 332 440 436 657
rect 492 667 596 716
rect 492 453 521 667
rect 567 453 596 667
rect 492 440 596 453
rect 652 703 756 716
rect 652 453 681 703
rect 727 453 756 703
rect 652 440 756 453
<< ndiffc >>
rect 41 81 87 127
rect 201 184 247 230
rect 361 81 407 127
rect 521 205 567 251
rect 681 81 727 255
<< pdiffc >>
rect 41 539 87 585
rect 361 657 407 703
rect 521 453 567 667
rect 681 453 727 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 116 397 172 440
rect 91 379 172 397
rect 276 396 332 440
rect 436 396 492 440
rect 91 333 104 379
rect 150 333 172 379
rect 91 312 172 333
rect 116 268 172 312
rect 251 377 332 396
rect 251 331 271 377
rect 317 331 332 377
rect 251 311 332 331
rect 380 377 492 396
rect 380 331 393 377
rect 439 373 492 377
rect 596 373 652 440
rect 439 331 652 373
rect 380 330 652 331
rect 380 311 492 330
rect 276 268 332 311
rect 436 268 492 311
rect 596 268 652 330
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
<< polycontact >>
rect 104 333 150 379
rect 271 331 317 377
rect 393 331 439 377
<< metal1 >>
rect 0 724 784 844
rect 361 703 407 724
rect 681 703 727 724
rect 361 646 407 657
rect 521 667 607 678
rect 41 585 424 600
rect 87 554 424 585
rect 41 528 87 539
rect 41 379 172 397
rect 41 333 104 379
rect 150 333 172 379
rect 41 312 172 333
rect 251 377 332 508
rect 251 331 271 377
rect 317 331 332 377
rect 251 311 332 331
rect 378 396 424 554
rect 567 453 607 667
rect 378 377 439 396
rect 378 331 393 377
rect 378 311 439 331
rect 378 230 424 311
rect 188 184 201 230
rect 247 184 424 230
rect 521 251 607 453
rect 681 430 727 453
rect 567 205 607 251
rect 521 184 607 205
rect 681 255 727 290
rect 41 127 87 138
rect 41 60 87 81
rect 361 127 407 138
rect 361 60 407 81
rect 681 60 727 81
rect 0 -60 784 60
<< labels >>
flabel metal1 s 0 724 784 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 784 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 251 311 332 508 0 FreeSans 200 0 0 0 B
port 5 nsew signal input
flabel metal1 41 312 172 397 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 521 184 607 678 0 FreeSans 200 0 0 0 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 784 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
