magic
tech gf180mcuD
magscale 1 10
timestamp 1751633659
<< nwell >>
rect -86 354 870 870
<< pwell >>
rect -86 -86 870 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
<< ndiff >>
rect 28 223 116 268
rect 28 81 41 223
rect 87 81 116 223
rect 28 68 116 81
rect 172 255 276 268
rect 172 209 201 255
rect 247 209 276 255
rect 172 68 276 209
rect 332 236 436 268
rect 332 81 361 236
rect 407 81 436 236
rect 332 68 436 81
rect 492 255 596 268
rect 492 209 521 255
rect 567 209 596 255
rect 492 68 596 209
rect 652 255 756 268
rect 652 81 681 255
rect 727 81 756 255
rect 652 68 756 81
<< pdiff >>
rect 28 703 116 716
rect 28 482 41 703
rect 87 482 116 703
rect 28 440 116 482
rect 172 666 276 716
rect 172 453 201 666
rect 247 453 276 666
rect 172 440 276 453
rect 332 703 436 716
rect 332 470 361 703
rect 407 470 436 703
rect 332 440 436 470
rect 492 666 596 716
rect 492 453 521 666
rect 567 453 596 666
rect 492 440 596 453
rect 652 703 756 716
rect 652 453 681 703
rect 727 453 756 703
rect 652 440 756 453
<< ndiffc >>
rect 41 81 87 223
rect 201 209 247 255
rect 361 81 407 236
rect 521 209 567 255
rect 681 81 727 255
<< pdiffc >>
rect 41 482 87 703
rect 201 453 247 666
rect 361 470 407 703
rect 521 453 567 666
rect 681 453 727 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 116 398 172 440
rect 96 387 172 398
rect 276 398 332 440
rect 436 420 492 440
rect 596 420 652 440
rect 436 398 652 420
rect 276 387 652 398
rect 96 384 652 387
rect 96 338 109 384
rect 155 358 652 384
rect 155 338 492 358
rect 96 336 492 338
rect 96 325 332 336
rect 116 268 172 325
rect 276 268 332 325
rect 436 268 492 336
rect 596 268 652 358
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
<< polycontact >>
rect 109 338 155 384
<< metal1 >>
rect 0 724 784 844
rect 41 703 87 724
rect 361 703 407 724
rect 41 471 87 482
rect 201 666 247 677
rect 681 703 727 724
rect 361 459 407 470
rect 521 666 567 677
rect 201 451 247 453
rect 41 384 155 425
rect 41 338 109 384
rect 41 318 155 338
rect 201 387 270 451
rect 521 387 567 453
rect 681 435 727 453
rect 201 341 567 387
rect 201 255 270 341
rect 41 223 87 247
rect 247 252 270 255
rect 521 255 567 341
rect 201 198 247 209
rect 361 236 407 247
rect 41 60 87 81
rect 521 198 567 209
rect 681 255 727 279
rect 361 60 407 81
rect 681 60 727 81
rect 0 -60 784 60
<< labels >>
flabel metal1 s 0 724 784 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 784 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 201 252 270 451 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 41 318 155 425 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 784 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
