magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 352 982 870
<< pwell >>
rect -86 -86 982 352
<< metal1 >>
rect 0 724 896 844
rect 49 645 95 724
rect 132 308 204 562
rect 356 308 428 674
rect 521 506 567 724
rect 501 60 547 153
rect 690 111 774 676
rect 0 -60 896 60
<< obsm1 >>
rect 253 258 299 665
rect 589 258 635 397
rect 49 211 635 258
rect 49 161 95 211
<< labels >>
rlabel metal1 s 132 308 204 562 6 A1
port 1 nsew default input
rlabel metal1 s 356 308 428 674 6 A2
port 2 nsew default input
rlabel metal1 s 690 111 774 676 6 Z
port 3 nsew default output
rlabel metal1 s 521 506 567 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 49 645 95 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 724 896 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel nwell s -86 352 982 870 6 VNW
port 5 nsew power bidirectional
rlabel pwell s -86 -86 982 352 6 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 0 -60 896 60 8 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 501 60 547 153 6 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 896 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1211902
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1208972
<< end >>
