magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 407 5238 870
rect -86 352 575 407
rect 943 352 5238 407
<< pwell >>
rect 575 352 943 407
rect -86 -86 5238 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 1064 68 1184 232
rect 1288 68 1408 232
rect 1512 68 1632 232
rect 1736 68 1856 232
rect 1960 68 2080 232
rect 2184 68 2304 232
rect 2408 68 2528 232
rect 2632 68 2752 232
rect 2856 68 2976 232
rect 3080 68 3200 232
rect 3304 68 3424 232
rect 3528 68 3648 232
rect 3752 68 3872 232
rect 3976 68 4096 232
rect 4200 68 4320 232
rect 4424 68 4544 232
rect 4648 68 4768 232
rect 4872 68 4992 232
<< mvpmos >>
rect 172 527 272 716
rect 376 527 476 716
rect 660 527 760 716
rect 1184 481 1284 716
rect 1388 481 1488 716
rect 1592 481 1692 716
rect 1796 481 1896 716
rect 2000 481 2100 716
rect 2204 481 2304 716
rect 2408 481 2508 716
rect 2612 481 2712 716
rect 2816 481 2916 716
rect 3020 481 3120 716
rect 3224 481 3324 716
rect 3428 481 3528 716
rect 3632 481 3732 716
rect 3836 481 3936 716
rect 4040 481 4140 716
rect 4244 481 4344 716
rect 4448 481 4548 716
rect 4652 481 4752 716
<< mvndiff >>
rect 752 274 824 287
rect 752 232 765 274
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 68 124 173
rect 244 128 348 232
rect 244 82 273 128
rect 319 82 348 128
rect 244 68 348 82
rect 468 169 572 232
rect 468 123 497 169
rect 543 123 572 169
rect 468 68 572 123
rect 692 228 765 232
rect 811 228 824 274
rect 692 68 824 228
rect 932 95 1064 232
rect 932 49 945 95
rect 991 68 1064 95
rect 1184 219 1288 232
rect 1184 173 1213 219
rect 1259 173 1288 219
rect 1184 68 1288 173
rect 1408 127 1512 232
rect 1408 81 1437 127
rect 1483 81 1512 127
rect 1408 68 1512 81
rect 1632 219 1736 232
rect 1632 173 1661 219
rect 1707 173 1736 219
rect 1632 68 1736 173
rect 1856 127 1960 232
rect 1856 81 1885 127
rect 1931 81 1960 127
rect 1856 68 1960 81
rect 2080 219 2184 232
rect 2080 173 2109 219
rect 2155 173 2184 219
rect 2080 68 2184 173
rect 2304 127 2408 232
rect 2304 81 2333 127
rect 2379 81 2408 127
rect 2304 68 2408 81
rect 2528 219 2632 232
rect 2528 173 2557 219
rect 2603 173 2632 219
rect 2528 68 2632 173
rect 2752 127 2856 232
rect 2752 81 2781 127
rect 2827 81 2856 127
rect 2752 68 2856 81
rect 2976 219 3080 232
rect 2976 173 3005 219
rect 3051 173 3080 219
rect 2976 68 3080 173
rect 3200 127 3304 232
rect 3200 81 3229 127
rect 3275 81 3304 127
rect 3200 68 3304 81
rect 3424 219 3528 232
rect 3424 173 3453 219
rect 3499 173 3528 219
rect 3424 68 3528 173
rect 3648 127 3752 232
rect 3648 81 3677 127
rect 3723 81 3752 127
rect 3648 68 3752 81
rect 3872 219 3976 232
rect 3872 173 3901 219
rect 3947 173 3976 219
rect 3872 68 3976 173
rect 4096 127 4200 232
rect 4096 81 4125 127
rect 4171 81 4200 127
rect 4096 68 4200 81
rect 4320 219 4424 232
rect 4320 173 4349 219
rect 4395 173 4424 219
rect 4320 68 4424 173
rect 4544 127 4648 232
rect 4544 81 4573 127
rect 4619 81 4648 127
rect 4544 68 4648 81
rect 4768 219 4872 232
rect 4768 173 4797 219
rect 4843 173 4872 219
rect 4768 68 4872 173
rect 4992 127 5080 232
rect 4992 81 5021 127
rect 5067 81 5080 127
rect 4992 68 5080 81
rect 991 49 1004 68
rect 932 36 1004 49
<< mvpdiff >>
rect 84 602 172 716
rect 84 556 97 602
rect 143 556 172 602
rect 84 527 172 556
rect 272 698 376 716
rect 272 652 301 698
rect 347 652 376 698
rect 272 527 376 652
rect 476 678 660 716
rect 476 632 548 678
rect 594 632 660 678
rect 476 527 660 632
rect 760 586 848 716
rect 760 540 789 586
rect 835 540 848 586
rect 760 527 848 540
rect 1096 665 1184 716
rect 1096 619 1109 665
rect 1155 619 1184 665
rect 1096 481 1184 619
rect 1284 665 1388 716
rect 1284 525 1313 665
rect 1359 525 1388 665
rect 1284 481 1388 525
rect 1488 665 1592 716
rect 1488 619 1517 665
rect 1563 619 1592 665
rect 1488 481 1592 619
rect 1692 665 1796 716
rect 1692 525 1721 665
rect 1767 525 1796 665
rect 1692 481 1796 525
rect 1896 665 2000 716
rect 1896 619 1925 665
rect 1971 619 2000 665
rect 1896 481 2000 619
rect 2100 665 2204 716
rect 2100 525 2129 665
rect 2175 525 2204 665
rect 2100 481 2204 525
rect 2304 665 2408 716
rect 2304 619 2333 665
rect 2379 619 2408 665
rect 2304 481 2408 619
rect 2508 665 2612 716
rect 2508 525 2537 665
rect 2583 525 2612 665
rect 2508 481 2612 525
rect 2712 703 2816 716
rect 2712 657 2741 703
rect 2787 657 2816 703
rect 2712 481 2816 657
rect 2916 665 3020 716
rect 2916 525 2945 665
rect 2991 525 3020 665
rect 2916 481 3020 525
rect 3120 703 3224 716
rect 3120 657 3149 703
rect 3195 657 3224 703
rect 3120 481 3224 657
rect 3324 665 3428 716
rect 3324 525 3353 665
rect 3399 525 3428 665
rect 3324 481 3428 525
rect 3528 703 3632 716
rect 3528 657 3557 703
rect 3603 657 3632 703
rect 3528 481 3632 657
rect 3732 665 3836 716
rect 3732 525 3761 665
rect 3807 525 3836 665
rect 3732 481 3836 525
rect 3936 703 4040 716
rect 3936 657 3965 703
rect 4011 657 4040 703
rect 3936 481 4040 657
rect 4140 665 4244 716
rect 4140 525 4169 665
rect 4215 525 4244 665
rect 4140 481 4244 525
rect 4344 703 4448 716
rect 4344 657 4373 703
rect 4419 657 4448 703
rect 4344 481 4448 657
rect 4548 665 4652 716
rect 4548 525 4577 665
rect 4623 525 4652 665
rect 4548 481 4652 525
rect 4752 665 4840 716
rect 4752 619 4781 665
rect 4827 619 4840 665
rect 4752 481 4840 619
<< mvndiffc >>
rect 49 173 95 219
rect 273 82 319 128
rect 497 123 543 169
rect 765 228 811 274
rect 945 49 991 95
rect 1213 173 1259 219
rect 1437 81 1483 127
rect 1661 173 1707 219
rect 1885 81 1931 127
rect 2109 173 2155 219
rect 2333 81 2379 127
rect 2557 173 2603 219
rect 2781 81 2827 127
rect 3005 173 3051 219
rect 3229 81 3275 127
rect 3453 173 3499 219
rect 3677 81 3723 127
rect 3901 173 3947 219
rect 4125 81 4171 127
rect 4349 173 4395 219
rect 4573 81 4619 127
rect 4797 173 4843 219
rect 5021 81 5067 127
<< mvpdiffc >>
rect 97 556 143 602
rect 301 652 347 698
rect 548 632 594 678
rect 789 540 835 586
rect 1109 619 1155 665
rect 1313 525 1359 665
rect 1517 619 1563 665
rect 1721 525 1767 665
rect 1925 619 1971 665
rect 2129 525 2175 665
rect 2333 619 2379 665
rect 2537 525 2583 665
rect 2741 657 2787 703
rect 2945 525 2991 665
rect 3149 657 3195 703
rect 3353 525 3399 665
rect 3557 657 3603 703
rect 3761 525 3807 665
rect 3965 657 4011 703
rect 4169 525 4215 665
rect 4373 657 4419 703
rect 4577 525 4623 665
rect 4781 619 4827 665
<< polysilicon >>
rect 172 716 272 760
rect 376 716 476 760
rect 660 716 760 760
rect 1184 716 1284 760
rect 1388 716 1488 760
rect 1592 716 1692 760
rect 1796 716 1896 760
rect 2000 716 2100 760
rect 2204 716 2304 760
rect 2408 716 2508 760
rect 2612 716 2712 760
rect 2816 716 2916 760
rect 3020 716 3120 760
rect 3224 716 3324 760
rect 3428 716 3528 760
rect 3632 716 3732 760
rect 3836 716 3936 760
rect 4040 716 4140 760
rect 4244 716 4344 760
rect 4448 716 4548 760
rect 4652 716 4752 760
rect 172 413 272 527
rect 376 413 476 527
rect 660 493 760 527
rect 660 447 673 493
rect 719 447 760 493
rect 660 434 760 447
rect 1184 415 1284 481
rect 124 412 612 413
rect 124 366 185 412
rect 231 373 612 412
rect 1184 399 1211 415
rect 231 366 244 373
rect 124 232 244 366
rect 348 311 468 324
rect 348 265 381 311
rect 427 265 468 311
rect 348 232 468 265
rect 572 288 612 373
rect 1064 369 1211 399
rect 1257 399 1284 415
rect 1388 415 1488 481
rect 1388 399 1415 415
rect 1257 369 1415 399
rect 1461 399 1488 415
rect 1592 415 1692 481
rect 1592 399 1619 415
rect 1461 369 1619 399
rect 1665 399 1692 415
rect 1796 415 1896 481
rect 1796 399 1823 415
rect 1665 369 1823 399
rect 1869 399 1896 415
rect 2000 415 2100 481
rect 2000 399 2027 415
rect 1869 369 2027 399
rect 2073 399 2100 415
rect 2204 415 2304 481
rect 2204 399 2231 415
rect 2073 369 2231 399
rect 2277 369 2304 415
rect 2408 439 2508 481
rect 2408 393 2449 439
rect 2495 420 2508 439
rect 2612 439 2712 481
rect 2612 420 2638 439
rect 2495 393 2638 420
rect 2684 420 2712 439
rect 2816 439 2916 481
rect 2816 420 2843 439
rect 2684 393 2843 420
rect 2889 420 2916 439
rect 3020 439 3120 481
rect 3020 420 3045 439
rect 2889 393 3045 420
rect 3091 420 3120 439
rect 3224 439 3324 481
rect 3224 420 3249 439
rect 3091 393 3249 420
rect 3295 420 3324 439
rect 3428 439 3528 481
rect 3428 420 3441 439
rect 3295 393 3441 420
rect 3487 420 3528 439
rect 3632 420 3732 481
rect 3836 439 3936 481
rect 3836 420 3877 439
rect 3487 393 3877 420
rect 3923 420 3936 439
rect 4040 439 4140 481
rect 4040 420 4067 439
rect 3923 393 4067 420
rect 4113 420 4140 439
rect 4244 439 4344 481
rect 4244 420 4271 439
rect 4113 393 4271 420
rect 4317 420 4344 439
rect 4448 439 4548 481
rect 4448 420 4475 439
rect 4317 393 4475 420
rect 4521 420 4548 439
rect 4652 439 4752 481
rect 4652 420 4682 439
rect 4521 393 4682 420
rect 4728 393 4752 439
rect 2408 380 4752 393
rect 1064 349 2304 369
rect 572 232 692 288
rect 1064 232 1184 349
rect 1288 232 1408 349
rect 1512 232 1632 349
rect 1736 232 1856 349
rect 1960 232 2080 349
rect 2184 232 2304 349
rect 2408 319 4992 332
rect 2408 273 2443 319
rect 2489 292 2667 319
rect 2489 273 2528 292
rect 2408 232 2528 273
rect 2632 273 2667 292
rect 2713 292 2892 319
rect 2713 273 2752 292
rect 2632 232 2752 273
rect 2856 273 2892 292
rect 2938 292 3118 319
rect 2938 273 2976 292
rect 2856 232 2976 273
rect 3080 273 3118 292
rect 3164 292 3317 319
rect 3164 273 3200 292
rect 3080 232 3200 273
rect 3304 273 3317 292
rect 3363 292 3813 319
rect 3363 273 3424 292
rect 3304 232 3424 273
rect 3528 232 3648 292
rect 3752 273 3813 292
rect 3859 292 4013 319
rect 3859 273 3872 292
rect 3752 232 3872 273
rect 3976 273 4013 292
rect 4059 292 4236 319
rect 4059 273 4096 292
rect 3976 232 4096 273
rect 4200 273 4236 292
rect 4282 292 4462 319
rect 4282 273 4320 292
rect 4200 232 4320 273
rect 4424 273 4462 292
rect 4508 292 4682 319
rect 4508 273 4544 292
rect 4424 232 4544 273
rect 4648 273 4682 292
rect 4728 292 4992 319
rect 4728 273 4768 292
rect 4648 232 4768 273
rect 4872 232 4992 292
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 1064 24 1184 68
rect 1288 24 1408 68
rect 1512 24 1632 68
rect 1736 24 1856 68
rect 1960 24 2080 68
rect 2184 24 2304 68
rect 2408 24 2528 68
rect 2632 24 2752 68
rect 2856 24 2976 68
rect 3080 24 3200 68
rect 3304 24 3424 68
rect 3528 24 3648 68
rect 3752 24 3872 68
rect 3976 24 4096 68
rect 4200 24 4320 68
rect 4424 24 4544 68
rect 4648 24 4768 68
rect 4872 24 4992 68
<< polycontact >>
rect 673 447 719 493
rect 185 366 231 412
rect 381 265 427 311
rect 1211 369 1257 415
rect 1415 369 1461 415
rect 1619 369 1665 415
rect 1823 369 1869 415
rect 2027 369 2073 415
rect 2231 369 2277 415
rect 2449 393 2495 439
rect 2638 393 2684 439
rect 2843 393 2889 439
rect 3045 393 3091 439
rect 3249 393 3295 439
rect 3441 393 3487 439
rect 3877 393 3923 439
rect 4067 393 4113 439
rect 4271 393 4317 439
rect 4475 393 4521 439
rect 4682 393 4728 439
rect 2443 273 2489 319
rect 2667 273 2713 319
rect 2892 273 2938 319
rect 3118 273 3164 319
rect 3317 273 3363 319
rect 3813 273 3859 319
rect 4013 273 4059 319
rect 4236 273 4282 319
rect 4462 273 4508 319
rect 4682 273 4728 319
<< metal1 >>
rect 0 724 5152 844
rect 290 698 358 724
rect 290 652 301 698
rect 347 652 358 698
rect 537 632 548 678
rect 594 632 965 678
rect 84 556 97 602
rect 143 556 427 602
rect 381 504 427 556
rect 778 540 789 586
rect 835 540 846 586
rect 381 493 730 504
rect 381 447 673 493
rect 719 447 730 493
rect 74 412 318 430
rect 74 366 185 412
rect 231 366 318 412
rect 74 354 318 366
rect 381 311 427 447
rect 778 401 846 540
rect 38 219 427 265
rect 497 355 846 401
rect 919 552 965 632
rect 1098 665 1166 724
rect 1098 619 1109 665
rect 1155 619 1166 665
rect 1098 608 1166 619
rect 1302 665 1370 676
rect 1302 552 1313 665
rect 919 525 1313 552
rect 1359 552 1370 665
rect 1506 665 1574 724
rect 1506 619 1517 665
rect 1563 619 1574 665
rect 1506 608 1574 619
rect 1710 665 1778 676
rect 1710 552 1721 665
rect 1359 525 1721 552
rect 1767 552 1778 665
rect 1914 665 1982 724
rect 1914 619 1925 665
rect 1971 619 1982 665
rect 1914 608 1982 619
rect 2118 665 2186 676
rect 2118 552 2129 665
rect 1767 525 2129 552
rect 2175 552 2186 665
rect 2322 665 2390 724
rect 2730 703 2798 724
rect 2322 619 2333 665
rect 2379 619 2390 665
rect 2322 608 2390 619
rect 2526 665 2594 676
rect 2175 525 2402 552
rect 919 506 2402 525
rect 2526 525 2537 665
rect 2583 594 2594 665
rect 2730 657 2741 703
rect 2787 657 2798 703
rect 3138 703 3206 724
rect 2934 665 3002 676
rect 2934 594 2945 665
rect 2583 525 2945 594
rect 2991 594 3002 665
rect 3138 657 3149 703
rect 3195 657 3206 703
rect 3546 703 3614 724
rect 3342 665 3410 676
rect 3342 594 3353 665
rect 2991 525 3353 594
rect 3399 594 3410 665
rect 3546 657 3557 703
rect 3603 657 3614 703
rect 3954 703 4022 724
rect 3750 665 3818 676
rect 3750 594 3761 665
rect 3399 525 3761 594
rect 3807 594 3818 665
rect 3954 657 3965 703
rect 4011 657 4022 703
rect 4362 703 4430 724
rect 4158 665 4226 676
rect 4158 594 4169 665
rect 3807 525 4169 594
rect 4215 594 4226 665
rect 4362 657 4373 703
rect 4419 657 4430 703
rect 4566 665 4634 676
rect 4566 594 4577 665
rect 4215 525 4577 594
rect 4623 525 4634 665
rect 4770 665 4838 724
rect 4770 619 4781 665
rect 4827 619 4838 665
rect 4770 608 4838 619
rect 2526 506 4634 525
rect 38 173 49 219
rect 95 173 106 219
rect 38 170 106 173
rect 497 169 543 355
rect 919 309 965 506
rect 2356 439 2402 506
rect 1025 415 2296 430
rect 1025 369 1211 415
rect 1257 369 1415 415
rect 1461 369 1619 415
rect 1665 369 1823 415
rect 1869 369 2027 415
rect 2073 369 2231 415
rect 2277 369 2296 415
rect 2356 393 2449 439
rect 2495 393 2638 439
rect 2684 393 2843 439
rect 2889 393 3045 439
rect 3091 393 3249 439
rect 3295 393 3441 439
rect 3487 393 3498 439
rect 1025 354 2296 369
rect 754 274 965 309
rect 754 228 765 274
rect 811 263 965 274
rect 2356 273 2443 319
rect 2489 273 2667 319
rect 2713 273 2892 319
rect 2938 273 3118 319
rect 3164 273 3317 319
rect 3363 273 3375 319
rect 811 228 822 263
rect 2356 219 2402 273
rect 3580 227 3700 506
rect 3866 393 3877 439
rect 3923 393 4067 439
rect 4113 393 4271 439
rect 4317 393 4475 439
rect 4521 393 4682 439
rect 4728 393 4741 439
rect 3802 273 3813 319
rect 3859 273 4013 319
rect 4059 273 4236 319
rect 4282 273 4462 319
rect 4508 273 4682 319
rect 4728 273 4741 319
rect 1139 187 1213 219
rect 262 128 330 131
rect 262 82 273 128
rect 319 82 330 128
rect 843 173 1213 187
rect 1259 173 1661 219
rect 1707 173 2109 219
rect 2155 173 2402 219
rect 2546 219 4854 227
rect 2546 173 2557 219
rect 2603 173 3005 219
rect 3051 173 3453 219
rect 3499 173 3901 219
rect 3947 173 4349 219
rect 4395 173 4797 219
rect 4843 173 4854 219
rect 843 152 1189 173
rect 543 141 1189 152
rect 543 123 888 141
rect 497 106 888 123
rect 262 60 330 82
rect 934 60 945 95
rect 0 49 945 60
rect 991 60 1002 95
rect 1426 81 1437 127
rect 1483 81 1494 127
rect 1426 60 1494 81
rect 1874 81 1885 127
rect 1931 81 1942 127
rect 1874 60 1942 81
rect 2322 81 2333 127
rect 2379 81 2390 127
rect 2322 60 2390 81
rect 2770 81 2781 127
rect 2827 81 2838 127
rect 2770 60 2838 81
rect 3218 81 3229 127
rect 3275 81 3286 127
rect 3218 60 3286 81
rect 3666 81 3677 127
rect 3723 81 3734 127
rect 3666 60 3734 81
rect 4114 81 4125 127
rect 4171 81 4182 127
rect 4114 60 4182 81
rect 4562 81 4573 127
rect 4619 81 4630 127
rect 4562 60 4630 81
rect 5010 81 5021 127
rect 5067 81 5078 127
rect 5010 60 5078 81
rect 991 49 5152 60
rect 0 -60 5152 49
<< labels >>
flabel metal1 s 0 724 5152 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 262 127 330 131 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 1025 354 2296 430 0 FreeSans 400 0 0 0 I
port 2 nsew default input
flabel metal1 s 4566 594 4634 676 0 FreeSans 400 0 0 0 Z
port 3 nsew default output
flabel metal1 s 74 354 318 430 0 FreeSans 600 0 0 0 EN
port 1 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 4158 594 4226 676 1 Z
port 3 nsew default output
rlabel metal1 s 3750 594 3818 676 1 Z
port 3 nsew default output
rlabel metal1 s 3342 594 3410 676 1 Z
port 3 nsew default output
rlabel metal1 s 2934 594 3002 676 1 Z
port 3 nsew default output
rlabel metal1 s 2526 594 2594 676 1 Z
port 3 nsew default output
rlabel metal1 s 2526 506 4634 594 1 Z
port 3 nsew default output
rlabel metal1 s 3580 227 3700 506 1 Z
port 3 nsew default output
rlabel metal1 s 2546 173 4854 227 1 Z
port 3 nsew default output
rlabel metal1 s 4770 657 4838 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4362 657 4430 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3954 657 4022 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3546 657 3614 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3138 657 3206 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2730 657 2798 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2322 657 2390 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1914 657 1982 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1506 657 1574 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1098 657 1166 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 657 358 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4770 652 4838 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2322 652 2390 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1914 652 1982 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1506 652 1574 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1098 652 1166 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 652 358 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4770 608 4838 652 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2322 608 2390 652 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1914 608 1982 652 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1506 608 1574 652 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1098 608 1166 652 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5010 95 5078 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4562 95 4630 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4114 95 4182 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3666 95 3734 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3218 95 3286 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2770 95 2838 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2322 95 2390 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1874 95 1942 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1426 95 1494 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 95 330 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5010 60 5078 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4562 60 4630 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4114 60 4182 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3666 60 3734 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3218 60 3286 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2770 60 2838 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2322 60 2390 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1874 60 1942 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1426 60 1494 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 95 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5152 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5152 784
string GDS_END 1427884
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1417274
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
