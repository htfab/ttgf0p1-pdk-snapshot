magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect 464 29129 5755 29130
rect 322 23868 5755 29129
rect 322 18380 5591 19962
rect 322 17408 5723 18380
rect 322 17407 629 17408
rect 120 15337 750 15918
rect 1464 15337 2094 15670
rect 120 12914 2094 15337
rect 1449 9405 2303 9582
rect 1449 9389 2930 9405
rect 621 9182 2930 9389
rect 100 8392 2930 9182
rect 620 8391 1475 8392
rect 2300 8391 2930 8392
rect 621 8310 1475 8391
rect 2301 7761 2930 8391
rect 3188 2700 3233 2702
<< mvnmos >>
rect 881 22317 1001 23679
rect 1501 22317 1621 23679
rect 2120 22317 2240 23679
rect 2740 22317 2860 23679
rect 3358 22317 3478 23679
rect 3978 22317 4098 23679
rect 4597 22317 4717 23679
rect 5217 22317 5337 23679
rect 881 20313 1001 21675
rect 1501 20313 1621 21675
rect 2120 20313 2240 21675
rect 2740 20313 2860 21675
rect 3358 20313 3478 21675
rect 3978 20313 4098 21675
rect 4597 20313 4717 21675
rect 5217 20313 5337 21675
rect 855 17143 975 17257
rect 1079 17143 1199 17257
rect 1303 17143 1423 17257
rect 1527 17143 1647 17257
rect 2094 17143 2214 17257
rect 2318 17143 2438 17257
rect 2542 17143 2662 17257
rect 2766 17143 2886 17257
rect 3332 17143 3452 17257
rect 3556 17143 3676 17257
rect 3780 17143 3900 17257
rect 4004 17143 4124 17257
rect 4571 17143 4691 17257
rect 4795 17143 4915 17257
rect 5019 17143 5139 17257
rect 5243 17143 5363 17257
rect 1043 15476 1163 15704
rect 375 9898 495 12620
rect 823 10351 943 12619
rect 1271 10351 1391 12619
rect 1719 10351 1839 12619
rect 986 9619 1106 9811
rect 1704 9719 1824 9911
rect 2556 9543 2676 9997
rect 876 7978 996 8170
rect 1100 7978 1220 8170
rect 1704 7957 1824 8149
rect 1928 7957 2048 8149
<< mvpmos >>
rect 769 27951 889 28633
rect 993 27951 1113 28633
rect 1389 27951 1509 28633
rect 1613 27951 1733 28633
rect 2008 27951 2128 28633
rect 2232 27951 2352 28633
rect 2628 27951 2748 28633
rect 2852 27951 2972 28633
rect 3246 27951 3366 28633
rect 3470 27951 3590 28633
rect 3866 27951 3986 28633
rect 4090 27951 4210 28633
rect 4485 27951 4605 28633
rect 4709 27951 4829 28633
rect 5069 27951 5189 28633
rect 5294 27951 5414 28633
rect 769 27176 889 27858
rect 993 27176 1113 27858
rect 1389 27176 1509 27858
rect 1613 27176 1733 27858
rect 2008 27176 2128 27858
rect 2232 27176 2352 27858
rect 2628 27176 2748 27858
rect 2852 27176 2972 27858
rect 3246 27176 3366 27858
rect 3470 27176 3590 27858
rect 3866 27176 3986 27858
rect 4090 27176 4210 27858
rect 4485 27176 4605 27858
rect 4709 27176 4829 27858
rect 5069 27176 5189 27858
rect 5294 27176 5414 27858
rect 883 25595 1003 26957
rect 1499 25595 1619 26957
rect 2122 25595 2242 26957
rect 2738 25595 2858 26957
rect 3360 25595 3480 26957
rect 3976 25595 4096 26957
rect 4599 25595 4719 26957
rect 5215 25595 5335 26957
rect 881 24008 1001 25370
rect 1501 24008 1621 25370
rect 2120 24008 2240 25370
rect 2740 24008 2860 25370
rect 3358 24008 3478 25370
rect 3978 24008 4098 25370
rect 4597 24008 4717 25370
rect 5217 24008 5337 25370
rect 881 18458 1001 19820
rect 1501 18458 1621 19820
rect 2120 18458 2240 19820
rect 2740 18458 2860 19820
rect 3358 18458 3478 19820
rect 3978 18458 4098 19820
rect 4597 18458 4717 19820
rect 5217 18458 5337 19820
rect 812 17548 932 17845
rect 1064 17548 1184 17845
rect 1318 17548 1438 17845
rect 1570 17548 1690 17845
rect 2051 17548 2171 17845
rect 2303 17548 2423 17845
rect 2557 17548 2677 17845
rect 2809 17548 2929 17845
rect 3289 17548 3409 17845
rect 3541 17548 3661 17845
rect 3795 17548 3915 17845
rect 4047 17548 4167 17845
rect 4528 17548 4648 17845
rect 4780 17548 4900 17845
rect 5034 17548 5154 17845
rect 5285 17548 5405 17845
rect 375 13056 495 15778
rect 928 14900 1048 15197
rect 1201 14900 1321 15197
rect 823 13056 943 14418
rect 1271 13056 1391 14418
rect 1719 13056 1839 15324
rect 876 9019 996 9247
rect 1100 9019 1220 9247
rect 1704 9212 1824 9440
rect 1928 9212 2048 9440
rect 876 8451 996 8643
rect 1100 8451 1220 8643
rect 1704 8533 1824 8725
rect 1928 8533 2048 8725
rect 2556 7903 2676 9265
<< mvndiff >>
rect 793 23666 881 23679
rect 793 23620 806 23666
rect 852 23620 881 23666
rect 793 23558 881 23620
rect 793 23512 806 23558
rect 852 23512 881 23558
rect 793 23450 881 23512
rect 793 23404 806 23450
rect 852 23404 881 23450
rect 793 23342 881 23404
rect 793 23296 806 23342
rect 852 23296 881 23342
rect 793 23234 881 23296
rect 793 23188 806 23234
rect 852 23188 881 23234
rect 793 23126 881 23188
rect 793 23080 806 23126
rect 852 23080 881 23126
rect 793 23018 881 23080
rect 793 22972 806 23018
rect 852 22972 881 23018
rect 793 22911 881 22972
rect 793 22865 806 22911
rect 852 22865 881 22911
rect 793 22804 881 22865
rect 793 22758 806 22804
rect 852 22758 881 22804
rect 793 22697 881 22758
rect 793 22651 806 22697
rect 852 22651 881 22697
rect 793 22590 881 22651
rect 793 22544 806 22590
rect 852 22544 881 22590
rect 793 22483 881 22544
rect 793 22437 806 22483
rect 852 22437 881 22483
rect 793 22376 881 22437
rect 793 22330 806 22376
rect 852 22330 881 22376
rect 793 22317 881 22330
rect 1001 23666 1089 23679
rect 1001 23620 1030 23666
rect 1076 23620 1089 23666
rect 1001 23558 1089 23620
rect 1001 23512 1030 23558
rect 1076 23512 1089 23558
rect 1001 23450 1089 23512
rect 1001 23404 1030 23450
rect 1076 23404 1089 23450
rect 1001 23342 1089 23404
rect 1001 23296 1030 23342
rect 1076 23296 1089 23342
rect 1001 23234 1089 23296
rect 1001 23188 1030 23234
rect 1076 23188 1089 23234
rect 1001 23126 1089 23188
rect 1001 23080 1030 23126
rect 1076 23080 1089 23126
rect 1001 23018 1089 23080
rect 1001 22972 1030 23018
rect 1076 22972 1089 23018
rect 1001 22911 1089 22972
rect 1001 22865 1030 22911
rect 1076 22865 1089 22911
rect 1001 22804 1089 22865
rect 1001 22758 1030 22804
rect 1076 22758 1089 22804
rect 1001 22697 1089 22758
rect 1001 22651 1030 22697
rect 1076 22651 1089 22697
rect 1001 22590 1089 22651
rect 1001 22544 1030 22590
rect 1076 22544 1089 22590
rect 1001 22483 1089 22544
rect 1001 22437 1030 22483
rect 1076 22437 1089 22483
rect 1001 22376 1089 22437
rect 1001 22330 1030 22376
rect 1076 22330 1089 22376
rect 1001 22317 1089 22330
rect 1413 23666 1501 23679
rect 1413 23620 1426 23666
rect 1472 23620 1501 23666
rect 1413 23558 1501 23620
rect 1413 23512 1426 23558
rect 1472 23512 1501 23558
rect 1413 23450 1501 23512
rect 1413 23404 1426 23450
rect 1472 23404 1501 23450
rect 1413 23342 1501 23404
rect 1413 23296 1426 23342
rect 1472 23296 1501 23342
rect 1413 23234 1501 23296
rect 1413 23188 1426 23234
rect 1472 23188 1501 23234
rect 1413 23126 1501 23188
rect 1413 23080 1426 23126
rect 1472 23080 1501 23126
rect 1413 23018 1501 23080
rect 1413 22972 1426 23018
rect 1472 22972 1501 23018
rect 1413 22911 1501 22972
rect 1413 22865 1426 22911
rect 1472 22865 1501 22911
rect 1413 22804 1501 22865
rect 1413 22758 1426 22804
rect 1472 22758 1501 22804
rect 1413 22697 1501 22758
rect 1413 22651 1426 22697
rect 1472 22651 1501 22697
rect 1413 22590 1501 22651
rect 1413 22544 1426 22590
rect 1472 22544 1501 22590
rect 1413 22483 1501 22544
rect 1413 22437 1426 22483
rect 1472 22437 1501 22483
rect 1413 22376 1501 22437
rect 1413 22330 1426 22376
rect 1472 22330 1501 22376
rect 1413 22317 1501 22330
rect 1621 23666 1709 23679
rect 1621 23620 1650 23666
rect 1696 23620 1709 23666
rect 1621 23558 1709 23620
rect 1621 23512 1650 23558
rect 1696 23512 1709 23558
rect 1621 23450 1709 23512
rect 1621 23404 1650 23450
rect 1696 23404 1709 23450
rect 1621 23342 1709 23404
rect 1621 23296 1650 23342
rect 1696 23296 1709 23342
rect 1621 23234 1709 23296
rect 1621 23188 1650 23234
rect 1696 23188 1709 23234
rect 1621 23126 1709 23188
rect 1621 23080 1650 23126
rect 1696 23080 1709 23126
rect 1621 23018 1709 23080
rect 1621 22972 1650 23018
rect 1696 22972 1709 23018
rect 1621 22911 1709 22972
rect 1621 22865 1650 22911
rect 1696 22865 1709 22911
rect 1621 22804 1709 22865
rect 1621 22758 1650 22804
rect 1696 22758 1709 22804
rect 1621 22697 1709 22758
rect 1621 22651 1650 22697
rect 1696 22651 1709 22697
rect 1621 22590 1709 22651
rect 1621 22544 1650 22590
rect 1696 22544 1709 22590
rect 1621 22483 1709 22544
rect 1621 22437 1650 22483
rect 1696 22437 1709 22483
rect 1621 22376 1709 22437
rect 1621 22330 1650 22376
rect 1696 22330 1709 22376
rect 1621 22317 1709 22330
rect 2032 23666 2120 23679
rect 2032 23620 2045 23666
rect 2091 23620 2120 23666
rect 2032 23558 2120 23620
rect 2032 23512 2045 23558
rect 2091 23512 2120 23558
rect 2032 23450 2120 23512
rect 2032 23404 2045 23450
rect 2091 23404 2120 23450
rect 2032 23342 2120 23404
rect 2032 23296 2045 23342
rect 2091 23296 2120 23342
rect 2032 23234 2120 23296
rect 2032 23188 2045 23234
rect 2091 23188 2120 23234
rect 2032 23126 2120 23188
rect 2032 23080 2045 23126
rect 2091 23080 2120 23126
rect 2032 23018 2120 23080
rect 2032 22972 2045 23018
rect 2091 22972 2120 23018
rect 2032 22911 2120 22972
rect 2032 22865 2045 22911
rect 2091 22865 2120 22911
rect 2032 22804 2120 22865
rect 2032 22758 2045 22804
rect 2091 22758 2120 22804
rect 2032 22697 2120 22758
rect 2032 22651 2045 22697
rect 2091 22651 2120 22697
rect 2032 22590 2120 22651
rect 2032 22544 2045 22590
rect 2091 22544 2120 22590
rect 2032 22483 2120 22544
rect 2032 22437 2045 22483
rect 2091 22437 2120 22483
rect 2032 22376 2120 22437
rect 2032 22330 2045 22376
rect 2091 22330 2120 22376
rect 2032 22317 2120 22330
rect 2240 23666 2328 23679
rect 2240 23620 2269 23666
rect 2315 23620 2328 23666
rect 2240 23558 2328 23620
rect 2240 23512 2269 23558
rect 2315 23512 2328 23558
rect 2240 23450 2328 23512
rect 2240 23404 2269 23450
rect 2315 23404 2328 23450
rect 2240 23342 2328 23404
rect 2240 23296 2269 23342
rect 2315 23296 2328 23342
rect 2240 23234 2328 23296
rect 2240 23188 2269 23234
rect 2315 23188 2328 23234
rect 2240 23126 2328 23188
rect 2240 23080 2269 23126
rect 2315 23080 2328 23126
rect 2240 23018 2328 23080
rect 2240 22972 2269 23018
rect 2315 22972 2328 23018
rect 2240 22911 2328 22972
rect 2240 22865 2269 22911
rect 2315 22865 2328 22911
rect 2240 22804 2328 22865
rect 2240 22758 2269 22804
rect 2315 22758 2328 22804
rect 2240 22697 2328 22758
rect 2240 22651 2269 22697
rect 2315 22651 2328 22697
rect 2240 22590 2328 22651
rect 2240 22544 2269 22590
rect 2315 22544 2328 22590
rect 2240 22483 2328 22544
rect 2240 22437 2269 22483
rect 2315 22437 2328 22483
rect 2240 22376 2328 22437
rect 2240 22330 2269 22376
rect 2315 22330 2328 22376
rect 2240 22317 2328 22330
rect 2652 23666 2740 23679
rect 2652 23620 2665 23666
rect 2711 23620 2740 23666
rect 2652 23558 2740 23620
rect 2652 23512 2665 23558
rect 2711 23512 2740 23558
rect 2652 23450 2740 23512
rect 2652 23404 2665 23450
rect 2711 23404 2740 23450
rect 2652 23342 2740 23404
rect 2652 23296 2665 23342
rect 2711 23296 2740 23342
rect 2652 23234 2740 23296
rect 2652 23188 2665 23234
rect 2711 23188 2740 23234
rect 2652 23126 2740 23188
rect 2652 23080 2665 23126
rect 2711 23080 2740 23126
rect 2652 23018 2740 23080
rect 2652 22972 2665 23018
rect 2711 22972 2740 23018
rect 2652 22911 2740 22972
rect 2652 22865 2665 22911
rect 2711 22865 2740 22911
rect 2652 22804 2740 22865
rect 2652 22758 2665 22804
rect 2711 22758 2740 22804
rect 2652 22697 2740 22758
rect 2652 22651 2665 22697
rect 2711 22651 2740 22697
rect 2652 22590 2740 22651
rect 2652 22544 2665 22590
rect 2711 22544 2740 22590
rect 2652 22483 2740 22544
rect 2652 22437 2665 22483
rect 2711 22437 2740 22483
rect 2652 22376 2740 22437
rect 2652 22330 2665 22376
rect 2711 22330 2740 22376
rect 2652 22317 2740 22330
rect 2860 23666 2948 23679
rect 2860 23620 2889 23666
rect 2935 23620 2948 23666
rect 2860 23558 2948 23620
rect 2860 23512 2889 23558
rect 2935 23512 2948 23558
rect 2860 23450 2948 23512
rect 2860 23404 2889 23450
rect 2935 23404 2948 23450
rect 2860 23342 2948 23404
rect 2860 23296 2889 23342
rect 2935 23296 2948 23342
rect 2860 23234 2948 23296
rect 2860 23188 2889 23234
rect 2935 23188 2948 23234
rect 2860 23126 2948 23188
rect 2860 23080 2889 23126
rect 2935 23080 2948 23126
rect 2860 23018 2948 23080
rect 2860 22972 2889 23018
rect 2935 22972 2948 23018
rect 2860 22911 2948 22972
rect 2860 22865 2889 22911
rect 2935 22865 2948 22911
rect 2860 22804 2948 22865
rect 2860 22758 2889 22804
rect 2935 22758 2948 22804
rect 2860 22697 2948 22758
rect 2860 22651 2889 22697
rect 2935 22651 2948 22697
rect 2860 22590 2948 22651
rect 2860 22544 2889 22590
rect 2935 22544 2948 22590
rect 2860 22483 2948 22544
rect 2860 22437 2889 22483
rect 2935 22437 2948 22483
rect 2860 22376 2948 22437
rect 2860 22330 2889 22376
rect 2935 22330 2948 22376
rect 2860 22317 2948 22330
rect 3270 23666 3358 23679
rect 3270 23620 3283 23666
rect 3329 23620 3358 23666
rect 3270 23558 3358 23620
rect 3270 23512 3283 23558
rect 3329 23512 3358 23558
rect 3270 23450 3358 23512
rect 3270 23404 3283 23450
rect 3329 23404 3358 23450
rect 3270 23342 3358 23404
rect 3270 23296 3283 23342
rect 3329 23296 3358 23342
rect 3270 23234 3358 23296
rect 3270 23188 3283 23234
rect 3329 23188 3358 23234
rect 3270 23126 3358 23188
rect 3270 23080 3283 23126
rect 3329 23080 3358 23126
rect 3270 23018 3358 23080
rect 3270 22972 3283 23018
rect 3329 22972 3358 23018
rect 3270 22911 3358 22972
rect 3270 22865 3283 22911
rect 3329 22865 3358 22911
rect 3270 22804 3358 22865
rect 3270 22758 3283 22804
rect 3329 22758 3358 22804
rect 3270 22697 3358 22758
rect 3270 22651 3283 22697
rect 3329 22651 3358 22697
rect 3270 22590 3358 22651
rect 3270 22544 3283 22590
rect 3329 22544 3358 22590
rect 3270 22483 3358 22544
rect 3270 22437 3283 22483
rect 3329 22437 3358 22483
rect 3270 22376 3358 22437
rect 3270 22330 3283 22376
rect 3329 22330 3358 22376
rect 3270 22317 3358 22330
rect 3478 23666 3566 23679
rect 3478 23620 3507 23666
rect 3553 23620 3566 23666
rect 3478 23558 3566 23620
rect 3478 23512 3507 23558
rect 3553 23512 3566 23558
rect 3478 23450 3566 23512
rect 3478 23404 3507 23450
rect 3553 23404 3566 23450
rect 3478 23342 3566 23404
rect 3478 23296 3507 23342
rect 3553 23296 3566 23342
rect 3478 23234 3566 23296
rect 3478 23188 3507 23234
rect 3553 23188 3566 23234
rect 3478 23126 3566 23188
rect 3478 23080 3507 23126
rect 3553 23080 3566 23126
rect 3478 23018 3566 23080
rect 3478 22972 3507 23018
rect 3553 22972 3566 23018
rect 3478 22911 3566 22972
rect 3478 22865 3507 22911
rect 3553 22865 3566 22911
rect 3478 22804 3566 22865
rect 3478 22758 3507 22804
rect 3553 22758 3566 22804
rect 3478 22697 3566 22758
rect 3478 22651 3507 22697
rect 3553 22651 3566 22697
rect 3478 22590 3566 22651
rect 3478 22544 3507 22590
rect 3553 22544 3566 22590
rect 3478 22483 3566 22544
rect 3478 22437 3507 22483
rect 3553 22437 3566 22483
rect 3478 22376 3566 22437
rect 3478 22330 3507 22376
rect 3553 22330 3566 22376
rect 3478 22317 3566 22330
rect 3890 23666 3978 23679
rect 3890 23620 3903 23666
rect 3949 23620 3978 23666
rect 3890 23558 3978 23620
rect 3890 23512 3903 23558
rect 3949 23512 3978 23558
rect 3890 23450 3978 23512
rect 3890 23404 3903 23450
rect 3949 23404 3978 23450
rect 3890 23342 3978 23404
rect 3890 23296 3903 23342
rect 3949 23296 3978 23342
rect 3890 23234 3978 23296
rect 3890 23188 3903 23234
rect 3949 23188 3978 23234
rect 3890 23126 3978 23188
rect 3890 23080 3903 23126
rect 3949 23080 3978 23126
rect 3890 23018 3978 23080
rect 3890 22972 3903 23018
rect 3949 22972 3978 23018
rect 3890 22911 3978 22972
rect 3890 22865 3903 22911
rect 3949 22865 3978 22911
rect 3890 22804 3978 22865
rect 3890 22758 3903 22804
rect 3949 22758 3978 22804
rect 3890 22697 3978 22758
rect 3890 22651 3903 22697
rect 3949 22651 3978 22697
rect 3890 22590 3978 22651
rect 3890 22544 3903 22590
rect 3949 22544 3978 22590
rect 3890 22483 3978 22544
rect 3890 22437 3903 22483
rect 3949 22437 3978 22483
rect 3890 22376 3978 22437
rect 3890 22330 3903 22376
rect 3949 22330 3978 22376
rect 3890 22317 3978 22330
rect 4098 23666 4186 23679
rect 4098 23620 4127 23666
rect 4173 23620 4186 23666
rect 4098 23558 4186 23620
rect 4098 23512 4127 23558
rect 4173 23512 4186 23558
rect 4098 23450 4186 23512
rect 4098 23404 4127 23450
rect 4173 23404 4186 23450
rect 4098 23342 4186 23404
rect 4098 23296 4127 23342
rect 4173 23296 4186 23342
rect 4098 23234 4186 23296
rect 4098 23188 4127 23234
rect 4173 23188 4186 23234
rect 4098 23126 4186 23188
rect 4098 23080 4127 23126
rect 4173 23080 4186 23126
rect 4098 23018 4186 23080
rect 4098 22972 4127 23018
rect 4173 22972 4186 23018
rect 4098 22911 4186 22972
rect 4098 22865 4127 22911
rect 4173 22865 4186 22911
rect 4098 22804 4186 22865
rect 4098 22758 4127 22804
rect 4173 22758 4186 22804
rect 4098 22697 4186 22758
rect 4098 22651 4127 22697
rect 4173 22651 4186 22697
rect 4098 22590 4186 22651
rect 4098 22544 4127 22590
rect 4173 22544 4186 22590
rect 4098 22483 4186 22544
rect 4098 22437 4127 22483
rect 4173 22437 4186 22483
rect 4098 22376 4186 22437
rect 4098 22330 4127 22376
rect 4173 22330 4186 22376
rect 4098 22317 4186 22330
rect 4509 23666 4597 23679
rect 4509 23620 4522 23666
rect 4568 23620 4597 23666
rect 4509 23558 4597 23620
rect 4509 23512 4522 23558
rect 4568 23512 4597 23558
rect 4509 23450 4597 23512
rect 4509 23404 4522 23450
rect 4568 23404 4597 23450
rect 4509 23342 4597 23404
rect 4509 23296 4522 23342
rect 4568 23296 4597 23342
rect 4509 23234 4597 23296
rect 4509 23188 4522 23234
rect 4568 23188 4597 23234
rect 4509 23126 4597 23188
rect 4509 23080 4522 23126
rect 4568 23080 4597 23126
rect 4509 23018 4597 23080
rect 4509 22972 4522 23018
rect 4568 22972 4597 23018
rect 4509 22911 4597 22972
rect 4509 22865 4522 22911
rect 4568 22865 4597 22911
rect 4509 22804 4597 22865
rect 4509 22758 4522 22804
rect 4568 22758 4597 22804
rect 4509 22697 4597 22758
rect 4509 22651 4522 22697
rect 4568 22651 4597 22697
rect 4509 22590 4597 22651
rect 4509 22544 4522 22590
rect 4568 22544 4597 22590
rect 4509 22483 4597 22544
rect 4509 22437 4522 22483
rect 4568 22437 4597 22483
rect 4509 22376 4597 22437
rect 4509 22330 4522 22376
rect 4568 22330 4597 22376
rect 4509 22317 4597 22330
rect 4717 23666 4805 23679
rect 4717 23620 4746 23666
rect 4792 23620 4805 23666
rect 4717 23558 4805 23620
rect 4717 23512 4746 23558
rect 4792 23512 4805 23558
rect 4717 23450 4805 23512
rect 4717 23404 4746 23450
rect 4792 23404 4805 23450
rect 4717 23342 4805 23404
rect 4717 23296 4746 23342
rect 4792 23296 4805 23342
rect 4717 23234 4805 23296
rect 4717 23188 4746 23234
rect 4792 23188 4805 23234
rect 4717 23126 4805 23188
rect 4717 23080 4746 23126
rect 4792 23080 4805 23126
rect 4717 23018 4805 23080
rect 4717 22972 4746 23018
rect 4792 22972 4805 23018
rect 4717 22911 4805 22972
rect 4717 22865 4746 22911
rect 4792 22865 4805 22911
rect 4717 22804 4805 22865
rect 4717 22758 4746 22804
rect 4792 22758 4805 22804
rect 4717 22697 4805 22758
rect 4717 22651 4746 22697
rect 4792 22651 4805 22697
rect 4717 22590 4805 22651
rect 4717 22544 4746 22590
rect 4792 22544 4805 22590
rect 4717 22483 4805 22544
rect 4717 22437 4746 22483
rect 4792 22437 4805 22483
rect 4717 22376 4805 22437
rect 4717 22330 4746 22376
rect 4792 22330 4805 22376
rect 4717 22317 4805 22330
rect 5129 23666 5217 23679
rect 5129 23620 5142 23666
rect 5188 23620 5217 23666
rect 5129 23558 5217 23620
rect 5129 23512 5142 23558
rect 5188 23512 5217 23558
rect 5129 23450 5217 23512
rect 5129 23404 5142 23450
rect 5188 23404 5217 23450
rect 5129 23342 5217 23404
rect 5129 23296 5142 23342
rect 5188 23296 5217 23342
rect 5129 23234 5217 23296
rect 5129 23188 5142 23234
rect 5188 23188 5217 23234
rect 5129 23126 5217 23188
rect 5129 23080 5142 23126
rect 5188 23080 5217 23126
rect 5129 23018 5217 23080
rect 5129 22972 5142 23018
rect 5188 22972 5217 23018
rect 5129 22911 5217 22972
rect 5129 22865 5142 22911
rect 5188 22865 5217 22911
rect 5129 22804 5217 22865
rect 5129 22758 5142 22804
rect 5188 22758 5217 22804
rect 5129 22697 5217 22758
rect 5129 22651 5142 22697
rect 5188 22651 5217 22697
rect 5129 22590 5217 22651
rect 5129 22544 5142 22590
rect 5188 22544 5217 22590
rect 5129 22483 5217 22544
rect 5129 22437 5142 22483
rect 5188 22437 5217 22483
rect 5129 22376 5217 22437
rect 5129 22330 5142 22376
rect 5188 22330 5217 22376
rect 5129 22317 5217 22330
rect 5337 23666 5425 23679
rect 5337 23620 5366 23666
rect 5412 23620 5425 23666
rect 5337 23558 5425 23620
rect 5337 23512 5366 23558
rect 5412 23512 5425 23558
rect 5337 23450 5425 23512
rect 5337 23404 5366 23450
rect 5412 23404 5425 23450
rect 5337 23342 5425 23404
rect 5337 23296 5366 23342
rect 5412 23296 5425 23342
rect 5337 23234 5425 23296
rect 5337 23188 5366 23234
rect 5412 23188 5425 23234
rect 5337 23126 5425 23188
rect 5337 23080 5366 23126
rect 5412 23080 5425 23126
rect 5337 23018 5425 23080
rect 5337 22972 5366 23018
rect 5412 22972 5425 23018
rect 5337 22911 5425 22972
rect 5337 22865 5366 22911
rect 5412 22865 5425 22911
rect 5337 22804 5425 22865
rect 5337 22758 5366 22804
rect 5412 22758 5425 22804
rect 5337 22697 5425 22758
rect 5337 22651 5366 22697
rect 5412 22651 5425 22697
rect 5337 22590 5425 22651
rect 5337 22544 5366 22590
rect 5412 22544 5425 22590
rect 5337 22483 5425 22544
rect 5337 22437 5366 22483
rect 5412 22437 5425 22483
rect 5337 22376 5425 22437
rect 5337 22330 5366 22376
rect 5412 22330 5425 22376
rect 5337 22317 5425 22330
rect 793 21662 881 21675
rect 793 21616 806 21662
rect 852 21616 881 21662
rect 793 21554 881 21616
rect 793 21508 806 21554
rect 852 21508 881 21554
rect 793 21446 881 21508
rect 793 21400 806 21446
rect 852 21400 881 21446
rect 793 21338 881 21400
rect 793 21292 806 21338
rect 852 21292 881 21338
rect 793 21230 881 21292
rect 793 21184 806 21230
rect 852 21184 881 21230
rect 793 21122 881 21184
rect 793 21076 806 21122
rect 852 21076 881 21122
rect 793 21014 881 21076
rect 793 20968 806 21014
rect 852 20968 881 21014
rect 793 20907 881 20968
rect 793 20861 806 20907
rect 852 20861 881 20907
rect 793 20800 881 20861
rect 793 20754 806 20800
rect 852 20754 881 20800
rect 793 20693 881 20754
rect 793 20647 806 20693
rect 852 20647 881 20693
rect 793 20586 881 20647
rect 793 20540 806 20586
rect 852 20540 881 20586
rect 793 20479 881 20540
rect 793 20433 806 20479
rect 852 20433 881 20479
rect 793 20372 881 20433
rect 793 20326 806 20372
rect 852 20326 881 20372
rect 793 20313 881 20326
rect 1001 21662 1089 21675
rect 1001 21616 1030 21662
rect 1076 21616 1089 21662
rect 1001 21554 1089 21616
rect 1001 21508 1030 21554
rect 1076 21508 1089 21554
rect 1001 21446 1089 21508
rect 1001 21400 1030 21446
rect 1076 21400 1089 21446
rect 1001 21338 1089 21400
rect 1001 21292 1030 21338
rect 1076 21292 1089 21338
rect 1001 21230 1089 21292
rect 1001 21184 1030 21230
rect 1076 21184 1089 21230
rect 1001 21122 1089 21184
rect 1001 21076 1030 21122
rect 1076 21076 1089 21122
rect 1001 21014 1089 21076
rect 1001 20968 1030 21014
rect 1076 20968 1089 21014
rect 1001 20907 1089 20968
rect 1001 20861 1030 20907
rect 1076 20861 1089 20907
rect 1001 20800 1089 20861
rect 1001 20754 1030 20800
rect 1076 20754 1089 20800
rect 1001 20693 1089 20754
rect 1001 20647 1030 20693
rect 1076 20647 1089 20693
rect 1001 20586 1089 20647
rect 1001 20540 1030 20586
rect 1076 20540 1089 20586
rect 1001 20479 1089 20540
rect 1001 20433 1030 20479
rect 1076 20433 1089 20479
rect 1001 20372 1089 20433
rect 1001 20326 1030 20372
rect 1076 20326 1089 20372
rect 1001 20313 1089 20326
rect 1413 21662 1501 21675
rect 1413 21616 1426 21662
rect 1472 21616 1501 21662
rect 1413 21554 1501 21616
rect 1413 21508 1426 21554
rect 1472 21508 1501 21554
rect 1413 21446 1501 21508
rect 1413 21400 1426 21446
rect 1472 21400 1501 21446
rect 1413 21338 1501 21400
rect 1413 21292 1426 21338
rect 1472 21292 1501 21338
rect 1413 21230 1501 21292
rect 1413 21184 1426 21230
rect 1472 21184 1501 21230
rect 1413 21122 1501 21184
rect 1413 21076 1426 21122
rect 1472 21076 1501 21122
rect 1413 21014 1501 21076
rect 1413 20968 1426 21014
rect 1472 20968 1501 21014
rect 1413 20907 1501 20968
rect 1413 20861 1426 20907
rect 1472 20861 1501 20907
rect 1413 20800 1501 20861
rect 1413 20754 1426 20800
rect 1472 20754 1501 20800
rect 1413 20693 1501 20754
rect 1413 20647 1426 20693
rect 1472 20647 1501 20693
rect 1413 20586 1501 20647
rect 1413 20540 1426 20586
rect 1472 20540 1501 20586
rect 1413 20479 1501 20540
rect 1413 20433 1426 20479
rect 1472 20433 1501 20479
rect 1413 20372 1501 20433
rect 1413 20326 1426 20372
rect 1472 20326 1501 20372
rect 1413 20313 1501 20326
rect 1621 21662 1709 21675
rect 1621 21616 1650 21662
rect 1696 21616 1709 21662
rect 1621 21554 1709 21616
rect 1621 21508 1650 21554
rect 1696 21508 1709 21554
rect 1621 21446 1709 21508
rect 1621 21400 1650 21446
rect 1696 21400 1709 21446
rect 1621 21338 1709 21400
rect 1621 21292 1650 21338
rect 1696 21292 1709 21338
rect 1621 21230 1709 21292
rect 1621 21184 1650 21230
rect 1696 21184 1709 21230
rect 1621 21122 1709 21184
rect 1621 21076 1650 21122
rect 1696 21076 1709 21122
rect 1621 21014 1709 21076
rect 1621 20968 1650 21014
rect 1696 20968 1709 21014
rect 1621 20907 1709 20968
rect 1621 20861 1650 20907
rect 1696 20861 1709 20907
rect 1621 20800 1709 20861
rect 1621 20754 1650 20800
rect 1696 20754 1709 20800
rect 1621 20693 1709 20754
rect 1621 20647 1650 20693
rect 1696 20647 1709 20693
rect 1621 20586 1709 20647
rect 1621 20540 1650 20586
rect 1696 20540 1709 20586
rect 1621 20479 1709 20540
rect 1621 20433 1650 20479
rect 1696 20433 1709 20479
rect 1621 20372 1709 20433
rect 1621 20326 1650 20372
rect 1696 20326 1709 20372
rect 1621 20313 1709 20326
rect 2032 21662 2120 21675
rect 2032 21616 2045 21662
rect 2091 21616 2120 21662
rect 2032 21554 2120 21616
rect 2032 21508 2045 21554
rect 2091 21508 2120 21554
rect 2032 21446 2120 21508
rect 2032 21400 2045 21446
rect 2091 21400 2120 21446
rect 2032 21338 2120 21400
rect 2032 21292 2045 21338
rect 2091 21292 2120 21338
rect 2032 21230 2120 21292
rect 2032 21184 2045 21230
rect 2091 21184 2120 21230
rect 2032 21122 2120 21184
rect 2032 21076 2045 21122
rect 2091 21076 2120 21122
rect 2032 21014 2120 21076
rect 2032 20968 2045 21014
rect 2091 20968 2120 21014
rect 2032 20907 2120 20968
rect 2032 20861 2045 20907
rect 2091 20861 2120 20907
rect 2032 20800 2120 20861
rect 2032 20754 2045 20800
rect 2091 20754 2120 20800
rect 2032 20693 2120 20754
rect 2032 20647 2045 20693
rect 2091 20647 2120 20693
rect 2032 20586 2120 20647
rect 2032 20540 2045 20586
rect 2091 20540 2120 20586
rect 2032 20479 2120 20540
rect 2032 20433 2045 20479
rect 2091 20433 2120 20479
rect 2032 20372 2120 20433
rect 2032 20326 2045 20372
rect 2091 20326 2120 20372
rect 2032 20313 2120 20326
rect 2240 21662 2328 21675
rect 2240 21616 2269 21662
rect 2315 21616 2328 21662
rect 2240 21554 2328 21616
rect 2240 21508 2269 21554
rect 2315 21508 2328 21554
rect 2240 21446 2328 21508
rect 2240 21400 2269 21446
rect 2315 21400 2328 21446
rect 2240 21338 2328 21400
rect 2240 21292 2269 21338
rect 2315 21292 2328 21338
rect 2240 21230 2328 21292
rect 2240 21184 2269 21230
rect 2315 21184 2328 21230
rect 2240 21122 2328 21184
rect 2240 21076 2269 21122
rect 2315 21076 2328 21122
rect 2240 21014 2328 21076
rect 2240 20968 2269 21014
rect 2315 20968 2328 21014
rect 2240 20907 2328 20968
rect 2240 20861 2269 20907
rect 2315 20861 2328 20907
rect 2240 20800 2328 20861
rect 2240 20754 2269 20800
rect 2315 20754 2328 20800
rect 2240 20693 2328 20754
rect 2240 20647 2269 20693
rect 2315 20647 2328 20693
rect 2240 20586 2328 20647
rect 2240 20540 2269 20586
rect 2315 20540 2328 20586
rect 2240 20479 2328 20540
rect 2240 20433 2269 20479
rect 2315 20433 2328 20479
rect 2240 20372 2328 20433
rect 2240 20326 2269 20372
rect 2315 20326 2328 20372
rect 2240 20313 2328 20326
rect 2652 21662 2740 21675
rect 2652 21616 2665 21662
rect 2711 21616 2740 21662
rect 2652 21554 2740 21616
rect 2652 21508 2665 21554
rect 2711 21508 2740 21554
rect 2652 21446 2740 21508
rect 2652 21400 2665 21446
rect 2711 21400 2740 21446
rect 2652 21338 2740 21400
rect 2652 21292 2665 21338
rect 2711 21292 2740 21338
rect 2652 21230 2740 21292
rect 2652 21184 2665 21230
rect 2711 21184 2740 21230
rect 2652 21122 2740 21184
rect 2652 21076 2665 21122
rect 2711 21076 2740 21122
rect 2652 21014 2740 21076
rect 2652 20968 2665 21014
rect 2711 20968 2740 21014
rect 2652 20907 2740 20968
rect 2652 20861 2665 20907
rect 2711 20861 2740 20907
rect 2652 20800 2740 20861
rect 2652 20754 2665 20800
rect 2711 20754 2740 20800
rect 2652 20693 2740 20754
rect 2652 20647 2665 20693
rect 2711 20647 2740 20693
rect 2652 20586 2740 20647
rect 2652 20540 2665 20586
rect 2711 20540 2740 20586
rect 2652 20479 2740 20540
rect 2652 20433 2665 20479
rect 2711 20433 2740 20479
rect 2652 20372 2740 20433
rect 2652 20326 2665 20372
rect 2711 20326 2740 20372
rect 2652 20313 2740 20326
rect 2860 21662 2948 21675
rect 2860 21616 2889 21662
rect 2935 21616 2948 21662
rect 2860 21554 2948 21616
rect 2860 21508 2889 21554
rect 2935 21508 2948 21554
rect 2860 21446 2948 21508
rect 2860 21400 2889 21446
rect 2935 21400 2948 21446
rect 2860 21338 2948 21400
rect 2860 21292 2889 21338
rect 2935 21292 2948 21338
rect 2860 21230 2948 21292
rect 2860 21184 2889 21230
rect 2935 21184 2948 21230
rect 2860 21122 2948 21184
rect 2860 21076 2889 21122
rect 2935 21076 2948 21122
rect 2860 21014 2948 21076
rect 2860 20968 2889 21014
rect 2935 20968 2948 21014
rect 2860 20907 2948 20968
rect 2860 20861 2889 20907
rect 2935 20861 2948 20907
rect 2860 20800 2948 20861
rect 2860 20754 2889 20800
rect 2935 20754 2948 20800
rect 2860 20693 2948 20754
rect 2860 20647 2889 20693
rect 2935 20647 2948 20693
rect 2860 20586 2948 20647
rect 2860 20540 2889 20586
rect 2935 20540 2948 20586
rect 2860 20479 2948 20540
rect 2860 20433 2889 20479
rect 2935 20433 2948 20479
rect 2860 20372 2948 20433
rect 2860 20326 2889 20372
rect 2935 20326 2948 20372
rect 2860 20313 2948 20326
rect 3270 21662 3358 21675
rect 3270 21616 3283 21662
rect 3329 21616 3358 21662
rect 3270 21554 3358 21616
rect 3270 21508 3283 21554
rect 3329 21508 3358 21554
rect 3270 21446 3358 21508
rect 3270 21400 3283 21446
rect 3329 21400 3358 21446
rect 3270 21338 3358 21400
rect 3270 21292 3283 21338
rect 3329 21292 3358 21338
rect 3270 21230 3358 21292
rect 3270 21184 3283 21230
rect 3329 21184 3358 21230
rect 3270 21122 3358 21184
rect 3270 21076 3283 21122
rect 3329 21076 3358 21122
rect 3270 21014 3358 21076
rect 3270 20968 3283 21014
rect 3329 20968 3358 21014
rect 3270 20907 3358 20968
rect 3270 20861 3283 20907
rect 3329 20861 3358 20907
rect 3270 20800 3358 20861
rect 3270 20754 3283 20800
rect 3329 20754 3358 20800
rect 3270 20693 3358 20754
rect 3270 20647 3283 20693
rect 3329 20647 3358 20693
rect 3270 20586 3358 20647
rect 3270 20540 3283 20586
rect 3329 20540 3358 20586
rect 3270 20479 3358 20540
rect 3270 20433 3283 20479
rect 3329 20433 3358 20479
rect 3270 20372 3358 20433
rect 3270 20326 3283 20372
rect 3329 20326 3358 20372
rect 3270 20313 3358 20326
rect 3478 21662 3566 21675
rect 3478 21616 3507 21662
rect 3553 21616 3566 21662
rect 3478 21554 3566 21616
rect 3478 21508 3507 21554
rect 3553 21508 3566 21554
rect 3478 21446 3566 21508
rect 3478 21400 3507 21446
rect 3553 21400 3566 21446
rect 3478 21338 3566 21400
rect 3478 21292 3507 21338
rect 3553 21292 3566 21338
rect 3478 21230 3566 21292
rect 3478 21184 3507 21230
rect 3553 21184 3566 21230
rect 3478 21122 3566 21184
rect 3478 21076 3507 21122
rect 3553 21076 3566 21122
rect 3478 21014 3566 21076
rect 3478 20968 3507 21014
rect 3553 20968 3566 21014
rect 3478 20907 3566 20968
rect 3478 20861 3507 20907
rect 3553 20861 3566 20907
rect 3478 20800 3566 20861
rect 3478 20754 3507 20800
rect 3553 20754 3566 20800
rect 3478 20693 3566 20754
rect 3478 20647 3507 20693
rect 3553 20647 3566 20693
rect 3478 20586 3566 20647
rect 3478 20540 3507 20586
rect 3553 20540 3566 20586
rect 3478 20479 3566 20540
rect 3478 20433 3507 20479
rect 3553 20433 3566 20479
rect 3478 20372 3566 20433
rect 3478 20326 3507 20372
rect 3553 20326 3566 20372
rect 3478 20313 3566 20326
rect 3890 21662 3978 21675
rect 3890 21616 3903 21662
rect 3949 21616 3978 21662
rect 3890 21554 3978 21616
rect 3890 21508 3903 21554
rect 3949 21508 3978 21554
rect 3890 21446 3978 21508
rect 3890 21400 3903 21446
rect 3949 21400 3978 21446
rect 3890 21338 3978 21400
rect 3890 21292 3903 21338
rect 3949 21292 3978 21338
rect 3890 21230 3978 21292
rect 3890 21184 3903 21230
rect 3949 21184 3978 21230
rect 3890 21122 3978 21184
rect 3890 21076 3903 21122
rect 3949 21076 3978 21122
rect 3890 21014 3978 21076
rect 3890 20968 3903 21014
rect 3949 20968 3978 21014
rect 3890 20907 3978 20968
rect 3890 20861 3903 20907
rect 3949 20861 3978 20907
rect 3890 20800 3978 20861
rect 3890 20754 3903 20800
rect 3949 20754 3978 20800
rect 3890 20693 3978 20754
rect 3890 20647 3903 20693
rect 3949 20647 3978 20693
rect 3890 20586 3978 20647
rect 3890 20540 3903 20586
rect 3949 20540 3978 20586
rect 3890 20479 3978 20540
rect 3890 20433 3903 20479
rect 3949 20433 3978 20479
rect 3890 20372 3978 20433
rect 3890 20326 3903 20372
rect 3949 20326 3978 20372
rect 3890 20313 3978 20326
rect 4098 21662 4186 21675
rect 4098 21616 4127 21662
rect 4173 21616 4186 21662
rect 4098 21554 4186 21616
rect 4098 21508 4127 21554
rect 4173 21508 4186 21554
rect 4098 21446 4186 21508
rect 4098 21400 4127 21446
rect 4173 21400 4186 21446
rect 4098 21338 4186 21400
rect 4098 21292 4127 21338
rect 4173 21292 4186 21338
rect 4098 21230 4186 21292
rect 4098 21184 4127 21230
rect 4173 21184 4186 21230
rect 4098 21122 4186 21184
rect 4098 21076 4127 21122
rect 4173 21076 4186 21122
rect 4098 21014 4186 21076
rect 4098 20968 4127 21014
rect 4173 20968 4186 21014
rect 4098 20907 4186 20968
rect 4098 20861 4127 20907
rect 4173 20861 4186 20907
rect 4098 20800 4186 20861
rect 4098 20754 4127 20800
rect 4173 20754 4186 20800
rect 4098 20693 4186 20754
rect 4098 20647 4127 20693
rect 4173 20647 4186 20693
rect 4098 20586 4186 20647
rect 4098 20540 4127 20586
rect 4173 20540 4186 20586
rect 4098 20479 4186 20540
rect 4098 20433 4127 20479
rect 4173 20433 4186 20479
rect 4098 20372 4186 20433
rect 4098 20326 4127 20372
rect 4173 20326 4186 20372
rect 4098 20313 4186 20326
rect 4509 21662 4597 21675
rect 4509 21616 4522 21662
rect 4568 21616 4597 21662
rect 4509 21554 4597 21616
rect 4509 21508 4522 21554
rect 4568 21508 4597 21554
rect 4509 21446 4597 21508
rect 4509 21400 4522 21446
rect 4568 21400 4597 21446
rect 4509 21338 4597 21400
rect 4509 21292 4522 21338
rect 4568 21292 4597 21338
rect 4509 21230 4597 21292
rect 4509 21184 4522 21230
rect 4568 21184 4597 21230
rect 4509 21122 4597 21184
rect 4509 21076 4522 21122
rect 4568 21076 4597 21122
rect 4509 21014 4597 21076
rect 4509 20968 4522 21014
rect 4568 20968 4597 21014
rect 4509 20907 4597 20968
rect 4509 20861 4522 20907
rect 4568 20861 4597 20907
rect 4509 20800 4597 20861
rect 4509 20754 4522 20800
rect 4568 20754 4597 20800
rect 4509 20693 4597 20754
rect 4509 20647 4522 20693
rect 4568 20647 4597 20693
rect 4509 20586 4597 20647
rect 4509 20540 4522 20586
rect 4568 20540 4597 20586
rect 4509 20479 4597 20540
rect 4509 20433 4522 20479
rect 4568 20433 4597 20479
rect 4509 20372 4597 20433
rect 4509 20326 4522 20372
rect 4568 20326 4597 20372
rect 4509 20313 4597 20326
rect 4717 21662 4805 21675
rect 4717 21616 4746 21662
rect 4792 21616 4805 21662
rect 4717 21554 4805 21616
rect 4717 21508 4746 21554
rect 4792 21508 4805 21554
rect 4717 21446 4805 21508
rect 4717 21400 4746 21446
rect 4792 21400 4805 21446
rect 4717 21338 4805 21400
rect 4717 21292 4746 21338
rect 4792 21292 4805 21338
rect 4717 21230 4805 21292
rect 4717 21184 4746 21230
rect 4792 21184 4805 21230
rect 4717 21122 4805 21184
rect 4717 21076 4746 21122
rect 4792 21076 4805 21122
rect 4717 21014 4805 21076
rect 4717 20968 4746 21014
rect 4792 20968 4805 21014
rect 4717 20907 4805 20968
rect 4717 20861 4746 20907
rect 4792 20861 4805 20907
rect 4717 20800 4805 20861
rect 4717 20754 4746 20800
rect 4792 20754 4805 20800
rect 4717 20693 4805 20754
rect 4717 20647 4746 20693
rect 4792 20647 4805 20693
rect 4717 20586 4805 20647
rect 4717 20540 4746 20586
rect 4792 20540 4805 20586
rect 4717 20479 4805 20540
rect 4717 20433 4746 20479
rect 4792 20433 4805 20479
rect 4717 20372 4805 20433
rect 4717 20326 4746 20372
rect 4792 20326 4805 20372
rect 4717 20313 4805 20326
rect 5129 21662 5217 21675
rect 5129 21616 5142 21662
rect 5188 21616 5217 21662
rect 5129 21554 5217 21616
rect 5129 21508 5142 21554
rect 5188 21508 5217 21554
rect 5129 21446 5217 21508
rect 5129 21400 5142 21446
rect 5188 21400 5217 21446
rect 5129 21338 5217 21400
rect 5129 21292 5142 21338
rect 5188 21292 5217 21338
rect 5129 21230 5217 21292
rect 5129 21184 5142 21230
rect 5188 21184 5217 21230
rect 5129 21122 5217 21184
rect 5129 21076 5142 21122
rect 5188 21076 5217 21122
rect 5129 21014 5217 21076
rect 5129 20968 5142 21014
rect 5188 20968 5217 21014
rect 5129 20907 5217 20968
rect 5129 20861 5142 20907
rect 5188 20861 5217 20907
rect 5129 20800 5217 20861
rect 5129 20754 5142 20800
rect 5188 20754 5217 20800
rect 5129 20693 5217 20754
rect 5129 20647 5142 20693
rect 5188 20647 5217 20693
rect 5129 20586 5217 20647
rect 5129 20540 5142 20586
rect 5188 20540 5217 20586
rect 5129 20479 5217 20540
rect 5129 20433 5142 20479
rect 5188 20433 5217 20479
rect 5129 20372 5217 20433
rect 5129 20326 5142 20372
rect 5188 20326 5217 20372
rect 5129 20313 5217 20326
rect 5337 21662 5425 21675
rect 5337 21616 5366 21662
rect 5412 21616 5425 21662
rect 5337 21554 5425 21616
rect 5337 21508 5366 21554
rect 5412 21508 5425 21554
rect 5337 21446 5425 21508
rect 5337 21400 5366 21446
rect 5412 21400 5425 21446
rect 5337 21338 5425 21400
rect 5337 21292 5366 21338
rect 5412 21292 5425 21338
rect 5337 21230 5425 21292
rect 5337 21184 5366 21230
rect 5412 21184 5425 21230
rect 5337 21122 5425 21184
rect 5337 21076 5366 21122
rect 5412 21076 5425 21122
rect 5337 21014 5425 21076
rect 5337 20968 5366 21014
rect 5412 20968 5425 21014
rect 5337 20907 5425 20968
rect 5337 20861 5366 20907
rect 5412 20861 5425 20907
rect 5337 20800 5425 20861
rect 5337 20754 5366 20800
rect 5412 20754 5425 20800
rect 5337 20693 5425 20754
rect 5337 20647 5366 20693
rect 5412 20647 5425 20693
rect 5337 20586 5425 20647
rect 5337 20540 5366 20586
rect 5412 20540 5425 20586
rect 5337 20479 5425 20540
rect 5337 20433 5366 20479
rect 5412 20433 5425 20479
rect 5337 20372 5425 20433
rect 5337 20326 5366 20372
rect 5412 20326 5425 20372
rect 5337 20313 5425 20326
rect 767 17223 855 17257
rect 767 17177 780 17223
rect 826 17177 855 17223
rect 767 17143 855 17177
rect 975 17223 1079 17257
rect 975 17177 1004 17223
rect 1050 17177 1079 17223
rect 975 17143 1079 17177
rect 1199 17223 1303 17257
rect 1199 17177 1228 17223
rect 1274 17177 1303 17223
rect 1199 17143 1303 17177
rect 1423 17223 1527 17257
rect 1423 17177 1452 17223
rect 1498 17177 1527 17223
rect 1423 17143 1527 17177
rect 1647 17223 1735 17257
rect 1647 17177 1676 17223
rect 1722 17177 1735 17223
rect 1647 17143 1735 17177
rect 2006 17223 2094 17257
rect 2006 17177 2019 17223
rect 2065 17177 2094 17223
rect 2006 17143 2094 17177
rect 2214 17223 2318 17257
rect 2214 17177 2243 17223
rect 2289 17177 2318 17223
rect 2214 17143 2318 17177
rect 2438 17223 2542 17257
rect 2438 17177 2467 17223
rect 2513 17177 2542 17223
rect 2438 17143 2542 17177
rect 2662 17223 2766 17257
rect 2662 17177 2691 17223
rect 2737 17177 2766 17223
rect 2662 17143 2766 17177
rect 2886 17223 2974 17257
rect 2886 17177 2915 17223
rect 2961 17177 2974 17223
rect 2886 17143 2974 17177
rect 3244 17223 3332 17257
rect 3244 17177 3257 17223
rect 3303 17177 3332 17223
rect 3244 17143 3332 17177
rect 3452 17223 3556 17257
rect 3452 17177 3481 17223
rect 3527 17177 3556 17223
rect 3452 17143 3556 17177
rect 3676 17223 3780 17257
rect 3676 17177 3705 17223
rect 3751 17177 3780 17223
rect 3676 17143 3780 17177
rect 3900 17223 4004 17257
rect 3900 17177 3929 17223
rect 3975 17177 4004 17223
rect 3900 17143 4004 17177
rect 4124 17223 4212 17257
rect 4124 17177 4153 17223
rect 4199 17177 4212 17223
rect 4124 17143 4212 17177
rect 4483 17223 4571 17257
rect 4483 17177 4496 17223
rect 4542 17177 4571 17223
rect 4483 17143 4571 17177
rect 4691 17223 4795 17257
rect 4691 17177 4720 17223
rect 4766 17177 4795 17223
rect 4691 17143 4795 17177
rect 4915 17223 5019 17257
rect 4915 17177 4944 17223
rect 4990 17177 5019 17223
rect 4915 17143 5019 17177
rect 5139 17223 5243 17257
rect 5139 17177 5168 17223
rect 5214 17177 5243 17223
rect 5139 17143 5243 17177
rect 5363 17223 5451 17257
rect 5363 17177 5392 17223
rect 5438 17177 5451 17223
rect 5363 17143 5451 17177
rect 904 15591 1043 15704
rect 904 15545 948 15591
rect 994 15545 1043 15591
rect 904 15476 1043 15545
rect 1163 15591 1301 15704
rect 1163 15545 1211 15591
rect 1257 15545 1301 15591
rect 1163 15476 1301 15545
rect 287 12607 375 12620
rect 287 9911 300 12607
rect 346 9911 375 12607
rect 287 9898 375 9911
rect 495 12607 583 12620
rect 495 9911 524 12607
rect 570 9911 583 12607
rect 735 12606 823 12619
rect 735 12560 748 12606
rect 794 12560 823 12606
rect 735 12502 823 12560
rect 735 12456 748 12502
rect 794 12456 823 12502
rect 735 12398 823 12456
rect 735 12352 748 12398
rect 794 12352 823 12398
rect 735 12294 823 12352
rect 735 12248 748 12294
rect 794 12248 823 12294
rect 735 12190 823 12248
rect 735 12144 748 12190
rect 794 12144 823 12190
rect 735 12086 823 12144
rect 735 12040 748 12086
rect 794 12040 823 12086
rect 735 11982 823 12040
rect 735 11936 748 11982
rect 794 11936 823 11982
rect 735 11878 823 11936
rect 735 11832 748 11878
rect 794 11832 823 11878
rect 735 11774 823 11832
rect 735 11728 748 11774
rect 794 11728 823 11774
rect 735 11670 823 11728
rect 735 11624 748 11670
rect 794 11624 823 11670
rect 735 11565 823 11624
rect 735 11519 748 11565
rect 794 11519 823 11565
rect 735 11460 823 11519
rect 735 11414 748 11460
rect 794 11414 823 11460
rect 735 11355 823 11414
rect 735 11309 748 11355
rect 794 11309 823 11355
rect 735 11250 823 11309
rect 735 11204 748 11250
rect 794 11204 823 11250
rect 735 11145 823 11204
rect 735 11099 748 11145
rect 794 11099 823 11145
rect 735 11040 823 11099
rect 735 10994 748 11040
rect 794 10994 823 11040
rect 735 10935 823 10994
rect 735 10889 748 10935
rect 794 10889 823 10935
rect 735 10830 823 10889
rect 735 10784 748 10830
rect 794 10784 823 10830
rect 735 10725 823 10784
rect 735 10679 748 10725
rect 794 10679 823 10725
rect 735 10620 823 10679
rect 735 10574 748 10620
rect 794 10574 823 10620
rect 735 10515 823 10574
rect 735 10469 748 10515
rect 794 10469 823 10515
rect 735 10410 823 10469
rect 735 10364 748 10410
rect 794 10364 823 10410
rect 735 10351 823 10364
rect 943 12606 1031 12619
rect 943 12560 972 12606
rect 1018 12560 1031 12606
rect 943 12502 1031 12560
rect 943 12456 972 12502
rect 1018 12456 1031 12502
rect 943 12398 1031 12456
rect 943 12352 972 12398
rect 1018 12352 1031 12398
rect 943 12294 1031 12352
rect 943 12248 972 12294
rect 1018 12248 1031 12294
rect 943 12190 1031 12248
rect 943 12144 972 12190
rect 1018 12144 1031 12190
rect 943 12086 1031 12144
rect 943 12040 972 12086
rect 1018 12040 1031 12086
rect 943 11982 1031 12040
rect 943 11936 972 11982
rect 1018 11936 1031 11982
rect 943 11878 1031 11936
rect 943 11832 972 11878
rect 1018 11832 1031 11878
rect 943 11774 1031 11832
rect 943 11728 972 11774
rect 1018 11728 1031 11774
rect 943 11670 1031 11728
rect 943 11624 972 11670
rect 1018 11624 1031 11670
rect 943 11565 1031 11624
rect 943 11519 972 11565
rect 1018 11519 1031 11565
rect 943 11460 1031 11519
rect 943 11414 972 11460
rect 1018 11414 1031 11460
rect 943 11355 1031 11414
rect 943 11309 972 11355
rect 1018 11309 1031 11355
rect 943 11250 1031 11309
rect 943 11204 972 11250
rect 1018 11204 1031 11250
rect 943 11145 1031 11204
rect 943 11099 972 11145
rect 1018 11099 1031 11145
rect 943 11040 1031 11099
rect 943 10994 972 11040
rect 1018 10994 1031 11040
rect 943 10935 1031 10994
rect 943 10889 972 10935
rect 1018 10889 1031 10935
rect 943 10830 1031 10889
rect 943 10784 972 10830
rect 1018 10784 1031 10830
rect 943 10725 1031 10784
rect 943 10679 972 10725
rect 1018 10679 1031 10725
rect 943 10620 1031 10679
rect 943 10574 972 10620
rect 1018 10574 1031 10620
rect 943 10515 1031 10574
rect 943 10469 972 10515
rect 1018 10469 1031 10515
rect 943 10410 1031 10469
rect 943 10364 972 10410
rect 1018 10364 1031 10410
rect 943 10351 1031 10364
rect 1183 12606 1271 12619
rect 1183 12560 1196 12606
rect 1242 12560 1271 12606
rect 1183 12502 1271 12560
rect 1183 12456 1196 12502
rect 1242 12456 1271 12502
rect 1183 12398 1271 12456
rect 1183 12352 1196 12398
rect 1242 12352 1271 12398
rect 1183 12294 1271 12352
rect 1183 12248 1196 12294
rect 1242 12248 1271 12294
rect 1183 12190 1271 12248
rect 1183 12144 1196 12190
rect 1242 12144 1271 12190
rect 1183 12086 1271 12144
rect 1183 12040 1196 12086
rect 1242 12040 1271 12086
rect 1183 11982 1271 12040
rect 1183 11936 1196 11982
rect 1242 11936 1271 11982
rect 1183 11878 1271 11936
rect 1183 11832 1196 11878
rect 1242 11832 1271 11878
rect 1183 11774 1271 11832
rect 1183 11728 1196 11774
rect 1242 11728 1271 11774
rect 1183 11670 1271 11728
rect 1183 11624 1196 11670
rect 1242 11624 1271 11670
rect 1183 11565 1271 11624
rect 1183 11519 1196 11565
rect 1242 11519 1271 11565
rect 1183 11460 1271 11519
rect 1183 11414 1196 11460
rect 1242 11414 1271 11460
rect 1183 11355 1271 11414
rect 1183 11309 1196 11355
rect 1242 11309 1271 11355
rect 1183 11250 1271 11309
rect 1183 11204 1196 11250
rect 1242 11204 1271 11250
rect 1183 11145 1271 11204
rect 1183 11099 1196 11145
rect 1242 11099 1271 11145
rect 1183 11040 1271 11099
rect 1183 10994 1196 11040
rect 1242 10994 1271 11040
rect 1183 10935 1271 10994
rect 1183 10889 1196 10935
rect 1242 10889 1271 10935
rect 1183 10830 1271 10889
rect 1183 10784 1196 10830
rect 1242 10784 1271 10830
rect 1183 10725 1271 10784
rect 1183 10679 1196 10725
rect 1242 10679 1271 10725
rect 1183 10620 1271 10679
rect 1183 10574 1196 10620
rect 1242 10574 1271 10620
rect 1183 10515 1271 10574
rect 1183 10469 1196 10515
rect 1242 10469 1271 10515
rect 1183 10410 1271 10469
rect 1183 10364 1196 10410
rect 1242 10364 1271 10410
rect 1183 10351 1271 10364
rect 1391 12606 1479 12619
rect 1391 12560 1420 12606
rect 1466 12560 1479 12606
rect 1391 12502 1479 12560
rect 1391 12456 1420 12502
rect 1466 12456 1479 12502
rect 1391 12398 1479 12456
rect 1391 12352 1420 12398
rect 1466 12352 1479 12398
rect 1391 12294 1479 12352
rect 1391 12248 1420 12294
rect 1466 12248 1479 12294
rect 1391 12190 1479 12248
rect 1391 12144 1420 12190
rect 1466 12144 1479 12190
rect 1391 12086 1479 12144
rect 1391 12040 1420 12086
rect 1466 12040 1479 12086
rect 1391 11982 1479 12040
rect 1391 11936 1420 11982
rect 1466 11936 1479 11982
rect 1391 11878 1479 11936
rect 1391 11832 1420 11878
rect 1466 11832 1479 11878
rect 1391 11774 1479 11832
rect 1391 11728 1420 11774
rect 1466 11728 1479 11774
rect 1391 11670 1479 11728
rect 1391 11624 1420 11670
rect 1466 11624 1479 11670
rect 1391 11565 1479 11624
rect 1391 11519 1420 11565
rect 1466 11519 1479 11565
rect 1391 11460 1479 11519
rect 1391 11414 1420 11460
rect 1466 11414 1479 11460
rect 1391 11355 1479 11414
rect 1391 11309 1420 11355
rect 1466 11309 1479 11355
rect 1391 11250 1479 11309
rect 1391 11204 1420 11250
rect 1466 11204 1479 11250
rect 1391 11145 1479 11204
rect 1391 11099 1420 11145
rect 1466 11099 1479 11145
rect 1391 11040 1479 11099
rect 1391 10994 1420 11040
rect 1466 10994 1479 11040
rect 1391 10935 1479 10994
rect 1391 10889 1420 10935
rect 1466 10889 1479 10935
rect 1391 10830 1479 10889
rect 1391 10784 1420 10830
rect 1466 10784 1479 10830
rect 1391 10725 1479 10784
rect 1391 10679 1420 10725
rect 1466 10679 1479 10725
rect 1391 10620 1479 10679
rect 1391 10574 1420 10620
rect 1466 10574 1479 10620
rect 1391 10515 1479 10574
rect 1391 10469 1420 10515
rect 1466 10469 1479 10515
rect 1391 10410 1479 10469
rect 1391 10364 1420 10410
rect 1466 10364 1479 10410
rect 1391 10351 1479 10364
rect 1631 12606 1719 12619
rect 1631 12560 1644 12606
rect 1690 12560 1719 12606
rect 1631 12502 1719 12560
rect 1631 12456 1644 12502
rect 1690 12456 1719 12502
rect 1631 12398 1719 12456
rect 1631 12352 1644 12398
rect 1690 12352 1719 12398
rect 1631 12294 1719 12352
rect 1631 12248 1644 12294
rect 1690 12248 1719 12294
rect 1631 12190 1719 12248
rect 1631 12144 1644 12190
rect 1690 12144 1719 12190
rect 1631 12086 1719 12144
rect 1631 12040 1644 12086
rect 1690 12040 1719 12086
rect 1631 11982 1719 12040
rect 1631 11936 1644 11982
rect 1690 11936 1719 11982
rect 1631 11878 1719 11936
rect 1631 11832 1644 11878
rect 1690 11832 1719 11878
rect 1631 11774 1719 11832
rect 1631 11728 1644 11774
rect 1690 11728 1719 11774
rect 1631 11670 1719 11728
rect 1631 11624 1644 11670
rect 1690 11624 1719 11670
rect 1631 11565 1719 11624
rect 1631 11519 1644 11565
rect 1690 11519 1719 11565
rect 1631 11460 1719 11519
rect 1631 11414 1644 11460
rect 1690 11414 1719 11460
rect 1631 11355 1719 11414
rect 1631 11309 1644 11355
rect 1690 11309 1719 11355
rect 1631 11250 1719 11309
rect 1631 11204 1644 11250
rect 1690 11204 1719 11250
rect 1631 11145 1719 11204
rect 1631 11099 1644 11145
rect 1690 11099 1719 11145
rect 1631 11040 1719 11099
rect 1631 10994 1644 11040
rect 1690 10994 1719 11040
rect 1631 10935 1719 10994
rect 1631 10889 1644 10935
rect 1690 10889 1719 10935
rect 1631 10830 1719 10889
rect 1631 10784 1644 10830
rect 1690 10784 1719 10830
rect 1631 10725 1719 10784
rect 1631 10679 1644 10725
rect 1690 10679 1719 10725
rect 1631 10620 1719 10679
rect 1631 10574 1644 10620
rect 1690 10574 1719 10620
rect 1631 10515 1719 10574
rect 1631 10469 1644 10515
rect 1690 10469 1719 10515
rect 1631 10410 1719 10469
rect 1631 10364 1644 10410
rect 1690 10364 1719 10410
rect 1631 10351 1719 10364
rect 1839 12606 1927 12619
rect 1839 12560 1868 12606
rect 1914 12560 1927 12606
rect 1839 12502 1927 12560
rect 1839 12456 1868 12502
rect 1914 12456 1927 12502
rect 1839 12398 1927 12456
rect 1839 12352 1868 12398
rect 1914 12352 1927 12398
rect 1839 12294 1927 12352
rect 1839 12248 1868 12294
rect 1914 12248 1927 12294
rect 1839 12190 1927 12248
rect 1839 12144 1868 12190
rect 1914 12144 1927 12190
rect 1839 12086 1927 12144
rect 1839 12040 1868 12086
rect 1914 12040 1927 12086
rect 1839 11982 1927 12040
rect 1839 11936 1868 11982
rect 1914 11936 1927 11982
rect 1839 11878 1927 11936
rect 1839 11832 1868 11878
rect 1914 11832 1927 11878
rect 1839 11774 1927 11832
rect 1839 11728 1868 11774
rect 1914 11728 1927 11774
rect 1839 11670 1927 11728
rect 1839 11624 1868 11670
rect 1914 11624 1927 11670
rect 1839 11565 1927 11624
rect 1839 11519 1868 11565
rect 1914 11519 1927 11565
rect 1839 11460 1927 11519
rect 1839 11414 1868 11460
rect 1914 11414 1927 11460
rect 1839 11355 1927 11414
rect 1839 11309 1868 11355
rect 1914 11309 1927 11355
rect 1839 11250 1927 11309
rect 1839 11204 1868 11250
rect 1914 11204 1927 11250
rect 1839 11145 1927 11204
rect 1839 11099 1868 11145
rect 1914 11099 1927 11145
rect 1839 11040 1927 11099
rect 1839 10994 1868 11040
rect 1914 10994 1927 11040
rect 1839 10935 1927 10994
rect 1839 10889 1868 10935
rect 1914 10889 1927 10935
rect 1839 10830 1927 10889
rect 1839 10784 1868 10830
rect 1914 10784 1927 10830
rect 1839 10725 1927 10784
rect 1839 10679 1868 10725
rect 1914 10679 1927 10725
rect 1839 10620 1927 10679
rect 1839 10574 1868 10620
rect 1914 10574 1927 10620
rect 1839 10515 1927 10574
rect 1839 10469 1868 10515
rect 1914 10469 1927 10515
rect 1839 10410 1927 10469
rect 1839 10364 1868 10410
rect 1914 10364 1927 10410
rect 1839 10351 1927 10364
rect 2468 9984 2556 9997
rect 2468 9938 2481 9984
rect 2527 9938 2556 9984
rect 495 9898 583 9911
rect 1616 9898 1704 9911
rect 1616 9852 1629 9898
rect 1675 9852 1704 9898
rect 898 9798 986 9811
rect 898 9752 911 9798
rect 957 9752 986 9798
rect 898 9678 986 9752
rect 898 9632 911 9678
rect 957 9632 986 9678
rect 898 9619 986 9632
rect 1106 9798 1194 9811
rect 1106 9752 1135 9798
rect 1181 9752 1194 9798
rect 1106 9678 1194 9752
rect 1616 9778 1704 9852
rect 1616 9732 1629 9778
rect 1675 9732 1704 9778
rect 1616 9719 1704 9732
rect 1824 9898 1912 9911
rect 1824 9852 1853 9898
rect 1899 9852 1912 9898
rect 1824 9778 1912 9852
rect 1824 9732 1853 9778
rect 1899 9732 1912 9778
rect 1824 9719 1912 9732
rect 2468 9856 2556 9938
rect 2468 9810 2481 9856
rect 2527 9810 2556 9856
rect 2468 9729 2556 9810
rect 1106 9632 1135 9678
rect 1181 9632 1194 9678
rect 1106 9619 1194 9632
rect 2468 9683 2481 9729
rect 2527 9683 2556 9729
rect 2468 9602 2556 9683
rect 2468 9556 2481 9602
rect 2527 9556 2556 9602
rect 2468 9543 2556 9556
rect 2676 9984 2764 9997
rect 2676 9938 2705 9984
rect 2751 9938 2764 9984
rect 2676 9856 2764 9938
rect 2676 9810 2705 9856
rect 2751 9810 2764 9856
rect 2676 9729 2764 9810
rect 2676 9683 2705 9729
rect 2751 9683 2764 9729
rect 2676 9602 2764 9683
rect 2676 9556 2705 9602
rect 2751 9556 2764 9602
rect 2676 9543 2764 9556
rect 788 8157 876 8170
rect 788 8111 801 8157
rect 847 8111 876 8157
rect 788 8037 876 8111
rect 788 7991 801 8037
rect 847 7991 876 8037
rect 788 7978 876 7991
rect 996 8157 1100 8170
rect 996 8111 1025 8157
rect 1071 8111 1100 8157
rect 996 8037 1100 8111
rect 996 7991 1025 8037
rect 1071 7991 1100 8037
rect 996 7978 1100 7991
rect 1220 8157 1308 8170
rect 1220 8111 1249 8157
rect 1295 8111 1308 8157
rect 1220 8037 1308 8111
rect 1220 7991 1249 8037
rect 1295 7991 1308 8037
rect 1220 7978 1308 7991
rect 1616 8136 1704 8149
rect 1616 8090 1629 8136
rect 1675 8090 1704 8136
rect 1616 8016 1704 8090
rect 1616 7970 1629 8016
rect 1675 7970 1704 8016
rect 1616 7957 1704 7970
rect 1824 8136 1928 8149
rect 1824 8090 1853 8136
rect 1899 8090 1928 8136
rect 1824 8016 1928 8090
rect 1824 7970 1853 8016
rect 1899 7970 1928 8016
rect 1824 7957 1928 7970
rect 2048 8136 2136 8149
rect 2048 8090 2077 8136
rect 2123 8090 2136 8136
rect 2048 8016 2136 8090
rect 2048 7970 2077 8016
rect 2123 7970 2136 8016
rect 2048 7957 2136 7970
rect 5543 536 5627 555
rect 5543 208 5562 536
rect 5608 208 5627 536
rect 5543 189 5627 208
<< mvpdiff >>
rect 601 28588 769 28633
rect 601 28542 692 28588
rect 738 28542 769 28588
rect 601 28406 769 28542
rect 601 28360 692 28406
rect 738 28360 769 28406
rect 601 28225 769 28360
rect 601 28179 692 28225
rect 738 28179 769 28225
rect 601 28043 769 28179
rect 601 27997 692 28043
rect 738 27997 769 28043
rect 601 27951 769 27997
rect 889 28588 993 28633
rect 889 28542 918 28588
rect 964 28542 993 28588
rect 889 28406 993 28542
rect 889 28360 918 28406
rect 964 28360 993 28406
rect 889 28225 993 28360
rect 889 28179 918 28225
rect 964 28179 993 28225
rect 889 28043 993 28179
rect 889 27997 918 28043
rect 964 27997 993 28043
rect 889 27951 993 27997
rect 1113 28588 1389 28633
rect 1113 28542 1228 28588
rect 1274 28542 1389 28588
rect 1113 28406 1389 28542
rect 1113 28360 1228 28406
rect 1274 28360 1389 28406
rect 1113 28225 1389 28360
rect 1113 28179 1228 28225
rect 1274 28179 1389 28225
rect 1113 28043 1389 28179
rect 1113 27997 1228 28043
rect 1274 27997 1389 28043
rect 1113 27951 1389 27997
rect 1509 28588 1613 28633
rect 1509 28542 1538 28588
rect 1584 28542 1613 28588
rect 1509 28406 1613 28542
rect 1509 28360 1538 28406
rect 1584 28360 1613 28406
rect 1509 28225 1613 28360
rect 1509 28179 1538 28225
rect 1584 28179 1613 28225
rect 1509 28043 1613 28179
rect 1509 27997 1538 28043
rect 1584 27997 1613 28043
rect 1509 27951 1613 27997
rect 1733 28588 2008 28633
rect 1733 28542 1764 28588
rect 1810 28542 1931 28588
rect 1977 28542 2008 28588
rect 1733 28406 2008 28542
rect 1733 28360 1764 28406
rect 1810 28360 1931 28406
rect 1977 28360 2008 28406
rect 1733 28225 2008 28360
rect 1733 28179 1764 28225
rect 1810 28179 1931 28225
rect 1977 28179 2008 28225
rect 1733 28043 2008 28179
rect 1733 27997 1764 28043
rect 1810 27997 1931 28043
rect 1977 27997 2008 28043
rect 1733 27951 2008 27997
rect 2128 28588 2232 28633
rect 2128 28542 2157 28588
rect 2203 28542 2232 28588
rect 2128 28406 2232 28542
rect 2128 28360 2157 28406
rect 2203 28360 2232 28406
rect 2128 28225 2232 28360
rect 2128 28179 2157 28225
rect 2203 28179 2232 28225
rect 2128 28043 2232 28179
rect 2128 27997 2157 28043
rect 2203 27997 2232 28043
rect 2128 27951 2232 27997
rect 2352 28588 2628 28633
rect 2352 28542 2467 28588
rect 2513 28542 2628 28588
rect 2352 28406 2628 28542
rect 2352 28360 2467 28406
rect 2513 28360 2628 28406
rect 2352 28225 2628 28360
rect 2352 28179 2467 28225
rect 2513 28179 2628 28225
rect 2352 28043 2628 28179
rect 2352 27997 2467 28043
rect 2513 27997 2628 28043
rect 2352 27951 2628 27997
rect 2748 28588 2852 28633
rect 2748 28542 2777 28588
rect 2823 28542 2852 28588
rect 2748 28406 2852 28542
rect 2748 28360 2777 28406
rect 2823 28360 2852 28406
rect 2748 28225 2852 28360
rect 2748 28179 2777 28225
rect 2823 28179 2852 28225
rect 2748 28043 2852 28179
rect 2748 27997 2777 28043
rect 2823 27997 2852 28043
rect 2748 27951 2852 27997
rect 2972 28588 3246 28633
rect 2972 28542 3003 28588
rect 3049 28542 3169 28588
rect 3215 28542 3246 28588
rect 2972 28406 3246 28542
rect 2972 28360 3003 28406
rect 3049 28360 3169 28406
rect 3215 28360 3246 28406
rect 2972 28225 3246 28360
rect 2972 28179 3003 28225
rect 3049 28179 3169 28225
rect 3215 28179 3246 28225
rect 2972 28043 3246 28179
rect 2972 27997 3003 28043
rect 3049 27997 3169 28043
rect 3215 27997 3246 28043
rect 2972 27951 3246 27997
rect 3366 28588 3470 28633
rect 3366 28542 3395 28588
rect 3441 28542 3470 28588
rect 3366 28406 3470 28542
rect 3366 28360 3395 28406
rect 3441 28360 3470 28406
rect 3366 28225 3470 28360
rect 3366 28179 3395 28225
rect 3441 28179 3470 28225
rect 3366 28043 3470 28179
rect 3366 27997 3395 28043
rect 3441 27997 3470 28043
rect 3366 27951 3470 27997
rect 3590 28588 3866 28633
rect 3590 28542 3705 28588
rect 3751 28542 3866 28588
rect 3590 28406 3866 28542
rect 3590 28360 3705 28406
rect 3751 28360 3866 28406
rect 3590 28225 3866 28360
rect 3590 28179 3705 28225
rect 3751 28179 3866 28225
rect 3590 28043 3866 28179
rect 3590 27997 3705 28043
rect 3751 27997 3866 28043
rect 3590 27951 3866 27997
rect 3986 28588 4090 28633
rect 3986 28542 4015 28588
rect 4061 28542 4090 28588
rect 3986 28406 4090 28542
rect 3986 28360 4015 28406
rect 4061 28360 4090 28406
rect 3986 28225 4090 28360
rect 3986 28179 4015 28225
rect 4061 28179 4090 28225
rect 3986 28043 4090 28179
rect 3986 27997 4015 28043
rect 4061 27997 4090 28043
rect 3986 27951 4090 27997
rect 4210 28588 4485 28633
rect 4210 28542 4241 28588
rect 4287 28542 4408 28588
rect 4454 28542 4485 28588
rect 4210 28406 4485 28542
rect 4210 28360 4241 28406
rect 4287 28360 4408 28406
rect 4454 28360 4485 28406
rect 4210 28225 4485 28360
rect 4210 28179 4241 28225
rect 4287 28179 4408 28225
rect 4454 28179 4485 28225
rect 4210 28043 4485 28179
rect 4210 27997 4241 28043
rect 4287 27997 4408 28043
rect 4454 27997 4485 28043
rect 4210 27951 4485 27997
rect 4605 28588 4709 28633
rect 4605 28542 4634 28588
rect 4680 28542 4709 28588
rect 4605 28406 4709 28542
rect 4605 28360 4634 28406
rect 4680 28360 4709 28406
rect 4605 28225 4709 28360
rect 4605 28179 4634 28225
rect 4680 28179 4709 28225
rect 4605 28043 4709 28179
rect 4605 27997 4634 28043
rect 4680 27997 4709 28043
rect 4605 27951 4709 27997
rect 4829 28588 5069 28633
rect 4829 28542 4944 28588
rect 4990 28542 5069 28588
rect 4829 28406 5069 28542
rect 4829 28360 4944 28406
rect 4990 28360 5069 28406
rect 4829 28225 5069 28360
rect 4829 28179 4944 28225
rect 4990 28179 5069 28225
rect 4829 28043 5069 28179
rect 4829 27997 4944 28043
rect 4990 27997 5069 28043
rect 4829 27951 5069 27997
rect 5189 28588 5294 28633
rect 5189 28542 5219 28588
rect 5265 28542 5294 28588
rect 5189 28406 5294 28542
rect 5189 28360 5219 28406
rect 5265 28360 5294 28406
rect 5189 28225 5294 28360
rect 5189 28179 5219 28225
rect 5265 28179 5294 28225
rect 5189 28043 5294 28179
rect 5189 27997 5219 28043
rect 5265 27997 5294 28043
rect 5189 27951 5294 27997
rect 5414 28588 5618 28633
rect 5414 28542 5480 28588
rect 5526 28542 5618 28588
rect 5414 28406 5618 28542
rect 5414 28360 5480 28406
rect 5526 28360 5618 28406
rect 5414 28225 5618 28360
rect 5414 28179 5480 28225
rect 5526 28179 5618 28225
rect 5414 28043 5618 28179
rect 5414 27997 5480 28043
rect 5526 27997 5618 28043
rect 5414 27951 5618 27997
rect 601 27812 769 27858
rect 601 27766 692 27812
rect 738 27766 769 27812
rect 601 27631 769 27766
rect 601 27585 692 27631
rect 738 27585 769 27631
rect 601 27450 769 27585
rect 601 27404 692 27450
rect 738 27404 769 27450
rect 601 27268 769 27404
rect 601 27222 692 27268
rect 738 27222 769 27268
rect 601 27176 769 27222
rect 889 27812 993 27858
rect 889 27766 918 27812
rect 964 27766 993 27812
rect 889 27631 993 27766
rect 889 27585 918 27631
rect 964 27585 993 27631
rect 889 27450 993 27585
rect 889 27404 918 27450
rect 964 27404 993 27450
rect 889 27268 993 27404
rect 889 27222 918 27268
rect 964 27222 993 27268
rect 889 27176 993 27222
rect 1113 27812 1389 27858
rect 1113 27766 1228 27812
rect 1274 27766 1389 27812
rect 1113 27631 1389 27766
rect 1113 27585 1228 27631
rect 1274 27585 1389 27631
rect 1113 27450 1389 27585
rect 1113 27404 1228 27450
rect 1274 27404 1389 27450
rect 1113 27268 1389 27404
rect 1113 27222 1228 27268
rect 1274 27222 1389 27268
rect 1113 27176 1389 27222
rect 1509 27812 1613 27858
rect 1509 27766 1538 27812
rect 1584 27766 1613 27812
rect 1509 27631 1613 27766
rect 1509 27585 1538 27631
rect 1584 27585 1613 27631
rect 1509 27450 1613 27585
rect 1509 27404 1538 27450
rect 1584 27404 1613 27450
rect 1509 27268 1613 27404
rect 1509 27222 1538 27268
rect 1584 27222 1613 27268
rect 1509 27176 1613 27222
rect 1733 27812 2008 27858
rect 1733 27766 1764 27812
rect 1810 27766 1931 27812
rect 1977 27766 2008 27812
rect 1733 27631 2008 27766
rect 1733 27585 1764 27631
rect 1810 27585 1931 27631
rect 1977 27585 2008 27631
rect 1733 27450 2008 27585
rect 1733 27404 1764 27450
rect 1810 27404 1931 27450
rect 1977 27404 2008 27450
rect 1733 27268 2008 27404
rect 1733 27222 1764 27268
rect 1810 27222 1931 27268
rect 1977 27222 2008 27268
rect 1733 27176 2008 27222
rect 2128 27812 2232 27858
rect 2128 27766 2157 27812
rect 2203 27766 2232 27812
rect 2128 27631 2232 27766
rect 2128 27585 2157 27631
rect 2203 27585 2232 27631
rect 2128 27450 2232 27585
rect 2128 27404 2157 27450
rect 2203 27404 2232 27450
rect 2128 27268 2232 27404
rect 2128 27222 2157 27268
rect 2203 27222 2232 27268
rect 2128 27176 2232 27222
rect 2352 27812 2628 27858
rect 2352 27766 2467 27812
rect 2513 27766 2628 27812
rect 2352 27631 2628 27766
rect 2352 27585 2467 27631
rect 2513 27585 2628 27631
rect 2352 27450 2628 27585
rect 2352 27404 2467 27450
rect 2513 27404 2628 27450
rect 2352 27268 2628 27404
rect 2352 27222 2467 27268
rect 2513 27222 2628 27268
rect 2352 27176 2628 27222
rect 2748 27812 2852 27858
rect 2748 27766 2777 27812
rect 2823 27766 2852 27812
rect 2748 27631 2852 27766
rect 2748 27585 2777 27631
rect 2823 27585 2852 27631
rect 2748 27450 2852 27585
rect 2748 27404 2777 27450
rect 2823 27404 2852 27450
rect 2748 27268 2852 27404
rect 2748 27222 2777 27268
rect 2823 27222 2852 27268
rect 2748 27176 2852 27222
rect 2972 27812 3246 27858
rect 2972 27766 3003 27812
rect 3049 27766 3169 27812
rect 3215 27766 3246 27812
rect 2972 27631 3246 27766
rect 2972 27585 3003 27631
rect 3049 27585 3169 27631
rect 3215 27585 3246 27631
rect 2972 27450 3246 27585
rect 2972 27404 3003 27450
rect 3049 27404 3169 27450
rect 3215 27404 3246 27450
rect 2972 27268 3246 27404
rect 2972 27222 3003 27268
rect 3049 27222 3169 27268
rect 3215 27222 3246 27268
rect 2972 27176 3246 27222
rect 3366 27812 3470 27858
rect 3366 27766 3395 27812
rect 3441 27766 3470 27812
rect 3366 27631 3470 27766
rect 3366 27585 3395 27631
rect 3441 27585 3470 27631
rect 3366 27450 3470 27585
rect 3366 27404 3395 27450
rect 3441 27404 3470 27450
rect 3366 27268 3470 27404
rect 3366 27222 3395 27268
rect 3441 27222 3470 27268
rect 3366 27176 3470 27222
rect 3590 27812 3866 27858
rect 3590 27766 3705 27812
rect 3751 27766 3866 27812
rect 3590 27631 3866 27766
rect 3590 27585 3705 27631
rect 3751 27585 3866 27631
rect 3590 27450 3866 27585
rect 3590 27404 3705 27450
rect 3751 27404 3866 27450
rect 3590 27268 3866 27404
rect 3590 27222 3705 27268
rect 3751 27222 3866 27268
rect 3590 27176 3866 27222
rect 3986 27812 4090 27858
rect 3986 27766 4015 27812
rect 4061 27766 4090 27812
rect 3986 27631 4090 27766
rect 3986 27585 4015 27631
rect 4061 27585 4090 27631
rect 3986 27450 4090 27585
rect 3986 27404 4015 27450
rect 4061 27404 4090 27450
rect 3986 27268 4090 27404
rect 3986 27222 4015 27268
rect 4061 27222 4090 27268
rect 3986 27176 4090 27222
rect 4210 27812 4485 27858
rect 4210 27766 4241 27812
rect 4287 27766 4408 27812
rect 4454 27766 4485 27812
rect 4210 27631 4485 27766
rect 4210 27585 4241 27631
rect 4287 27585 4408 27631
rect 4454 27585 4485 27631
rect 4210 27450 4485 27585
rect 4210 27404 4241 27450
rect 4287 27404 4408 27450
rect 4454 27404 4485 27450
rect 4210 27268 4485 27404
rect 4210 27222 4241 27268
rect 4287 27222 4408 27268
rect 4454 27222 4485 27268
rect 4210 27176 4485 27222
rect 4605 27812 4709 27858
rect 4605 27766 4634 27812
rect 4680 27766 4709 27812
rect 4605 27631 4709 27766
rect 4605 27585 4634 27631
rect 4680 27585 4709 27631
rect 4605 27450 4709 27585
rect 4605 27404 4634 27450
rect 4680 27404 4709 27450
rect 4605 27268 4709 27404
rect 4605 27222 4634 27268
rect 4680 27222 4709 27268
rect 4605 27176 4709 27222
rect 4829 27812 5069 27858
rect 4829 27766 4944 27812
rect 4990 27766 5069 27812
rect 4829 27631 5069 27766
rect 4829 27585 4944 27631
rect 4990 27585 5069 27631
rect 4829 27450 5069 27585
rect 4829 27404 4944 27450
rect 4990 27404 5069 27450
rect 4829 27268 5069 27404
rect 4829 27222 4944 27268
rect 4990 27222 5069 27268
rect 4829 27176 5069 27222
rect 5189 27812 5294 27858
rect 5189 27766 5219 27812
rect 5265 27766 5294 27812
rect 5189 27631 5294 27766
rect 5189 27585 5219 27631
rect 5265 27585 5294 27631
rect 5189 27450 5294 27585
rect 5189 27404 5219 27450
rect 5265 27404 5294 27450
rect 5189 27268 5294 27404
rect 5189 27222 5219 27268
rect 5265 27222 5294 27268
rect 5189 27176 5294 27222
rect 5414 27812 5618 27858
rect 5414 27766 5480 27812
rect 5526 27766 5618 27812
rect 5414 27631 5618 27766
rect 5414 27585 5480 27631
rect 5526 27585 5618 27631
rect 5414 27450 5618 27585
rect 5414 27404 5480 27450
rect 5526 27404 5618 27450
rect 5414 27268 5618 27404
rect 5414 27222 5480 27268
rect 5526 27222 5618 27268
rect 5414 27176 5618 27222
rect 795 26944 883 26957
rect 795 26898 808 26944
rect 854 26898 883 26944
rect 795 26836 883 26898
rect 795 26790 808 26836
rect 854 26790 883 26836
rect 795 26728 883 26790
rect 795 26682 808 26728
rect 854 26682 883 26728
rect 795 26620 883 26682
rect 795 26574 808 26620
rect 854 26574 883 26620
rect 795 26512 883 26574
rect 795 26466 808 26512
rect 854 26466 883 26512
rect 795 26404 883 26466
rect 795 26358 808 26404
rect 854 26358 883 26404
rect 795 26296 883 26358
rect 795 26250 808 26296
rect 854 26250 883 26296
rect 795 26189 883 26250
rect 795 26143 808 26189
rect 854 26143 883 26189
rect 795 26082 883 26143
rect 795 26036 808 26082
rect 854 26036 883 26082
rect 795 25975 883 26036
rect 795 25929 808 25975
rect 854 25929 883 25975
rect 795 25868 883 25929
rect 795 25822 808 25868
rect 854 25822 883 25868
rect 795 25761 883 25822
rect 795 25715 808 25761
rect 854 25715 883 25761
rect 795 25654 883 25715
rect 795 25608 808 25654
rect 854 25608 883 25654
rect 795 25595 883 25608
rect 1003 26944 1091 26957
rect 1003 26898 1032 26944
rect 1078 26898 1091 26944
rect 1003 26836 1091 26898
rect 1003 26790 1032 26836
rect 1078 26790 1091 26836
rect 1003 26728 1091 26790
rect 1003 26682 1032 26728
rect 1078 26682 1091 26728
rect 1003 26620 1091 26682
rect 1003 26574 1032 26620
rect 1078 26574 1091 26620
rect 1003 26512 1091 26574
rect 1003 26466 1032 26512
rect 1078 26466 1091 26512
rect 1003 26404 1091 26466
rect 1003 26358 1032 26404
rect 1078 26358 1091 26404
rect 1003 26296 1091 26358
rect 1003 26250 1032 26296
rect 1078 26250 1091 26296
rect 1003 26189 1091 26250
rect 1003 26143 1032 26189
rect 1078 26143 1091 26189
rect 1003 26082 1091 26143
rect 1003 26036 1032 26082
rect 1078 26036 1091 26082
rect 1003 25975 1091 26036
rect 1003 25929 1032 25975
rect 1078 25929 1091 25975
rect 1003 25868 1091 25929
rect 1003 25822 1032 25868
rect 1078 25822 1091 25868
rect 1003 25761 1091 25822
rect 1003 25715 1032 25761
rect 1078 25715 1091 25761
rect 1003 25654 1091 25715
rect 1003 25608 1032 25654
rect 1078 25608 1091 25654
rect 1003 25595 1091 25608
rect 1411 26944 1499 26957
rect 1411 26898 1424 26944
rect 1470 26898 1499 26944
rect 1411 26836 1499 26898
rect 1411 26790 1424 26836
rect 1470 26790 1499 26836
rect 1411 26728 1499 26790
rect 1411 26682 1424 26728
rect 1470 26682 1499 26728
rect 1411 26620 1499 26682
rect 1411 26574 1424 26620
rect 1470 26574 1499 26620
rect 1411 26512 1499 26574
rect 1411 26466 1424 26512
rect 1470 26466 1499 26512
rect 1411 26404 1499 26466
rect 1411 26358 1424 26404
rect 1470 26358 1499 26404
rect 1411 26296 1499 26358
rect 1411 26250 1424 26296
rect 1470 26250 1499 26296
rect 1411 26189 1499 26250
rect 1411 26143 1424 26189
rect 1470 26143 1499 26189
rect 1411 26082 1499 26143
rect 1411 26036 1424 26082
rect 1470 26036 1499 26082
rect 1411 25975 1499 26036
rect 1411 25929 1424 25975
rect 1470 25929 1499 25975
rect 1411 25868 1499 25929
rect 1411 25822 1424 25868
rect 1470 25822 1499 25868
rect 1411 25761 1499 25822
rect 1411 25715 1424 25761
rect 1470 25715 1499 25761
rect 1411 25654 1499 25715
rect 1411 25608 1424 25654
rect 1470 25608 1499 25654
rect 1411 25595 1499 25608
rect 1619 26944 1707 26957
rect 1619 26898 1648 26944
rect 1694 26898 1707 26944
rect 1619 26836 1707 26898
rect 1619 26790 1648 26836
rect 1694 26790 1707 26836
rect 1619 26728 1707 26790
rect 1619 26682 1648 26728
rect 1694 26682 1707 26728
rect 1619 26620 1707 26682
rect 1619 26574 1648 26620
rect 1694 26574 1707 26620
rect 1619 26512 1707 26574
rect 1619 26466 1648 26512
rect 1694 26466 1707 26512
rect 1619 26404 1707 26466
rect 1619 26358 1648 26404
rect 1694 26358 1707 26404
rect 1619 26296 1707 26358
rect 1619 26250 1648 26296
rect 1694 26250 1707 26296
rect 1619 26189 1707 26250
rect 1619 26143 1648 26189
rect 1694 26143 1707 26189
rect 1619 26082 1707 26143
rect 1619 26036 1648 26082
rect 1694 26036 1707 26082
rect 1619 25975 1707 26036
rect 1619 25929 1648 25975
rect 1694 25929 1707 25975
rect 1619 25868 1707 25929
rect 1619 25822 1648 25868
rect 1694 25822 1707 25868
rect 1619 25761 1707 25822
rect 1619 25715 1648 25761
rect 1694 25715 1707 25761
rect 1619 25654 1707 25715
rect 1619 25608 1648 25654
rect 1694 25608 1707 25654
rect 1619 25595 1707 25608
rect 2034 26944 2122 26957
rect 2034 26898 2047 26944
rect 2093 26898 2122 26944
rect 2034 26836 2122 26898
rect 2034 26790 2047 26836
rect 2093 26790 2122 26836
rect 2034 26728 2122 26790
rect 2034 26682 2047 26728
rect 2093 26682 2122 26728
rect 2034 26620 2122 26682
rect 2034 26574 2047 26620
rect 2093 26574 2122 26620
rect 2034 26512 2122 26574
rect 2034 26466 2047 26512
rect 2093 26466 2122 26512
rect 2034 26404 2122 26466
rect 2034 26358 2047 26404
rect 2093 26358 2122 26404
rect 2034 26296 2122 26358
rect 2034 26250 2047 26296
rect 2093 26250 2122 26296
rect 2034 26189 2122 26250
rect 2034 26143 2047 26189
rect 2093 26143 2122 26189
rect 2034 26082 2122 26143
rect 2034 26036 2047 26082
rect 2093 26036 2122 26082
rect 2034 25975 2122 26036
rect 2034 25929 2047 25975
rect 2093 25929 2122 25975
rect 2034 25868 2122 25929
rect 2034 25822 2047 25868
rect 2093 25822 2122 25868
rect 2034 25761 2122 25822
rect 2034 25715 2047 25761
rect 2093 25715 2122 25761
rect 2034 25654 2122 25715
rect 2034 25608 2047 25654
rect 2093 25608 2122 25654
rect 2034 25595 2122 25608
rect 2242 26944 2330 26957
rect 2242 26898 2271 26944
rect 2317 26898 2330 26944
rect 2242 26836 2330 26898
rect 2242 26790 2271 26836
rect 2317 26790 2330 26836
rect 2242 26728 2330 26790
rect 2242 26682 2271 26728
rect 2317 26682 2330 26728
rect 2242 26620 2330 26682
rect 2242 26574 2271 26620
rect 2317 26574 2330 26620
rect 2242 26512 2330 26574
rect 2242 26466 2271 26512
rect 2317 26466 2330 26512
rect 2242 26404 2330 26466
rect 2242 26358 2271 26404
rect 2317 26358 2330 26404
rect 2242 26296 2330 26358
rect 2242 26250 2271 26296
rect 2317 26250 2330 26296
rect 2242 26189 2330 26250
rect 2242 26143 2271 26189
rect 2317 26143 2330 26189
rect 2242 26082 2330 26143
rect 2242 26036 2271 26082
rect 2317 26036 2330 26082
rect 2242 25975 2330 26036
rect 2242 25929 2271 25975
rect 2317 25929 2330 25975
rect 2242 25868 2330 25929
rect 2242 25822 2271 25868
rect 2317 25822 2330 25868
rect 2242 25761 2330 25822
rect 2242 25715 2271 25761
rect 2317 25715 2330 25761
rect 2242 25654 2330 25715
rect 2242 25608 2271 25654
rect 2317 25608 2330 25654
rect 2242 25595 2330 25608
rect 2650 26944 2738 26957
rect 2650 26898 2663 26944
rect 2709 26898 2738 26944
rect 2650 26836 2738 26898
rect 2650 26790 2663 26836
rect 2709 26790 2738 26836
rect 2650 26728 2738 26790
rect 2650 26682 2663 26728
rect 2709 26682 2738 26728
rect 2650 26620 2738 26682
rect 2650 26574 2663 26620
rect 2709 26574 2738 26620
rect 2650 26512 2738 26574
rect 2650 26466 2663 26512
rect 2709 26466 2738 26512
rect 2650 26404 2738 26466
rect 2650 26358 2663 26404
rect 2709 26358 2738 26404
rect 2650 26296 2738 26358
rect 2650 26250 2663 26296
rect 2709 26250 2738 26296
rect 2650 26189 2738 26250
rect 2650 26143 2663 26189
rect 2709 26143 2738 26189
rect 2650 26082 2738 26143
rect 2650 26036 2663 26082
rect 2709 26036 2738 26082
rect 2650 25975 2738 26036
rect 2650 25929 2663 25975
rect 2709 25929 2738 25975
rect 2650 25868 2738 25929
rect 2650 25822 2663 25868
rect 2709 25822 2738 25868
rect 2650 25761 2738 25822
rect 2650 25715 2663 25761
rect 2709 25715 2738 25761
rect 2650 25654 2738 25715
rect 2650 25608 2663 25654
rect 2709 25608 2738 25654
rect 2650 25595 2738 25608
rect 2858 26944 2946 26957
rect 2858 26898 2887 26944
rect 2933 26898 2946 26944
rect 2858 26836 2946 26898
rect 2858 26790 2887 26836
rect 2933 26790 2946 26836
rect 2858 26728 2946 26790
rect 2858 26682 2887 26728
rect 2933 26682 2946 26728
rect 2858 26620 2946 26682
rect 2858 26574 2887 26620
rect 2933 26574 2946 26620
rect 2858 26512 2946 26574
rect 2858 26466 2887 26512
rect 2933 26466 2946 26512
rect 2858 26404 2946 26466
rect 2858 26358 2887 26404
rect 2933 26358 2946 26404
rect 2858 26296 2946 26358
rect 2858 26250 2887 26296
rect 2933 26250 2946 26296
rect 2858 26189 2946 26250
rect 2858 26143 2887 26189
rect 2933 26143 2946 26189
rect 2858 26082 2946 26143
rect 2858 26036 2887 26082
rect 2933 26036 2946 26082
rect 2858 25975 2946 26036
rect 2858 25929 2887 25975
rect 2933 25929 2946 25975
rect 2858 25868 2946 25929
rect 2858 25822 2887 25868
rect 2933 25822 2946 25868
rect 2858 25761 2946 25822
rect 2858 25715 2887 25761
rect 2933 25715 2946 25761
rect 2858 25654 2946 25715
rect 2858 25608 2887 25654
rect 2933 25608 2946 25654
rect 2858 25595 2946 25608
rect 3272 26944 3360 26957
rect 3272 26898 3285 26944
rect 3331 26898 3360 26944
rect 3272 26836 3360 26898
rect 3272 26790 3285 26836
rect 3331 26790 3360 26836
rect 3272 26728 3360 26790
rect 3272 26682 3285 26728
rect 3331 26682 3360 26728
rect 3272 26620 3360 26682
rect 3272 26574 3285 26620
rect 3331 26574 3360 26620
rect 3272 26512 3360 26574
rect 3272 26466 3285 26512
rect 3331 26466 3360 26512
rect 3272 26404 3360 26466
rect 3272 26358 3285 26404
rect 3331 26358 3360 26404
rect 3272 26296 3360 26358
rect 3272 26250 3285 26296
rect 3331 26250 3360 26296
rect 3272 26189 3360 26250
rect 3272 26143 3285 26189
rect 3331 26143 3360 26189
rect 3272 26082 3360 26143
rect 3272 26036 3285 26082
rect 3331 26036 3360 26082
rect 3272 25975 3360 26036
rect 3272 25929 3285 25975
rect 3331 25929 3360 25975
rect 3272 25868 3360 25929
rect 3272 25822 3285 25868
rect 3331 25822 3360 25868
rect 3272 25761 3360 25822
rect 3272 25715 3285 25761
rect 3331 25715 3360 25761
rect 3272 25654 3360 25715
rect 3272 25608 3285 25654
rect 3331 25608 3360 25654
rect 3272 25595 3360 25608
rect 3480 26944 3568 26957
rect 3480 26898 3509 26944
rect 3555 26898 3568 26944
rect 3480 26836 3568 26898
rect 3480 26790 3509 26836
rect 3555 26790 3568 26836
rect 3480 26728 3568 26790
rect 3480 26682 3509 26728
rect 3555 26682 3568 26728
rect 3480 26620 3568 26682
rect 3480 26574 3509 26620
rect 3555 26574 3568 26620
rect 3480 26512 3568 26574
rect 3480 26466 3509 26512
rect 3555 26466 3568 26512
rect 3480 26404 3568 26466
rect 3480 26358 3509 26404
rect 3555 26358 3568 26404
rect 3480 26296 3568 26358
rect 3480 26250 3509 26296
rect 3555 26250 3568 26296
rect 3480 26189 3568 26250
rect 3480 26143 3509 26189
rect 3555 26143 3568 26189
rect 3480 26082 3568 26143
rect 3480 26036 3509 26082
rect 3555 26036 3568 26082
rect 3480 25975 3568 26036
rect 3480 25929 3509 25975
rect 3555 25929 3568 25975
rect 3480 25868 3568 25929
rect 3480 25822 3509 25868
rect 3555 25822 3568 25868
rect 3480 25761 3568 25822
rect 3480 25715 3509 25761
rect 3555 25715 3568 25761
rect 3480 25654 3568 25715
rect 3480 25608 3509 25654
rect 3555 25608 3568 25654
rect 3480 25595 3568 25608
rect 3888 26944 3976 26957
rect 3888 26898 3901 26944
rect 3947 26898 3976 26944
rect 3888 26836 3976 26898
rect 3888 26790 3901 26836
rect 3947 26790 3976 26836
rect 3888 26728 3976 26790
rect 3888 26682 3901 26728
rect 3947 26682 3976 26728
rect 3888 26620 3976 26682
rect 3888 26574 3901 26620
rect 3947 26574 3976 26620
rect 3888 26512 3976 26574
rect 3888 26466 3901 26512
rect 3947 26466 3976 26512
rect 3888 26404 3976 26466
rect 3888 26358 3901 26404
rect 3947 26358 3976 26404
rect 3888 26296 3976 26358
rect 3888 26250 3901 26296
rect 3947 26250 3976 26296
rect 3888 26189 3976 26250
rect 3888 26143 3901 26189
rect 3947 26143 3976 26189
rect 3888 26082 3976 26143
rect 3888 26036 3901 26082
rect 3947 26036 3976 26082
rect 3888 25975 3976 26036
rect 3888 25929 3901 25975
rect 3947 25929 3976 25975
rect 3888 25868 3976 25929
rect 3888 25822 3901 25868
rect 3947 25822 3976 25868
rect 3888 25761 3976 25822
rect 3888 25715 3901 25761
rect 3947 25715 3976 25761
rect 3888 25654 3976 25715
rect 3888 25608 3901 25654
rect 3947 25608 3976 25654
rect 3888 25595 3976 25608
rect 4096 26944 4184 26957
rect 4096 26898 4125 26944
rect 4171 26898 4184 26944
rect 4096 26836 4184 26898
rect 4096 26790 4125 26836
rect 4171 26790 4184 26836
rect 4096 26728 4184 26790
rect 4096 26682 4125 26728
rect 4171 26682 4184 26728
rect 4096 26620 4184 26682
rect 4096 26574 4125 26620
rect 4171 26574 4184 26620
rect 4096 26512 4184 26574
rect 4096 26466 4125 26512
rect 4171 26466 4184 26512
rect 4096 26404 4184 26466
rect 4096 26358 4125 26404
rect 4171 26358 4184 26404
rect 4096 26296 4184 26358
rect 4096 26250 4125 26296
rect 4171 26250 4184 26296
rect 4096 26189 4184 26250
rect 4096 26143 4125 26189
rect 4171 26143 4184 26189
rect 4096 26082 4184 26143
rect 4096 26036 4125 26082
rect 4171 26036 4184 26082
rect 4096 25975 4184 26036
rect 4096 25929 4125 25975
rect 4171 25929 4184 25975
rect 4096 25868 4184 25929
rect 4096 25822 4125 25868
rect 4171 25822 4184 25868
rect 4096 25761 4184 25822
rect 4096 25715 4125 25761
rect 4171 25715 4184 25761
rect 4096 25654 4184 25715
rect 4096 25608 4125 25654
rect 4171 25608 4184 25654
rect 4096 25595 4184 25608
rect 4511 26944 4599 26957
rect 4511 26898 4524 26944
rect 4570 26898 4599 26944
rect 4511 26836 4599 26898
rect 4511 26790 4524 26836
rect 4570 26790 4599 26836
rect 4511 26728 4599 26790
rect 4511 26682 4524 26728
rect 4570 26682 4599 26728
rect 4511 26620 4599 26682
rect 4511 26574 4524 26620
rect 4570 26574 4599 26620
rect 4511 26512 4599 26574
rect 4511 26466 4524 26512
rect 4570 26466 4599 26512
rect 4511 26404 4599 26466
rect 4511 26358 4524 26404
rect 4570 26358 4599 26404
rect 4511 26296 4599 26358
rect 4511 26250 4524 26296
rect 4570 26250 4599 26296
rect 4511 26189 4599 26250
rect 4511 26143 4524 26189
rect 4570 26143 4599 26189
rect 4511 26082 4599 26143
rect 4511 26036 4524 26082
rect 4570 26036 4599 26082
rect 4511 25975 4599 26036
rect 4511 25929 4524 25975
rect 4570 25929 4599 25975
rect 4511 25868 4599 25929
rect 4511 25822 4524 25868
rect 4570 25822 4599 25868
rect 4511 25761 4599 25822
rect 4511 25715 4524 25761
rect 4570 25715 4599 25761
rect 4511 25654 4599 25715
rect 4511 25608 4524 25654
rect 4570 25608 4599 25654
rect 4511 25595 4599 25608
rect 4719 26944 4807 26957
rect 4719 26898 4748 26944
rect 4794 26898 4807 26944
rect 4719 26836 4807 26898
rect 4719 26790 4748 26836
rect 4794 26790 4807 26836
rect 4719 26728 4807 26790
rect 4719 26682 4748 26728
rect 4794 26682 4807 26728
rect 4719 26620 4807 26682
rect 4719 26574 4748 26620
rect 4794 26574 4807 26620
rect 4719 26512 4807 26574
rect 4719 26466 4748 26512
rect 4794 26466 4807 26512
rect 4719 26404 4807 26466
rect 4719 26358 4748 26404
rect 4794 26358 4807 26404
rect 4719 26296 4807 26358
rect 4719 26250 4748 26296
rect 4794 26250 4807 26296
rect 4719 26189 4807 26250
rect 4719 26143 4748 26189
rect 4794 26143 4807 26189
rect 4719 26082 4807 26143
rect 4719 26036 4748 26082
rect 4794 26036 4807 26082
rect 4719 25975 4807 26036
rect 4719 25929 4748 25975
rect 4794 25929 4807 25975
rect 4719 25868 4807 25929
rect 4719 25822 4748 25868
rect 4794 25822 4807 25868
rect 4719 25761 4807 25822
rect 4719 25715 4748 25761
rect 4794 25715 4807 25761
rect 4719 25654 4807 25715
rect 4719 25608 4748 25654
rect 4794 25608 4807 25654
rect 4719 25595 4807 25608
rect 5127 26944 5215 26957
rect 5127 26898 5140 26944
rect 5186 26898 5215 26944
rect 5127 26836 5215 26898
rect 5127 26790 5140 26836
rect 5186 26790 5215 26836
rect 5127 26728 5215 26790
rect 5127 26682 5140 26728
rect 5186 26682 5215 26728
rect 5127 26620 5215 26682
rect 5127 26574 5140 26620
rect 5186 26574 5215 26620
rect 5127 26512 5215 26574
rect 5127 26466 5140 26512
rect 5186 26466 5215 26512
rect 5127 26404 5215 26466
rect 5127 26358 5140 26404
rect 5186 26358 5215 26404
rect 5127 26296 5215 26358
rect 5127 26250 5140 26296
rect 5186 26250 5215 26296
rect 5127 26189 5215 26250
rect 5127 26143 5140 26189
rect 5186 26143 5215 26189
rect 5127 26082 5215 26143
rect 5127 26036 5140 26082
rect 5186 26036 5215 26082
rect 5127 25975 5215 26036
rect 5127 25929 5140 25975
rect 5186 25929 5215 25975
rect 5127 25868 5215 25929
rect 5127 25822 5140 25868
rect 5186 25822 5215 25868
rect 5127 25761 5215 25822
rect 5127 25715 5140 25761
rect 5186 25715 5215 25761
rect 5127 25654 5215 25715
rect 5127 25608 5140 25654
rect 5186 25608 5215 25654
rect 5127 25595 5215 25608
rect 5335 26944 5423 26957
rect 5335 26898 5364 26944
rect 5410 26898 5423 26944
rect 5335 26836 5423 26898
rect 5335 26790 5364 26836
rect 5410 26790 5423 26836
rect 5335 26728 5423 26790
rect 5335 26682 5364 26728
rect 5410 26682 5423 26728
rect 5335 26620 5423 26682
rect 5335 26574 5364 26620
rect 5410 26574 5423 26620
rect 5335 26512 5423 26574
rect 5335 26466 5364 26512
rect 5410 26466 5423 26512
rect 5335 26404 5423 26466
rect 5335 26358 5364 26404
rect 5410 26358 5423 26404
rect 5335 26296 5423 26358
rect 5335 26250 5364 26296
rect 5410 26250 5423 26296
rect 5335 26189 5423 26250
rect 5335 26143 5364 26189
rect 5410 26143 5423 26189
rect 5335 26082 5423 26143
rect 5335 26036 5364 26082
rect 5410 26036 5423 26082
rect 5335 25975 5423 26036
rect 5335 25929 5364 25975
rect 5410 25929 5423 25975
rect 5335 25868 5423 25929
rect 5335 25822 5364 25868
rect 5410 25822 5423 25868
rect 5335 25761 5423 25822
rect 5335 25715 5364 25761
rect 5410 25715 5423 25761
rect 5335 25654 5423 25715
rect 5335 25608 5364 25654
rect 5410 25608 5423 25654
rect 5335 25595 5423 25608
rect 793 25357 881 25370
rect 793 25311 806 25357
rect 852 25311 881 25357
rect 793 25249 881 25311
rect 793 25203 806 25249
rect 852 25203 881 25249
rect 793 25141 881 25203
rect 793 25095 806 25141
rect 852 25095 881 25141
rect 793 25033 881 25095
rect 793 24987 806 25033
rect 852 24987 881 25033
rect 793 24925 881 24987
rect 793 24879 806 24925
rect 852 24879 881 24925
rect 793 24817 881 24879
rect 793 24771 806 24817
rect 852 24771 881 24817
rect 793 24709 881 24771
rect 793 24663 806 24709
rect 852 24663 881 24709
rect 793 24602 881 24663
rect 793 24556 806 24602
rect 852 24556 881 24602
rect 793 24495 881 24556
rect 793 24449 806 24495
rect 852 24449 881 24495
rect 793 24388 881 24449
rect 793 24342 806 24388
rect 852 24342 881 24388
rect 793 24281 881 24342
rect 793 24235 806 24281
rect 852 24235 881 24281
rect 793 24174 881 24235
rect 793 24128 806 24174
rect 852 24128 881 24174
rect 793 24067 881 24128
rect 793 24021 806 24067
rect 852 24021 881 24067
rect 793 24008 881 24021
rect 1001 25357 1089 25370
rect 1001 25311 1030 25357
rect 1076 25311 1089 25357
rect 1001 25249 1089 25311
rect 1001 25203 1030 25249
rect 1076 25203 1089 25249
rect 1001 25141 1089 25203
rect 1001 25095 1030 25141
rect 1076 25095 1089 25141
rect 1001 25033 1089 25095
rect 1001 24987 1030 25033
rect 1076 24987 1089 25033
rect 1001 24925 1089 24987
rect 1001 24879 1030 24925
rect 1076 24879 1089 24925
rect 1001 24817 1089 24879
rect 1001 24771 1030 24817
rect 1076 24771 1089 24817
rect 1001 24709 1089 24771
rect 1001 24663 1030 24709
rect 1076 24663 1089 24709
rect 1413 25357 1501 25370
rect 1413 25311 1426 25357
rect 1472 25311 1501 25357
rect 1413 25249 1501 25311
rect 1413 25203 1426 25249
rect 1472 25203 1501 25249
rect 1413 25141 1501 25203
rect 1413 25095 1426 25141
rect 1472 25095 1501 25141
rect 1413 25033 1501 25095
rect 1413 24987 1426 25033
rect 1472 24987 1501 25033
rect 1413 24925 1501 24987
rect 1413 24879 1426 24925
rect 1472 24879 1501 24925
rect 1413 24817 1501 24879
rect 1413 24771 1426 24817
rect 1472 24771 1501 24817
rect 1413 24709 1501 24771
rect 1001 24602 1089 24663
rect 1001 24556 1030 24602
rect 1076 24556 1089 24602
rect 1001 24495 1089 24556
rect 1001 24449 1030 24495
rect 1076 24449 1089 24495
rect 1001 24388 1089 24449
rect 1413 24663 1426 24709
rect 1472 24663 1501 24709
rect 1413 24602 1501 24663
rect 1413 24556 1426 24602
rect 1472 24556 1501 24602
rect 1413 24495 1501 24556
rect 1413 24449 1426 24495
rect 1472 24449 1501 24495
rect 1001 24342 1030 24388
rect 1076 24342 1089 24388
rect 1001 24281 1089 24342
rect 1001 24235 1030 24281
rect 1076 24235 1089 24281
rect 1001 24174 1089 24235
rect 1001 24128 1030 24174
rect 1076 24128 1089 24174
rect 1001 24067 1089 24128
rect 1001 24021 1030 24067
rect 1076 24021 1089 24067
rect 1001 24008 1089 24021
rect 1413 24388 1501 24449
rect 1413 24342 1426 24388
rect 1472 24342 1501 24388
rect 1413 24281 1501 24342
rect 1413 24235 1426 24281
rect 1472 24235 1501 24281
rect 1413 24174 1501 24235
rect 1413 24128 1426 24174
rect 1472 24128 1501 24174
rect 1413 24067 1501 24128
rect 1413 24021 1426 24067
rect 1472 24021 1501 24067
rect 1413 24008 1501 24021
rect 1621 25357 1709 25370
rect 1621 25311 1650 25357
rect 1696 25311 1709 25357
rect 1621 25249 1709 25311
rect 1621 25203 1650 25249
rect 1696 25203 1709 25249
rect 1621 25141 1709 25203
rect 1621 25095 1650 25141
rect 1696 25095 1709 25141
rect 1621 25033 1709 25095
rect 1621 24987 1650 25033
rect 1696 24987 1709 25033
rect 1621 24925 1709 24987
rect 1621 24879 1650 24925
rect 1696 24879 1709 24925
rect 1621 24817 1709 24879
rect 1621 24771 1650 24817
rect 1696 24771 1709 24817
rect 1621 24709 1709 24771
rect 1621 24663 1650 24709
rect 1696 24663 1709 24709
rect 1621 24602 1709 24663
rect 1621 24556 1650 24602
rect 1696 24556 1709 24602
rect 1621 24495 1709 24556
rect 1621 24449 1650 24495
rect 1696 24449 1709 24495
rect 1621 24388 1709 24449
rect 1621 24342 1650 24388
rect 1696 24342 1709 24388
rect 1621 24281 1709 24342
rect 1621 24235 1650 24281
rect 1696 24235 1709 24281
rect 1621 24174 1709 24235
rect 1621 24128 1650 24174
rect 1696 24128 1709 24174
rect 1621 24067 1709 24128
rect 1621 24021 1650 24067
rect 1696 24021 1709 24067
rect 1621 24008 1709 24021
rect 2032 25357 2120 25370
rect 2032 25311 2045 25357
rect 2091 25311 2120 25357
rect 2032 25249 2120 25311
rect 2032 25203 2045 25249
rect 2091 25203 2120 25249
rect 2032 25141 2120 25203
rect 2032 25095 2045 25141
rect 2091 25095 2120 25141
rect 2032 25033 2120 25095
rect 2032 24987 2045 25033
rect 2091 24987 2120 25033
rect 2032 24925 2120 24987
rect 2032 24879 2045 24925
rect 2091 24879 2120 24925
rect 2032 24817 2120 24879
rect 2032 24771 2045 24817
rect 2091 24771 2120 24817
rect 2032 24709 2120 24771
rect 2032 24663 2045 24709
rect 2091 24663 2120 24709
rect 2032 24602 2120 24663
rect 2032 24556 2045 24602
rect 2091 24556 2120 24602
rect 2032 24495 2120 24556
rect 2032 24449 2045 24495
rect 2091 24449 2120 24495
rect 2032 24388 2120 24449
rect 2032 24342 2045 24388
rect 2091 24342 2120 24388
rect 2032 24281 2120 24342
rect 2032 24235 2045 24281
rect 2091 24235 2120 24281
rect 2032 24174 2120 24235
rect 2032 24128 2045 24174
rect 2091 24128 2120 24174
rect 2032 24067 2120 24128
rect 2032 24021 2045 24067
rect 2091 24021 2120 24067
rect 2032 24008 2120 24021
rect 2240 25357 2328 25370
rect 2240 25311 2269 25357
rect 2315 25311 2328 25357
rect 2240 25249 2328 25311
rect 2240 25203 2269 25249
rect 2315 25203 2328 25249
rect 2240 25141 2328 25203
rect 2240 25095 2269 25141
rect 2315 25095 2328 25141
rect 2240 25033 2328 25095
rect 2240 24987 2269 25033
rect 2315 24987 2328 25033
rect 2240 24925 2328 24987
rect 2240 24879 2269 24925
rect 2315 24879 2328 24925
rect 2240 24817 2328 24879
rect 2240 24771 2269 24817
rect 2315 24771 2328 24817
rect 2240 24709 2328 24771
rect 2240 24663 2269 24709
rect 2315 24663 2328 24709
rect 2652 25357 2740 25370
rect 2652 25311 2665 25357
rect 2711 25311 2740 25357
rect 2652 25249 2740 25311
rect 2652 25203 2665 25249
rect 2711 25203 2740 25249
rect 2652 25141 2740 25203
rect 2652 25095 2665 25141
rect 2711 25095 2740 25141
rect 2652 25033 2740 25095
rect 2652 24987 2665 25033
rect 2711 24987 2740 25033
rect 2652 24925 2740 24987
rect 2652 24879 2665 24925
rect 2711 24879 2740 24925
rect 2652 24817 2740 24879
rect 2652 24771 2665 24817
rect 2711 24771 2740 24817
rect 2652 24709 2740 24771
rect 2240 24602 2328 24663
rect 2240 24556 2269 24602
rect 2315 24556 2328 24602
rect 2240 24495 2328 24556
rect 2240 24449 2269 24495
rect 2315 24449 2328 24495
rect 2240 24388 2328 24449
rect 2652 24663 2665 24709
rect 2711 24663 2740 24709
rect 2652 24602 2740 24663
rect 2652 24556 2665 24602
rect 2711 24556 2740 24602
rect 2652 24495 2740 24556
rect 2652 24449 2665 24495
rect 2711 24449 2740 24495
rect 2240 24342 2269 24388
rect 2315 24342 2328 24388
rect 2240 24281 2328 24342
rect 2240 24235 2269 24281
rect 2315 24235 2328 24281
rect 2240 24174 2328 24235
rect 2240 24128 2269 24174
rect 2315 24128 2328 24174
rect 2240 24067 2328 24128
rect 2240 24021 2269 24067
rect 2315 24021 2328 24067
rect 2240 24008 2328 24021
rect 2652 24388 2740 24449
rect 2652 24342 2665 24388
rect 2711 24342 2740 24388
rect 2652 24281 2740 24342
rect 2652 24235 2665 24281
rect 2711 24235 2740 24281
rect 2652 24174 2740 24235
rect 2652 24128 2665 24174
rect 2711 24128 2740 24174
rect 2652 24067 2740 24128
rect 2652 24021 2665 24067
rect 2711 24021 2740 24067
rect 2652 24008 2740 24021
rect 2860 25357 2948 25370
rect 2860 25311 2889 25357
rect 2935 25311 2948 25357
rect 2860 25249 2948 25311
rect 2860 25203 2889 25249
rect 2935 25203 2948 25249
rect 2860 25141 2948 25203
rect 2860 25095 2889 25141
rect 2935 25095 2948 25141
rect 2860 25033 2948 25095
rect 2860 24987 2889 25033
rect 2935 24987 2948 25033
rect 2860 24925 2948 24987
rect 2860 24879 2889 24925
rect 2935 24879 2948 24925
rect 2860 24817 2948 24879
rect 2860 24771 2889 24817
rect 2935 24771 2948 24817
rect 2860 24709 2948 24771
rect 2860 24663 2889 24709
rect 2935 24663 2948 24709
rect 2860 24602 2948 24663
rect 2860 24556 2889 24602
rect 2935 24556 2948 24602
rect 2860 24495 2948 24556
rect 2860 24449 2889 24495
rect 2935 24449 2948 24495
rect 2860 24388 2948 24449
rect 2860 24342 2889 24388
rect 2935 24342 2948 24388
rect 2860 24281 2948 24342
rect 2860 24235 2889 24281
rect 2935 24235 2948 24281
rect 2860 24174 2948 24235
rect 2860 24128 2889 24174
rect 2935 24128 2948 24174
rect 2860 24067 2948 24128
rect 2860 24021 2889 24067
rect 2935 24021 2948 24067
rect 2860 24008 2948 24021
rect 3270 25357 3358 25370
rect 3270 25311 3283 25357
rect 3329 25311 3358 25357
rect 3270 25249 3358 25311
rect 3270 25203 3283 25249
rect 3329 25203 3358 25249
rect 3270 25141 3358 25203
rect 3270 25095 3283 25141
rect 3329 25095 3358 25141
rect 3270 25033 3358 25095
rect 3270 24987 3283 25033
rect 3329 24987 3358 25033
rect 3270 24925 3358 24987
rect 3270 24879 3283 24925
rect 3329 24879 3358 24925
rect 3270 24817 3358 24879
rect 3270 24771 3283 24817
rect 3329 24771 3358 24817
rect 3270 24709 3358 24771
rect 3270 24663 3283 24709
rect 3329 24663 3358 24709
rect 3270 24602 3358 24663
rect 3270 24556 3283 24602
rect 3329 24556 3358 24602
rect 3270 24495 3358 24556
rect 3270 24449 3283 24495
rect 3329 24449 3358 24495
rect 3270 24388 3358 24449
rect 3270 24342 3283 24388
rect 3329 24342 3358 24388
rect 3270 24281 3358 24342
rect 3270 24235 3283 24281
rect 3329 24235 3358 24281
rect 3270 24174 3358 24235
rect 3270 24128 3283 24174
rect 3329 24128 3358 24174
rect 3270 24067 3358 24128
rect 3270 24021 3283 24067
rect 3329 24021 3358 24067
rect 3270 24008 3358 24021
rect 3478 25357 3566 25370
rect 3478 25311 3507 25357
rect 3553 25311 3566 25357
rect 3478 25249 3566 25311
rect 3478 25203 3507 25249
rect 3553 25203 3566 25249
rect 3478 25141 3566 25203
rect 3478 25095 3507 25141
rect 3553 25095 3566 25141
rect 3478 25033 3566 25095
rect 3478 24987 3507 25033
rect 3553 24987 3566 25033
rect 3478 24925 3566 24987
rect 3478 24879 3507 24925
rect 3553 24879 3566 24925
rect 3478 24817 3566 24879
rect 3478 24771 3507 24817
rect 3553 24771 3566 24817
rect 3478 24709 3566 24771
rect 3478 24663 3507 24709
rect 3553 24663 3566 24709
rect 3890 25357 3978 25370
rect 3890 25311 3903 25357
rect 3949 25311 3978 25357
rect 3890 25249 3978 25311
rect 3890 25203 3903 25249
rect 3949 25203 3978 25249
rect 3890 25141 3978 25203
rect 3890 25095 3903 25141
rect 3949 25095 3978 25141
rect 3890 25033 3978 25095
rect 3890 24987 3903 25033
rect 3949 24987 3978 25033
rect 3890 24925 3978 24987
rect 3890 24879 3903 24925
rect 3949 24879 3978 24925
rect 3890 24817 3978 24879
rect 3890 24771 3903 24817
rect 3949 24771 3978 24817
rect 3890 24709 3978 24771
rect 3478 24602 3566 24663
rect 3478 24556 3507 24602
rect 3553 24556 3566 24602
rect 3478 24495 3566 24556
rect 3478 24449 3507 24495
rect 3553 24449 3566 24495
rect 3478 24388 3566 24449
rect 3890 24663 3903 24709
rect 3949 24663 3978 24709
rect 3890 24602 3978 24663
rect 3890 24556 3903 24602
rect 3949 24556 3978 24602
rect 3890 24495 3978 24556
rect 3890 24449 3903 24495
rect 3949 24449 3978 24495
rect 3478 24342 3507 24388
rect 3553 24342 3566 24388
rect 3478 24281 3566 24342
rect 3478 24235 3507 24281
rect 3553 24235 3566 24281
rect 3478 24174 3566 24235
rect 3478 24128 3507 24174
rect 3553 24128 3566 24174
rect 3478 24067 3566 24128
rect 3478 24021 3507 24067
rect 3553 24021 3566 24067
rect 3478 24008 3566 24021
rect 3890 24388 3978 24449
rect 3890 24342 3903 24388
rect 3949 24342 3978 24388
rect 3890 24281 3978 24342
rect 3890 24235 3903 24281
rect 3949 24235 3978 24281
rect 3890 24174 3978 24235
rect 3890 24128 3903 24174
rect 3949 24128 3978 24174
rect 3890 24067 3978 24128
rect 3890 24021 3903 24067
rect 3949 24021 3978 24067
rect 3890 24008 3978 24021
rect 4098 25357 4186 25370
rect 4098 25311 4127 25357
rect 4173 25311 4186 25357
rect 4098 25249 4186 25311
rect 4098 25203 4127 25249
rect 4173 25203 4186 25249
rect 4098 25141 4186 25203
rect 4098 25095 4127 25141
rect 4173 25095 4186 25141
rect 4098 25033 4186 25095
rect 4098 24987 4127 25033
rect 4173 24987 4186 25033
rect 4098 24925 4186 24987
rect 4098 24879 4127 24925
rect 4173 24879 4186 24925
rect 4098 24817 4186 24879
rect 4098 24771 4127 24817
rect 4173 24771 4186 24817
rect 4098 24709 4186 24771
rect 4098 24663 4127 24709
rect 4173 24663 4186 24709
rect 4098 24602 4186 24663
rect 4098 24556 4127 24602
rect 4173 24556 4186 24602
rect 4098 24495 4186 24556
rect 4098 24449 4127 24495
rect 4173 24449 4186 24495
rect 4098 24388 4186 24449
rect 4098 24342 4127 24388
rect 4173 24342 4186 24388
rect 4098 24281 4186 24342
rect 4098 24235 4127 24281
rect 4173 24235 4186 24281
rect 4098 24174 4186 24235
rect 4098 24128 4127 24174
rect 4173 24128 4186 24174
rect 4098 24067 4186 24128
rect 4098 24021 4127 24067
rect 4173 24021 4186 24067
rect 4098 24008 4186 24021
rect 4509 25357 4597 25370
rect 4509 25311 4522 25357
rect 4568 25311 4597 25357
rect 4509 25249 4597 25311
rect 4509 25203 4522 25249
rect 4568 25203 4597 25249
rect 4509 25141 4597 25203
rect 4509 25095 4522 25141
rect 4568 25095 4597 25141
rect 4509 25033 4597 25095
rect 4509 24987 4522 25033
rect 4568 24987 4597 25033
rect 4509 24925 4597 24987
rect 4509 24879 4522 24925
rect 4568 24879 4597 24925
rect 4509 24817 4597 24879
rect 4509 24771 4522 24817
rect 4568 24771 4597 24817
rect 4509 24709 4597 24771
rect 4509 24663 4522 24709
rect 4568 24663 4597 24709
rect 4509 24602 4597 24663
rect 4509 24556 4522 24602
rect 4568 24556 4597 24602
rect 4509 24495 4597 24556
rect 4509 24449 4522 24495
rect 4568 24449 4597 24495
rect 4509 24388 4597 24449
rect 4509 24342 4522 24388
rect 4568 24342 4597 24388
rect 4509 24281 4597 24342
rect 4509 24235 4522 24281
rect 4568 24235 4597 24281
rect 4509 24174 4597 24235
rect 4509 24128 4522 24174
rect 4568 24128 4597 24174
rect 4509 24067 4597 24128
rect 4509 24021 4522 24067
rect 4568 24021 4597 24067
rect 4509 24008 4597 24021
rect 4717 25357 4805 25370
rect 4717 25311 4746 25357
rect 4792 25311 4805 25357
rect 4717 25249 4805 25311
rect 4717 25203 4746 25249
rect 4792 25203 4805 25249
rect 4717 25141 4805 25203
rect 4717 25095 4746 25141
rect 4792 25095 4805 25141
rect 4717 25033 4805 25095
rect 4717 24987 4746 25033
rect 4792 24987 4805 25033
rect 4717 24925 4805 24987
rect 4717 24879 4746 24925
rect 4792 24879 4805 24925
rect 4717 24817 4805 24879
rect 4717 24771 4746 24817
rect 4792 24771 4805 24817
rect 4717 24709 4805 24771
rect 4717 24663 4746 24709
rect 4792 24663 4805 24709
rect 5129 25357 5217 25370
rect 5129 25311 5142 25357
rect 5188 25311 5217 25357
rect 5129 25249 5217 25311
rect 5129 25203 5142 25249
rect 5188 25203 5217 25249
rect 5129 25141 5217 25203
rect 5129 25095 5142 25141
rect 5188 25095 5217 25141
rect 5129 25033 5217 25095
rect 5129 24987 5142 25033
rect 5188 24987 5217 25033
rect 5129 24925 5217 24987
rect 5129 24879 5142 24925
rect 5188 24879 5217 24925
rect 5129 24817 5217 24879
rect 5129 24771 5142 24817
rect 5188 24771 5217 24817
rect 5129 24709 5217 24771
rect 4717 24602 4805 24663
rect 4717 24556 4746 24602
rect 4792 24556 4805 24602
rect 4717 24495 4805 24556
rect 4717 24449 4746 24495
rect 4792 24449 4805 24495
rect 4717 24388 4805 24449
rect 5129 24663 5142 24709
rect 5188 24663 5217 24709
rect 5129 24602 5217 24663
rect 5129 24556 5142 24602
rect 5188 24556 5217 24602
rect 5129 24495 5217 24556
rect 5129 24449 5142 24495
rect 5188 24449 5217 24495
rect 4717 24342 4746 24388
rect 4792 24342 4805 24388
rect 4717 24281 4805 24342
rect 4717 24235 4746 24281
rect 4792 24235 4805 24281
rect 4717 24174 4805 24235
rect 4717 24128 4746 24174
rect 4792 24128 4805 24174
rect 4717 24067 4805 24128
rect 4717 24021 4746 24067
rect 4792 24021 4805 24067
rect 4717 24008 4805 24021
rect 5129 24388 5217 24449
rect 5129 24342 5142 24388
rect 5188 24342 5217 24388
rect 5129 24281 5217 24342
rect 5129 24235 5142 24281
rect 5188 24235 5217 24281
rect 5129 24174 5217 24235
rect 5129 24128 5142 24174
rect 5188 24128 5217 24174
rect 5129 24067 5217 24128
rect 5129 24021 5142 24067
rect 5188 24021 5217 24067
rect 5129 24008 5217 24021
rect 5337 25357 5425 25370
rect 5337 25311 5366 25357
rect 5412 25311 5425 25357
rect 5337 25249 5425 25311
rect 5337 25203 5366 25249
rect 5412 25203 5425 25249
rect 5337 25141 5425 25203
rect 5337 25095 5366 25141
rect 5412 25095 5425 25141
rect 5337 25033 5425 25095
rect 5337 24987 5366 25033
rect 5412 24987 5425 25033
rect 5337 24925 5425 24987
rect 5337 24879 5366 24925
rect 5412 24879 5425 24925
rect 5337 24817 5425 24879
rect 5337 24771 5366 24817
rect 5412 24771 5425 24817
rect 5337 24709 5425 24771
rect 5337 24663 5366 24709
rect 5412 24663 5425 24709
rect 5337 24602 5425 24663
rect 5337 24556 5366 24602
rect 5412 24556 5425 24602
rect 5337 24495 5425 24556
rect 5337 24449 5366 24495
rect 5412 24449 5425 24495
rect 5337 24388 5425 24449
rect 5337 24342 5366 24388
rect 5412 24342 5425 24388
rect 5337 24281 5425 24342
rect 5337 24235 5366 24281
rect 5412 24235 5425 24281
rect 5337 24174 5425 24235
rect 5337 24128 5366 24174
rect 5412 24128 5425 24174
rect 5337 24067 5425 24128
rect 5337 24021 5366 24067
rect 5412 24021 5425 24067
rect 5337 24008 5425 24021
rect 793 19807 881 19820
rect 793 19761 806 19807
rect 852 19761 881 19807
rect 793 19699 881 19761
rect 793 19653 806 19699
rect 852 19653 881 19699
rect 793 19591 881 19653
rect 793 19545 806 19591
rect 852 19545 881 19591
rect 793 19483 881 19545
rect 793 19437 806 19483
rect 852 19437 881 19483
rect 793 19375 881 19437
rect 793 19329 806 19375
rect 852 19329 881 19375
rect 793 19267 881 19329
rect 793 19221 806 19267
rect 852 19221 881 19267
rect 793 19159 881 19221
rect 793 19113 806 19159
rect 852 19113 881 19159
rect 793 19052 881 19113
rect 793 19006 806 19052
rect 852 19006 881 19052
rect 793 18945 881 19006
rect 793 18899 806 18945
rect 852 18899 881 18945
rect 793 18838 881 18899
rect 793 18792 806 18838
rect 852 18792 881 18838
rect 793 18731 881 18792
rect 793 18685 806 18731
rect 852 18685 881 18731
rect 793 18624 881 18685
rect 793 18578 806 18624
rect 852 18578 881 18624
rect 793 18517 881 18578
rect 793 18471 806 18517
rect 852 18471 881 18517
rect 793 18458 881 18471
rect 1001 19807 1089 19820
rect 1001 19761 1030 19807
rect 1076 19761 1089 19807
rect 1001 19699 1089 19761
rect 1001 19653 1030 19699
rect 1076 19653 1089 19699
rect 1001 19591 1089 19653
rect 1001 19545 1030 19591
rect 1076 19545 1089 19591
rect 1001 19483 1089 19545
rect 1001 19437 1030 19483
rect 1076 19437 1089 19483
rect 1001 19375 1089 19437
rect 1001 19329 1030 19375
rect 1076 19329 1089 19375
rect 1001 19267 1089 19329
rect 1001 19221 1030 19267
rect 1076 19221 1089 19267
rect 1001 19159 1089 19221
rect 1001 19113 1030 19159
rect 1076 19113 1089 19159
rect 1001 19052 1089 19113
rect 1001 19006 1030 19052
rect 1076 19006 1089 19052
rect 1001 18945 1089 19006
rect 1001 18899 1030 18945
rect 1076 18899 1089 18945
rect 1001 18838 1089 18899
rect 1001 18792 1030 18838
rect 1076 18792 1089 18838
rect 1001 18731 1089 18792
rect 1001 18685 1030 18731
rect 1076 18685 1089 18731
rect 1001 18624 1089 18685
rect 1001 18578 1030 18624
rect 1076 18578 1089 18624
rect 1001 18517 1089 18578
rect 1001 18471 1030 18517
rect 1076 18471 1089 18517
rect 1001 18458 1089 18471
rect 1413 19807 1501 19820
rect 1413 19761 1426 19807
rect 1472 19761 1501 19807
rect 1413 19699 1501 19761
rect 1413 19653 1426 19699
rect 1472 19653 1501 19699
rect 1413 19591 1501 19653
rect 1413 19545 1426 19591
rect 1472 19545 1501 19591
rect 1413 19483 1501 19545
rect 1413 19437 1426 19483
rect 1472 19437 1501 19483
rect 1413 19375 1501 19437
rect 1413 19329 1426 19375
rect 1472 19329 1501 19375
rect 1413 19267 1501 19329
rect 1413 19221 1426 19267
rect 1472 19221 1501 19267
rect 1413 19159 1501 19221
rect 1413 19113 1426 19159
rect 1472 19113 1501 19159
rect 1413 19052 1501 19113
rect 1413 19006 1426 19052
rect 1472 19006 1501 19052
rect 1413 18945 1501 19006
rect 1413 18899 1426 18945
rect 1472 18899 1501 18945
rect 1413 18838 1501 18899
rect 1413 18792 1426 18838
rect 1472 18792 1501 18838
rect 1413 18731 1501 18792
rect 1413 18685 1426 18731
rect 1472 18685 1501 18731
rect 1413 18624 1501 18685
rect 1413 18578 1426 18624
rect 1472 18578 1501 18624
rect 1413 18517 1501 18578
rect 1413 18471 1426 18517
rect 1472 18471 1501 18517
rect 1413 18458 1501 18471
rect 1621 19807 1709 19820
rect 1621 19761 1650 19807
rect 1696 19761 1709 19807
rect 1621 19699 1709 19761
rect 1621 19653 1650 19699
rect 1696 19653 1709 19699
rect 1621 19591 1709 19653
rect 1621 19545 1650 19591
rect 1696 19545 1709 19591
rect 1621 19483 1709 19545
rect 1621 19437 1650 19483
rect 1696 19437 1709 19483
rect 1621 19375 1709 19437
rect 1621 19329 1650 19375
rect 1696 19329 1709 19375
rect 1621 19267 1709 19329
rect 1621 19221 1650 19267
rect 1696 19221 1709 19267
rect 1621 19159 1709 19221
rect 1621 19113 1650 19159
rect 1696 19113 1709 19159
rect 1621 19052 1709 19113
rect 1621 19006 1650 19052
rect 1696 19006 1709 19052
rect 1621 18945 1709 19006
rect 1621 18899 1650 18945
rect 1696 18899 1709 18945
rect 1621 18838 1709 18899
rect 1621 18792 1650 18838
rect 1696 18792 1709 18838
rect 1621 18731 1709 18792
rect 1621 18685 1650 18731
rect 1696 18685 1709 18731
rect 1621 18624 1709 18685
rect 1621 18578 1650 18624
rect 1696 18578 1709 18624
rect 1621 18517 1709 18578
rect 1621 18471 1650 18517
rect 1696 18471 1709 18517
rect 1621 18458 1709 18471
rect 2032 19807 2120 19820
rect 2032 19761 2045 19807
rect 2091 19761 2120 19807
rect 2032 19699 2120 19761
rect 2032 19653 2045 19699
rect 2091 19653 2120 19699
rect 2032 19591 2120 19653
rect 2032 19545 2045 19591
rect 2091 19545 2120 19591
rect 2032 19483 2120 19545
rect 2032 19437 2045 19483
rect 2091 19437 2120 19483
rect 2032 19375 2120 19437
rect 2032 19329 2045 19375
rect 2091 19329 2120 19375
rect 2032 19267 2120 19329
rect 2032 19221 2045 19267
rect 2091 19221 2120 19267
rect 2032 19159 2120 19221
rect 2032 19113 2045 19159
rect 2091 19113 2120 19159
rect 2032 19052 2120 19113
rect 2032 19006 2045 19052
rect 2091 19006 2120 19052
rect 2032 18945 2120 19006
rect 2032 18899 2045 18945
rect 2091 18899 2120 18945
rect 2032 18838 2120 18899
rect 2032 18792 2045 18838
rect 2091 18792 2120 18838
rect 2032 18731 2120 18792
rect 2032 18685 2045 18731
rect 2091 18685 2120 18731
rect 2032 18624 2120 18685
rect 2032 18578 2045 18624
rect 2091 18578 2120 18624
rect 2032 18517 2120 18578
rect 2032 18471 2045 18517
rect 2091 18471 2120 18517
rect 2032 18458 2120 18471
rect 2240 19807 2328 19820
rect 2240 19761 2269 19807
rect 2315 19761 2328 19807
rect 2240 19699 2328 19761
rect 2240 19653 2269 19699
rect 2315 19653 2328 19699
rect 2240 19591 2328 19653
rect 2240 19545 2269 19591
rect 2315 19545 2328 19591
rect 2240 19483 2328 19545
rect 2240 19437 2269 19483
rect 2315 19437 2328 19483
rect 2240 19375 2328 19437
rect 2240 19329 2269 19375
rect 2315 19329 2328 19375
rect 2240 19267 2328 19329
rect 2240 19221 2269 19267
rect 2315 19221 2328 19267
rect 2240 19159 2328 19221
rect 2240 19113 2269 19159
rect 2315 19113 2328 19159
rect 2240 19052 2328 19113
rect 2240 19006 2269 19052
rect 2315 19006 2328 19052
rect 2240 18945 2328 19006
rect 2240 18899 2269 18945
rect 2315 18899 2328 18945
rect 2240 18838 2328 18899
rect 2240 18792 2269 18838
rect 2315 18792 2328 18838
rect 2240 18731 2328 18792
rect 2240 18685 2269 18731
rect 2315 18685 2328 18731
rect 2240 18624 2328 18685
rect 2240 18578 2269 18624
rect 2315 18578 2328 18624
rect 2240 18517 2328 18578
rect 2240 18471 2269 18517
rect 2315 18471 2328 18517
rect 2240 18458 2328 18471
rect 2652 19807 2740 19820
rect 2652 19761 2665 19807
rect 2711 19761 2740 19807
rect 2652 19699 2740 19761
rect 2652 19653 2665 19699
rect 2711 19653 2740 19699
rect 2652 19591 2740 19653
rect 2652 19545 2665 19591
rect 2711 19545 2740 19591
rect 2652 19483 2740 19545
rect 2652 19437 2665 19483
rect 2711 19437 2740 19483
rect 2652 19375 2740 19437
rect 2652 19329 2665 19375
rect 2711 19329 2740 19375
rect 2652 19267 2740 19329
rect 2652 19221 2665 19267
rect 2711 19221 2740 19267
rect 2652 19159 2740 19221
rect 2652 19113 2665 19159
rect 2711 19113 2740 19159
rect 2652 19052 2740 19113
rect 2652 19006 2665 19052
rect 2711 19006 2740 19052
rect 2652 18945 2740 19006
rect 2652 18899 2665 18945
rect 2711 18899 2740 18945
rect 2652 18838 2740 18899
rect 2652 18792 2665 18838
rect 2711 18792 2740 18838
rect 2652 18731 2740 18792
rect 2652 18685 2665 18731
rect 2711 18685 2740 18731
rect 2652 18624 2740 18685
rect 2652 18578 2665 18624
rect 2711 18578 2740 18624
rect 2652 18517 2740 18578
rect 2652 18471 2665 18517
rect 2711 18471 2740 18517
rect 2652 18458 2740 18471
rect 2860 19807 2948 19820
rect 2860 19761 2889 19807
rect 2935 19761 2948 19807
rect 2860 19699 2948 19761
rect 2860 19653 2889 19699
rect 2935 19653 2948 19699
rect 2860 19591 2948 19653
rect 2860 19545 2889 19591
rect 2935 19545 2948 19591
rect 2860 19483 2948 19545
rect 2860 19437 2889 19483
rect 2935 19437 2948 19483
rect 2860 19375 2948 19437
rect 2860 19329 2889 19375
rect 2935 19329 2948 19375
rect 2860 19267 2948 19329
rect 2860 19221 2889 19267
rect 2935 19221 2948 19267
rect 2860 19159 2948 19221
rect 2860 19113 2889 19159
rect 2935 19113 2948 19159
rect 2860 19052 2948 19113
rect 2860 19006 2889 19052
rect 2935 19006 2948 19052
rect 2860 18945 2948 19006
rect 2860 18899 2889 18945
rect 2935 18899 2948 18945
rect 2860 18838 2948 18899
rect 2860 18792 2889 18838
rect 2935 18792 2948 18838
rect 2860 18731 2948 18792
rect 2860 18685 2889 18731
rect 2935 18685 2948 18731
rect 2860 18624 2948 18685
rect 2860 18578 2889 18624
rect 2935 18578 2948 18624
rect 2860 18517 2948 18578
rect 2860 18471 2889 18517
rect 2935 18471 2948 18517
rect 2860 18458 2948 18471
rect 3270 19807 3358 19820
rect 3270 19761 3283 19807
rect 3329 19761 3358 19807
rect 3270 19699 3358 19761
rect 3270 19653 3283 19699
rect 3329 19653 3358 19699
rect 3270 19591 3358 19653
rect 3270 19545 3283 19591
rect 3329 19545 3358 19591
rect 3270 19483 3358 19545
rect 3270 19437 3283 19483
rect 3329 19437 3358 19483
rect 3270 19375 3358 19437
rect 3270 19329 3283 19375
rect 3329 19329 3358 19375
rect 3270 19267 3358 19329
rect 3270 19221 3283 19267
rect 3329 19221 3358 19267
rect 3270 19159 3358 19221
rect 3270 19113 3283 19159
rect 3329 19113 3358 19159
rect 3270 19052 3358 19113
rect 3270 19006 3283 19052
rect 3329 19006 3358 19052
rect 3270 18945 3358 19006
rect 3270 18899 3283 18945
rect 3329 18899 3358 18945
rect 3270 18838 3358 18899
rect 3270 18792 3283 18838
rect 3329 18792 3358 18838
rect 3270 18731 3358 18792
rect 3270 18685 3283 18731
rect 3329 18685 3358 18731
rect 3270 18624 3358 18685
rect 3270 18578 3283 18624
rect 3329 18578 3358 18624
rect 3270 18517 3358 18578
rect 3270 18471 3283 18517
rect 3329 18471 3358 18517
rect 3270 18458 3358 18471
rect 3478 19807 3566 19820
rect 3478 19761 3507 19807
rect 3553 19761 3566 19807
rect 3478 19699 3566 19761
rect 3478 19653 3507 19699
rect 3553 19653 3566 19699
rect 3478 19591 3566 19653
rect 3478 19545 3507 19591
rect 3553 19545 3566 19591
rect 3478 19483 3566 19545
rect 3478 19437 3507 19483
rect 3553 19437 3566 19483
rect 3478 19375 3566 19437
rect 3478 19329 3507 19375
rect 3553 19329 3566 19375
rect 3478 19267 3566 19329
rect 3478 19221 3507 19267
rect 3553 19221 3566 19267
rect 3478 19159 3566 19221
rect 3478 19113 3507 19159
rect 3553 19113 3566 19159
rect 3478 19052 3566 19113
rect 3478 19006 3507 19052
rect 3553 19006 3566 19052
rect 3478 18945 3566 19006
rect 3478 18899 3507 18945
rect 3553 18899 3566 18945
rect 3478 18838 3566 18899
rect 3478 18792 3507 18838
rect 3553 18792 3566 18838
rect 3478 18731 3566 18792
rect 3478 18685 3507 18731
rect 3553 18685 3566 18731
rect 3478 18624 3566 18685
rect 3478 18578 3507 18624
rect 3553 18578 3566 18624
rect 3478 18517 3566 18578
rect 3478 18471 3507 18517
rect 3553 18471 3566 18517
rect 3478 18458 3566 18471
rect 3890 19807 3978 19820
rect 3890 19761 3903 19807
rect 3949 19761 3978 19807
rect 3890 19699 3978 19761
rect 3890 19653 3903 19699
rect 3949 19653 3978 19699
rect 3890 19591 3978 19653
rect 3890 19545 3903 19591
rect 3949 19545 3978 19591
rect 3890 19483 3978 19545
rect 3890 19437 3903 19483
rect 3949 19437 3978 19483
rect 3890 19375 3978 19437
rect 3890 19329 3903 19375
rect 3949 19329 3978 19375
rect 3890 19267 3978 19329
rect 3890 19221 3903 19267
rect 3949 19221 3978 19267
rect 3890 19159 3978 19221
rect 3890 19113 3903 19159
rect 3949 19113 3978 19159
rect 3890 19052 3978 19113
rect 3890 19006 3903 19052
rect 3949 19006 3978 19052
rect 3890 18945 3978 19006
rect 3890 18899 3903 18945
rect 3949 18899 3978 18945
rect 3890 18838 3978 18899
rect 3890 18792 3903 18838
rect 3949 18792 3978 18838
rect 3890 18731 3978 18792
rect 3890 18685 3903 18731
rect 3949 18685 3978 18731
rect 3890 18624 3978 18685
rect 3890 18578 3903 18624
rect 3949 18578 3978 18624
rect 3890 18517 3978 18578
rect 3890 18471 3903 18517
rect 3949 18471 3978 18517
rect 3890 18458 3978 18471
rect 4098 19807 4186 19820
rect 4098 19761 4127 19807
rect 4173 19761 4186 19807
rect 4098 19699 4186 19761
rect 4098 19653 4127 19699
rect 4173 19653 4186 19699
rect 4098 19591 4186 19653
rect 4098 19545 4127 19591
rect 4173 19545 4186 19591
rect 4098 19483 4186 19545
rect 4098 19437 4127 19483
rect 4173 19437 4186 19483
rect 4098 19375 4186 19437
rect 4098 19329 4127 19375
rect 4173 19329 4186 19375
rect 4098 19267 4186 19329
rect 4098 19221 4127 19267
rect 4173 19221 4186 19267
rect 4098 19159 4186 19221
rect 4098 19113 4127 19159
rect 4173 19113 4186 19159
rect 4098 19052 4186 19113
rect 4098 19006 4127 19052
rect 4173 19006 4186 19052
rect 4098 18945 4186 19006
rect 4098 18899 4127 18945
rect 4173 18899 4186 18945
rect 4098 18838 4186 18899
rect 4098 18792 4127 18838
rect 4173 18792 4186 18838
rect 4098 18731 4186 18792
rect 4098 18685 4127 18731
rect 4173 18685 4186 18731
rect 4098 18624 4186 18685
rect 4098 18578 4127 18624
rect 4173 18578 4186 18624
rect 4098 18517 4186 18578
rect 4098 18471 4127 18517
rect 4173 18471 4186 18517
rect 4098 18458 4186 18471
rect 4509 19807 4597 19820
rect 4509 19761 4522 19807
rect 4568 19761 4597 19807
rect 4509 19699 4597 19761
rect 4509 19653 4522 19699
rect 4568 19653 4597 19699
rect 4509 19591 4597 19653
rect 4509 19545 4522 19591
rect 4568 19545 4597 19591
rect 4509 19483 4597 19545
rect 4509 19437 4522 19483
rect 4568 19437 4597 19483
rect 4509 19375 4597 19437
rect 4509 19329 4522 19375
rect 4568 19329 4597 19375
rect 4509 19267 4597 19329
rect 4509 19221 4522 19267
rect 4568 19221 4597 19267
rect 4509 19159 4597 19221
rect 4509 19113 4522 19159
rect 4568 19113 4597 19159
rect 4509 19052 4597 19113
rect 4509 19006 4522 19052
rect 4568 19006 4597 19052
rect 4509 18945 4597 19006
rect 4509 18899 4522 18945
rect 4568 18899 4597 18945
rect 4509 18838 4597 18899
rect 4509 18792 4522 18838
rect 4568 18792 4597 18838
rect 4509 18731 4597 18792
rect 4509 18685 4522 18731
rect 4568 18685 4597 18731
rect 4509 18624 4597 18685
rect 4509 18578 4522 18624
rect 4568 18578 4597 18624
rect 4509 18517 4597 18578
rect 4509 18471 4522 18517
rect 4568 18471 4597 18517
rect 4509 18458 4597 18471
rect 4717 19807 4805 19820
rect 4717 19761 4746 19807
rect 4792 19761 4805 19807
rect 4717 19699 4805 19761
rect 4717 19653 4746 19699
rect 4792 19653 4805 19699
rect 4717 19591 4805 19653
rect 4717 19545 4746 19591
rect 4792 19545 4805 19591
rect 4717 19483 4805 19545
rect 4717 19437 4746 19483
rect 4792 19437 4805 19483
rect 4717 19375 4805 19437
rect 4717 19329 4746 19375
rect 4792 19329 4805 19375
rect 4717 19267 4805 19329
rect 4717 19221 4746 19267
rect 4792 19221 4805 19267
rect 4717 19159 4805 19221
rect 4717 19113 4746 19159
rect 4792 19113 4805 19159
rect 4717 19052 4805 19113
rect 4717 19006 4746 19052
rect 4792 19006 4805 19052
rect 4717 18945 4805 19006
rect 4717 18899 4746 18945
rect 4792 18899 4805 18945
rect 4717 18838 4805 18899
rect 4717 18792 4746 18838
rect 4792 18792 4805 18838
rect 4717 18731 4805 18792
rect 4717 18685 4746 18731
rect 4792 18685 4805 18731
rect 4717 18624 4805 18685
rect 4717 18578 4746 18624
rect 4792 18578 4805 18624
rect 4717 18517 4805 18578
rect 4717 18471 4746 18517
rect 4792 18471 4805 18517
rect 4717 18458 4805 18471
rect 5129 19807 5217 19820
rect 5129 19761 5142 19807
rect 5188 19761 5217 19807
rect 5129 19699 5217 19761
rect 5129 19653 5142 19699
rect 5188 19653 5217 19699
rect 5129 19591 5217 19653
rect 5129 19545 5142 19591
rect 5188 19545 5217 19591
rect 5129 19483 5217 19545
rect 5129 19437 5142 19483
rect 5188 19437 5217 19483
rect 5129 19375 5217 19437
rect 5129 19329 5142 19375
rect 5188 19329 5217 19375
rect 5129 19267 5217 19329
rect 5129 19221 5142 19267
rect 5188 19221 5217 19267
rect 5129 19159 5217 19221
rect 5129 19113 5142 19159
rect 5188 19113 5217 19159
rect 5129 19052 5217 19113
rect 5129 19006 5142 19052
rect 5188 19006 5217 19052
rect 5129 18945 5217 19006
rect 5129 18899 5142 18945
rect 5188 18899 5217 18945
rect 5129 18838 5217 18899
rect 5129 18792 5142 18838
rect 5188 18792 5217 18838
rect 5129 18731 5217 18792
rect 5129 18685 5142 18731
rect 5188 18685 5217 18731
rect 5129 18624 5217 18685
rect 5129 18578 5142 18624
rect 5188 18578 5217 18624
rect 5129 18517 5217 18578
rect 5129 18471 5142 18517
rect 5188 18471 5217 18517
rect 5129 18458 5217 18471
rect 5337 19807 5425 19820
rect 5337 19761 5366 19807
rect 5412 19761 5425 19807
rect 5337 19699 5425 19761
rect 5337 19653 5366 19699
rect 5412 19653 5425 19699
rect 5337 19591 5425 19653
rect 5337 19545 5366 19591
rect 5412 19545 5425 19591
rect 5337 19483 5425 19545
rect 5337 19437 5366 19483
rect 5412 19437 5425 19483
rect 5337 19375 5425 19437
rect 5337 19329 5366 19375
rect 5412 19329 5425 19375
rect 5337 19267 5425 19329
rect 5337 19221 5366 19267
rect 5412 19221 5425 19267
rect 5337 19159 5425 19221
rect 5337 19113 5366 19159
rect 5412 19113 5425 19159
rect 5337 19052 5425 19113
rect 5337 19006 5366 19052
rect 5412 19006 5425 19052
rect 5337 18945 5425 19006
rect 5337 18899 5366 18945
rect 5412 18899 5425 18945
rect 5337 18838 5425 18899
rect 5337 18792 5366 18838
rect 5412 18792 5425 18838
rect 5337 18731 5425 18792
rect 5337 18685 5366 18731
rect 5412 18685 5425 18731
rect 5337 18624 5425 18685
rect 5337 18578 5366 18624
rect 5412 18578 5425 18624
rect 5337 18517 5425 18578
rect 5337 18471 5366 18517
rect 5412 18471 5425 18517
rect 5337 18458 5425 18471
rect 631 17720 812 17845
rect 631 17674 725 17720
rect 771 17674 812 17720
rect 631 17548 812 17674
rect 932 17720 1064 17845
rect 932 17674 975 17720
rect 1021 17674 1064 17720
rect 932 17548 1064 17674
rect 1184 17720 1318 17845
rect 1184 17674 1228 17720
rect 1274 17674 1318 17720
rect 1184 17548 1318 17674
rect 1438 17720 1570 17845
rect 1438 17674 1481 17720
rect 1527 17674 1570 17720
rect 1438 17548 1570 17674
rect 1690 17720 2051 17845
rect 1690 17674 1731 17720
rect 1777 17674 1964 17720
rect 2010 17674 2051 17720
rect 1690 17548 2051 17674
rect 2171 17720 2303 17845
rect 2171 17674 2214 17720
rect 2260 17674 2303 17720
rect 2171 17548 2303 17674
rect 2423 17720 2557 17845
rect 2423 17674 2467 17720
rect 2513 17674 2557 17720
rect 2423 17548 2557 17674
rect 2677 17720 2809 17845
rect 2677 17674 2720 17720
rect 2766 17674 2809 17720
rect 2677 17548 2809 17674
rect 2929 17720 3289 17845
rect 2929 17674 2970 17720
rect 3016 17674 3202 17720
rect 3248 17674 3289 17720
rect 2929 17548 3289 17674
rect 3409 17720 3541 17845
rect 3409 17674 3452 17720
rect 3498 17674 3541 17720
rect 3409 17548 3541 17674
rect 3661 17720 3795 17845
rect 3661 17674 3705 17720
rect 3751 17674 3795 17720
rect 3661 17548 3795 17674
rect 3915 17720 4047 17845
rect 3915 17674 3958 17720
rect 4004 17674 4047 17720
rect 3915 17548 4047 17674
rect 4167 17720 4528 17845
rect 4167 17674 4208 17720
rect 4254 17674 4441 17720
rect 4487 17674 4528 17720
rect 4167 17548 4528 17674
rect 4648 17720 4780 17845
rect 4648 17674 4691 17720
rect 4737 17674 4780 17720
rect 4648 17548 4780 17674
rect 4900 17720 5034 17845
rect 4900 17674 4944 17720
rect 4990 17674 5034 17720
rect 4900 17548 5034 17674
rect 5154 17720 5285 17845
rect 5154 17674 5197 17720
rect 5243 17674 5285 17720
rect 5154 17548 5285 17674
rect 5405 17720 5587 17845
rect 5405 17674 5447 17720
rect 5493 17674 5587 17720
rect 5405 17548 5587 17674
rect 287 15765 375 15778
rect 287 13069 300 15765
rect 346 13069 375 15765
rect 287 13056 375 13069
rect 495 15765 583 15778
rect 495 13069 524 15765
rect 570 13069 583 15765
rect 1631 15311 1719 15324
rect 1631 15265 1644 15311
rect 1690 15265 1719 15311
rect 1631 15207 1719 15265
rect 810 15072 928 15197
rect 810 15026 853 15072
rect 899 15026 928 15072
rect 810 14900 928 15026
rect 1048 15072 1201 15197
rect 1048 15026 1117 15072
rect 1163 15026 1201 15072
rect 1048 14900 1201 15026
rect 1321 15072 1439 15197
rect 1321 15026 1350 15072
rect 1396 15026 1439 15072
rect 1321 14900 1439 15026
rect 1631 15161 1644 15207
rect 1690 15161 1719 15207
rect 1631 15103 1719 15161
rect 1631 15057 1644 15103
rect 1690 15057 1719 15103
rect 1631 14999 1719 15057
rect 1631 14953 1644 14999
rect 1690 14953 1719 14999
rect 1631 14895 1719 14953
rect 1631 14849 1644 14895
rect 1690 14849 1719 14895
rect 1631 14791 1719 14849
rect 1631 14745 1644 14791
rect 1690 14745 1719 14791
rect 1631 14687 1719 14745
rect 1631 14641 1644 14687
rect 1690 14641 1719 14687
rect 1631 14583 1719 14641
rect 1631 14537 1644 14583
rect 1690 14537 1719 14583
rect 1631 14479 1719 14537
rect 1631 14433 1644 14479
rect 1690 14433 1719 14479
rect 495 13056 583 13069
rect 735 14405 823 14418
rect 735 14359 748 14405
rect 794 14359 823 14405
rect 735 14298 823 14359
rect 735 14252 748 14298
rect 794 14252 823 14298
rect 735 14191 823 14252
rect 735 14145 748 14191
rect 794 14145 823 14191
rect 735 14084 823 14145
rect 735 14038 748 14084
rect 794 14038 823 14084
rect 735 13977 823 14038
rect 735 13931 748 13977
rect 794 13931 823 13977
rect 735 13870 823 13931
rect 735 13824 748 13870
rect 794 13824 823 13870
rect 735 13763 823 13824
rect 735 13717 748 13763
rect 794 13717 823 13763
rect 735 13655 823 13717
rect 735 13609 748 13655
rect 794 13609 823 13655
rect 735 13547 823 13609
rect 735 13501 748 13547
rect 794 13501 823 13547
rect 735 13439 823 13501
rect 735 13393 748 13439
rect 794 13393 823 13439
rect 735 13331 823 13393
rect 735 13285 748 13331
rect 794 13285 823 13331
rect 735 13223 823 13285
rect 735 13177 748 13223
rect 794 13177 823 13223
rect 735 13115 823 13177
rect 735 13069 748 13115
rect 794 13069 823 13115
rect 735 13056 823 13069
rect 943 14405 1031 14418
rect 943 14359 972 14405
rect 1018 14359 1031 14405
rect 943 14298 1031 14359
rect 943 14252 972 14298
rect 1018 14252 1031 14298
rect 943 14191 1031 14252
rect 943 14145 972 14191
rect 1018 14145 1031 14191
rect 943 14084 1031 14145
rect 943 14038 972 14084
rect 1018 14038 1031 14084
rect 943 13977 1031 14038
rect 943 13931 972 13977
rect 1018 13931 1031 13977
rect 943 13870 1031 13931
rect 943 13824 972 13870
rect 1018 13824 1031 13870
rect 943 13763 1031 13824
rect 943 13717 972 13763
rect 1018 13717 1031 13763
rect 943 13655 1031 13717
rect 943 13609 972 13655
rect 1018 13609 1031 13655
rect 943 13547 1031 13609
rect 943 13501 972 13547
rect 1018 13501 1031 13547
rect 943 13439 1031 13501
rect 943 13393 972 13439
rect 1018 13393 1031 13439
rect 943 13331 1031 13393
rect 943 13285 972 13331
rect 1018 13285 1031 13331
rect 943 13223 1031 13285
rect 943 13177 972 13223
rect 1018 13177 1031 13223
rect 943 13115 1031 13177
rect 943 13069 972 13115
rect 1018 13069 1031 13115
rect 943 13056 1031 13069
rect 1183 14405 1271 14418
rect 1183 14359 1196 14405
rect 1242 14359 1271 14405
rect 1183 14298 1271 14359
rect 1183 14252 1196 14298
rect 1242 14252 1271 14298
rect 1183 14191 1271 14252
rect 1183 14145 1196 14191
rect 1242 14145 1271 14191
rect 1183 14084 1271 14145
rect 1183 14038 1196 14084
rect 1242 14038 1271 14084
rect 1183 13977 1271 14038
rect 1183 13931 1196 13977
rect 1242 13931 1271 13977
rect 1183 13870 1271 13931
rect 1183 13824 1196 13870
rect 1242 13824 1271 13870
rect 1183 13763 1271 13824
rect 1183 13717 1196 13763
rect 1242 13717 1271 13763
rect 1183 13655 1271 13717
rect 1183 13609 1196 13655
rect 1242 13609 1271 13655
rect 1183 13547 1271 13609
rect 1183 13501 1196 13547
rect 1242 13501 1271 13547
rect 1183 13439 1271 13501
rect 1183 13393 1196 13439
rect 1242 13393 1271 13439
rect 1183 13331 1271 13393
rect 1183 13285 1196 13331
rect 1242 13285 1271 13331
rect 1183 13223 1271 13285
rect 1183 13177 1196 13223
rect 1242 13177 1271 13223
rect 1183 13115 1271 13177
rect 1183 13069 1196 13115
rect 1242 13069 1271 13115
rect 1183 13056 1271 13069
rect 1391 14405 1479 14418
rect 1391 14359 1420 14405
rect 1466 14359 1479 14405
rect 1391 14298 1479 14359
rect 1391 14252 1420 14298
rect 1466 14252 1479 14298
rect 1391 14191 1479 14252
rect 1391 14145 1420 14191
rect 1466 14145 1479 14191
rect 1391 14084 1479 14145
rect 1391 14038 1420 14084
rect 1466 14038 1479 14084
rect 1391 13977 1479 14038
rect 1391 13931 1420 13977
rect 1466 13931 1479 13977
rect 1391 13870 1479 13931
rect 1391 13824 1420 13870
rect 1466 13824 1479 13870
rect 1391 13763 1479 13824
rect 1391 13717 1420 13763
rect 1466 13717 1479 13763
rect 1391 13655 1479 13717
rect 1391 13609 1420 13655
rect 1466 13609 1479 13655
rect 1391 13547 1479 13609
rect 1391 13501 1420 13547
rect 1466 13501 1479 13547
rect 1391 13439 1479 13501
rect 1391 13393 1420 13439
rect 1466 13393 1479 13439
rect 1391 13331 1479 13393
rect 1391 13285 1420 13331
rect 1466 13285 1479 13331
rect 1391 13223 1479 13285
rect 1391 13177 1420 13223
rect 1466 13177 1479 13223
rect 1391 13115 1479 13177
rect 1391 13069 1420 13115
rect 1466 13069 1479 13115
rect 1391 13056 1479 13069
rect 1631 14375 1719 14433
rect 1631 14329 1644 14375
rect 1690 14329 1719 14375
rect 1631 14270 1719 14329
rect 1631 14224 1644 14270
rect 1690 14224 1719 14270
rect 1631 14165 1719 14224
rect 1631 14119 1644 14165
rect 1690 14119 1719 14165
rect 1631 14060 1719 14119
rect 1631 14014 1644 14060
rect 1690 14014 1719 14060
rect 1631 13955 1719 14014
rect 1631 13909 1644 13955
rect 1690 13909 1719 13955
rect 1631 13850 1719 13909
rect 1631 13804 1644 13850
rect 1690 13804 1719 13850
rect 1631 13745 1719 13804
rect 1631 13699 1644 13745
rect 1690 13699 1719 13745
rect 1631 13640 1719 13699
rect 1631 13594 1644 13640
rect 1690 13594 1719 13640
rect 1631 13535 1719 13594
rect 1631 13489 1644 13535
rect 1690 13489 1719 13535
rect 1631 13430 1719 13489
rect 1631 13384 1644 13430
rect 1690 13384 1719 13430
rect 1631 13325 1719 13384
rect 1631 13279 1644 13325
rect 1690 13279 1719 13325
rect 1631 13220 1719 13279
rect 1631 13174 1644 13220
rect 1690 13174 1719 13220
rect 1631 13115 1719 13174
rect 1631 13069 1644 13115
rect 1690 13069 1719 13115
rect 1631 13056 1719 13069
rect 1839 15311 1927 15324
rect 1839 15265 1868 15311
rect 1914 15265 1927 15311
rect 1839 15207 1927 15265
rect 1839 15161 1868 15207
rect 1914 15161 1927 15207
rect 1839 15103 1927 15161
rect 1839 15057 1868 15103
rect 1914 15057 1927 15103
rect 1839 14999 1927 15057
rect 1839 14953 1868 14999
rect 1914 14953 1927 14999
rect 1839 14895 1927 14953
rect 1839 14849 1868 14895
rect 1914 14849 1927 14895
rect 1839 14791 1927 14849
rect 1839 14745 1868 14791
rect 1914 14745 1927 14791
rect 1839 14687 1927 14745
rect 1839 14641 1868 14687
rect 1914 14641 1927 14687
rect 1839 14583 1927 14641
rect 1839 14537 1868 14583
rect 1914 14537 1927 14583
rect 1839 14479 1927 14537
rect 1839 14433 1868 14479
rect 1914 14433 1927 14479
rect 1839 14375 1927 14433
rect 1839 14329 1868 14375
rect 1914 14329 1927 14375
rect 1839 14270 1927 14329
rect 1839 14224 1868 14270
rect 1914 14224 1927 14270
rect 1839 14165 1927 14224
rect 1839 14119 1868 14165
rect 1914 14119 1927 14165
rect 1839 14060 1927 14119
rect 1839 14014 1868 14060
rect 1914 14014 1927 14060
rect 1839 13955 1927 14014
rect 1839 13909 1868 13955
rect 1914 13909 1927 13955
rect 1839 13850 1927 13909
rect 1839 13804 1868 13850
rect 1914 13804 1927 13850
rect 1839 13745 1927 13804
rect 1839 13699 1868 13745
rect 1914 13699 1927 13745
rect 1839 13640 1927 13699
rect 1839 13594 1868 13640
rect 1914 13594 1927 13640
rect 1839 13535 1927 13594
rect 1839 13489 1868 13535
rect 1914 13489 1927 13535
rect 1839 13430 1927 13489
rect 1839 13384 1868 13430
rect 1914 13384 1927 13430
rect 1839 13325 1927 13384
rect 1839 13279 1868 13325
rect 1914 13279 1927 13325
rect 1839 13220 1927 13279
rect 1839 13174 1868 13220
rect 1914 13174 1927 13220
rect 1839 13115 1927 13174
rect 1839 13069 1868 13115
rect 1914 13069 1927 13115
rect 1839 13056 1927 13069
rect 1616 9427 1704 9440
rect 1616 9381 1629 9427
rect 1675 9381 1704 9427
rect 1616 9271 1704 9381
rect 788 9234 876 9247
rect 788 9188 801 9234
rect 847 9188 876 9234
rect 788 9078 876 9188
rect 788 9032 801 9078
rect 847 9032 876 9078
rect 788 9019 876 9032
rect 996 9234 1100 9247
rect 996 9188 1025 9234
rect 1071 9188 1100 9234
rect 996 9078 1100 9188
rect 996 9032 1025 9078
rect 1071 9032 1100 9078
rect 996 9019 1100 9032
rect 1220 9234 1308 9247
rect 1220 9188 1249 9234
rect 1295 9188 1308 9234
rect 1616 9225 1629 9271
rect 1675 9225 1704 9271
rect 1616 9212 1704 9225
rect 1824 9427 1928 9440
rect 1824 9381 1853 9427
rect 1899 9381 1928 9427
rect 1824 9271 1928 9381
rect 1824 9225 1853 9271
rect 1899 9225 1928 9271
rect 1824 9212 1928 9225
rect 2048 9427 2136 9440
rect 2048 9381 2077 9427
rect 2123 9381 2136 9427
rect 2048 9271 2136 9381
rect 2048 9225 2077 9271
rect 2123 9225 2136 9271
rect 2048 9212 2136 9225
rect 2468 9252 2556 9265
rect 1220 9078 1308 9188
rect 2468 9206 2481 9252
rect 2527 9206 2556 9252
rect 2468 9145 2556 9206
rect 1220 9032 1249 9078
rect 1295 9032 1308 9078
rect 2468 9099 2481 9145
rect 2527 9099 2556 9145
rect 1220 9019 1308 9032
rect 2468 9038 2556 9099
rect 2468 8992 2481 9038
rect 2527 8992 2556 9038
rect 2468 8931 2556 8992
rect 2468 8885 2481 8931
rect 2527 8885 2556 8931
rect 2468 8824 2556 8885
rect 2468 8778 2481 8824
rect 2527 8778 2556 8824
rect 1616 8712 1704 8725
rect 1616 8666 1629 8712
rect 1675 8666 1704 8712
rect 788 8630 876 8643
rect 788 8584 801 8630
rect 847 8584 876 8630
rect 788 8510 876 8584
rect 788 8464 801 8510
rect 847 8464 876 8510
rect 788 8451 876 8464
rect 996 8630 1100 8643
rect 996 8584 1025 8630
rect 1071 8584 1100 8630
rect 996 8510 1100 8584
rect 996 8464 1025 8510
rect 1071 8464 1100 8510
rect 996 8451 1100 8464
rect 1220 8630 1308 8643
rect 1220 8584 1249 8630
rect 1295 8584 1308 8630
rect 1220 8510 1308 8584
rect 1616 8592 1704 8666
rect 1616 8546 1629 8592
rect 1675 8546 1704 8592
rect 1616 8533 1704 8546
rect 1824 8712 1928 8725
rect 1824 8666 1853 8712
rect 1899 8666 1928 8712
rect 1824 8592 1928 8666
rect 1824 8546 1853 8592
rect 1899 8546 1928 8592
rect 1824 8533 1928 8546
rect 2048 8712 2136 8725
rect 2048 8666 2077 8712
rect 2123 8666 2136 8712
rect 2048 8592 2136 8666
rect 2048 8546 2077 8592
rect 2123 8546 2136 8592
rect 2048 8533 2136 8546
rect 2468 8717 2556 8778
rect 2468 8671 2481 8717
rect 2527 8671 2556 8717
rect 2468 8610 2556 8671
rect 2468 8564 2481 8610
rect 2527 8564 2556 8610
rect 1220 8464 1249 8510
rect 1295 8464 1308 8510
rect 1220 8451 1308 8464
rect 2468 8502 2556 8564
rect 2468 8456 2481 8502
rect 2527 8456 2556 8502
rect 2468 8394 2556 8456
rect 2468 8348 2481 8394
rect 2527 8348 2556 8394
rect 2468 8286 2556 8348
rect 2468 8240 2481 8286
rect 2527 8240 2556 8286
rect 2468 8178 2556 8240
rect 2468 8132 2481 8178
rect 2527 8132 2556 8178
rect 2468 8070 2556 8132
rect 2468 8024 2481 8070
rect 2527 8024 2556 8070
rect 2468 7962 2556 8024
rect 2468 7916 2481 7962
rect 2527 7916 2556 7962
rect 2468 7903 2556 7916
rect 2676 9252 2764 9265
rect 2676 9206 2705 9252
rect 2751 9206 2764 9252
rect 2676 9145 2764 9206
rect 2676 9099 2705 9145
rect 2751 9099 2764 9145
rect 2676 9038 2764 9099
rect 2676 8992 2705 9038
rect 2751 8992 2764 9038
rect 2676 8931 2764 8992
rect 2676 8885 2705 8931
rect 2751 8885 2764 8931
rect 2676 8824 2764 8885
rect 2676 8778 2705 8824
rect 2751 8778 2764 8824
rect 2676 8717 2764 8778
rect 2676 8671 2705 8717
rect 2751 8671 2764 8717
rect 2676 8610 2764 8671
rect 2676 8564 2705 8610
rect 2751 8564 2764 8610
rect 2676 8502 2764 8564
rect 2676 8456 2705 8502
rect 2751 8456 2764 8502
rect 2676 8394 2764 8456
rect 2676 8348 2705 8394
rect 2751 8348 2764 8394
rect 2676 8286 2764 8348
rect 2676 8240 2705 8286
rect 2751 8240 2764 8286
rect 2676 8178 2764 8240
rect 2676 8132 2705 8178
rect 2751 8132 2764 8178
rect 2676 8070 2764 8132
rect 2676 8024 2705 8070
rect 2751 8024 2764 8070
rect 2676 7962 2764 8024
rect 2676 7916 2705 7962
rect 2751 7916 2764 7962
rect 2676 7903 2764 7916
<< mvndiffc >>
rect 806 23620 852 23666
rect 806 23512 852 23558
rect 806 23404 852 23450
rect 806 23296 852 23342
rect 806 23188 852 23234
rect 806 23080 852 23126
rect 806 22972 852 23018
rect 806 22865 852 22911
rect 806 22758 852 22804
rect 806 22651 852 22697
rect 806 22544 852 22590
rect 806 22437 852 22483
rect 806 22330 852 22376
rect 1030 23620 1076 23666
rect 1030 23512 1076 23558
rect 1030 23404 1076 23450
rect 1030 23296 1076 23342
rect 1030 23188 1076 23234
rect 1030 23080 1076 23126
rect 1030 22972 1076 23018
rect 1030 22865 1076 22911
rect 1030 22758 1076 22804
rect 1030 22651 1076 22697
rect 1030 22544 1076 22590
rect 1030 22437 1076 22483
rect 1030 22330 1076 22376
rect 1426 23620 1472 23666
rect 1426 23512 1472 23558
rect 1426 23404 1472 23450
rect 1426 23296 1472 23342
rect 1426 23188 1472 23234
rect 1426 23080 1472 23126
rect 1426 22972 1472 23018
rect 1426 22865 1472 22911
rect 1426 22758 1472 22804
rect 1426 22651 1472 22697
rect 1426 22544 1472 22590
rect 1426 22437 1472 22483
rect 1426 22330 1472 22376
rect 1650 23620 1696 23666
rect 1650 23512 1696 23558
rect 1650 23404 1696 23450
rect 1650 23296 1696 23342
rect 1650 23188 1696 23234
rect 1650 23080 1696 23126
rect 1650 22972 1696 23018
rect 1650 22865 1696 22911
rect 1650 22758 1696 22804
rect 1650 22651 1696 22697
rect 1650 22544 1696 22590
rect 1650 22437 1696 22483
rect 1650 22330 1696 22376
rect 2045 23620 2091 23666
rect 2045 23512 2091 23558
rect 2045 23404 2091 23450
rect 2045 23296 2091 23342
rect 2045 23188 2091 23234
rect 2045 23080 2091 23126
rect 2045 22972 2091 23018
rect 2045 22865 2091 22911
rect 2045 22758 2091 22804
rect 2045 22651 2091 22697
rect 2045 22544 2091 22590
rect 2045 22437 2091 22483
rect 2045 22330 2091 22376
rect 2269 23620 2315 23666
rect 2269 23512 2315 23558
rect 2269 23404 2315 23450
rect 2269 23296 2315 23342
rect 2269 23188 2315 23234
rect 2269 23080 2315 23126
rect 2269 22972 2315 23018
rect 2269 22865 2315 22911
rect 2269 22758 2315 22804
rect 2269 22651 2315 22697
rect 2269 22544 2315 22590
rect 2269 22437 2315 22483
rect 2269 22330 2315 22376
rect 2665 23620 2711 23666
rect 2665 23512 2711 23558
rect 2665 23404 2711 23450
rect 2665 23296 2711 23342
rect 2665 23188 2711 23234
rect 2665 23080 2711 23126
rect 2665 22972 2711 23018
rect 2665 22865 2711 22911
rect 2665 22758 2711 22804
rect 2665 22651 2711 22697
rect 2665 22544 2711 22590
rect 2665 22437 2711 22483
rect 2665 22330 2711 22376
rect 2889 23620 2935 23666
rect 2889 23512 2935 23558
rect 2889 23404 2935 23450
rect 2889 23296 2935 23342
rect 2889 23188 2935 23234
rect 2889 23080 2935 23126
rect 2889 22972 2935 23018
rect 2889 22865 2935 22911
rect 2889 22758 2935 22804
rect 2889 22651 2935 22697
rect 2889 22544 2935 22590
rect 2889 22437 2935 22483
rect 2889 22330 2935 22376
rect 3283 23620 3329 23666
rect 3283 23512 3329 23558
rect 3283 23404 3329 23450
rect 3283 23296 3329 23342
rect 3283 23188 3329 23234
rect 3283 23080 3329 23126
rect 3283 22972 3329 23018
rect 3283 22865 3329 22911
rect 3283 22758 3329 22804
rect 3283 22651 3329 22697
rect 3283 22544 3329 22590
rect 3283 22437 3329 22483
rect 3283 22330 3329 22376
rect 3507 23620 3553 23666
rect 3507 23512 3553 23558
rect 3507 23404 3553 23450
rect 3507 23296 3553 23342
rect 3507 23188 3553 23234
rect 3507 23080 3553 23126
rect 3507 22972 3553 23018
rect 3507 22865 3553 22911
rect 3507 22758 3553 22804
rect 3507 22651 3553 22697
rect 3507 22544 3553 22590
rect 3507 22437 3553 22483
rect 3507 22330 3553 22376
rect 3903 23620 3949 23666
rect 3903 23512 3949 23558
rect 3903 23404 3949 23450
rect 3903 23296 3949 23342
rect 3903 23188 3949 23234
rect 3903 23080 3949 23126
rect 3903 22972 3949 23018
rect 3903 22865 3949 22911
rect 3903 22758 3949 22804
rect 3903 22651 3949 22697
rect 3903 22544 3949 22590
rect 3903 22437 3949 22483
rect 3903 22330 3949 22376
rect 4127 23620 4173 23666
rect 4127 23512 4173 23558
rect 4127 23404 4173 23450
rect 4127 23296 4173 23342
rect 4127 23188 4173 23234
rect 4127 23080 4173 23126
rect 4127 22972 4173 23018
rect 4127 22865 4173 22911
rect 4127 22758 4173 22804
rect 4127 22651 4173 22697
rect 4127 22544 4173 22590
rect 4127 22437 4173 22483
rect 4127 22330 4173 22376
rect 4522 23620 4568 23666
rect 4522 23512 4568 23558
rect 4522 23404 4568 23450
rect 4522 23296 4568 23342
rect 4522 23188 4568 23234
rect 4522 23080 4568 23126
rect 4522 22972 4568 23018
rect 4522 22865 4568 22911
rect 4522 22758 4568 22804
rect 4522 22651 4568 22697
rect 4522 22544 4568 22590
rect 4522 22437 4568 22483
rect 4522 22330 4568 22376
rect 4746 23620 4792 23666
rect 4746 23512 4792 23558
rect 4746 23404 4792 23450
rect 4746 23296 4792 23342
rect 4746 23188 4792 23234
rect 4746 23080 4792 23126
rect 4746 22972 4792 23018
rect 4746 22865 4792 22911
rect 4746 22758 4792 22804
rect 4746 22651 4792 22697
rect 4746 22544 4792 22590
rect 4746 22437 4792 22483
rect 4746 22330 4792 22376
rect 5142 23620 5188 23666
rect 5142 23512 5188 23558
rect 5142 23404 5188 23450
rect 5142 23296 5188 23342
rect 5142 23188 5188 23234
rect 5142 23080 5188 23126
rect 5142 22972 5188 23018
rect 5142 22865 5188 22911
rect 5142 22758 5188 22804
rect 5142 22651 5188 22697
rect 5142 22544 5188 22590
rect 5142 22437 5188 22483
rect 5142 22330 5188 22376
rect 5366 23620 5412 23666
rect 5366 23512 5412 23558
rect 5366 23404 5412 23450
rect 5366 23296 5412 23342
rect 5366 23188 5412 23234
rect 5366 23080 5412 23126
rect 5366 22972 5412 23018
rect 5366 22865 5412 22911
rect 5366 22758 5412 22804
rect 5366 22651 5412 22697
rect 5366 22544 5412 22590
rect 5366 22437 5412 22483
rect 5366 22330 5412 22376
rect 806 21616 852 21662
rect 806 21508 852 21554
rect 806 21400 852 21446
rect 806 21292 852 21338
rect 806 21184 852 21230
rect 806 21076 852 21122
rect 806 20968 852 21014
rect 806 20861 852 20907
rect 806 20754 852 20800
rect 806 20647 852 20693
rect 806 20540 852 20586
rect 806 20433 852 20479
rect 806 20326 852 20372
rect 1030 21616 1076 21662
rect 1030 21508 1076 21554
rect 1030 21400 1076 21446
rect 1030 21292 1076 21338
rect 1030 21184 1076 21230
rect 1030 21076 1076 21122
rect 1030 20968 1076 21014
rect 1030 20861 1076 20907
rect 1030 20754 1076 20800
rect 1030 20647 1076 20693
rect 1030 20540 1076 20586
rect 1030 20433 1076 20479
rect 1030 20326 1076 20372
rect 1426 21616 1472 21662
rect 1426 21508 1472 21554
rect 1426 21400 1472 21446
rect 1426 21292 1472 21338
rect 1426 21184 1472 21230
rect 1426 21076 1472 21122
rect 1426 20968 1472 21014
rect 1426 20861 1472 20907
rect 1426 20754 1472 20800
rect 1426 20647 1472 20693
rect 1426 20540 1472 20586
rect 1426 20433 1472 20479
rect 1426 20326 1472 20372
rect 1650 21616 1696 21662
rect 1650 21508 1696 21554
rect 1650 21400 1696 21446
rect 1650 21292 1696 21338
rect 1650 21184 1696 21230
rect 1650 21076 1696 21122
rect 1650 20968 1696 21014
rect 1650 20861 1696 20907
rect 1650 20754 1696 20800
rect 1650 20647 1696 20693
rect 1650 20540 1696 20586
rect 1650 20433 1696 20479
rect 1650 20326 1696 20372
rect 2045 21616 2091 21662
rect 2045 21508 2091 21554
rect 2045 21400 2091 21446
rect 2045 21292 2091 21338
rect 2045 21184 2091 21230
rect 2045 21076 2091 21122
rect 2045 20968 2091 21014
rect 2045 20861 2091 20907
rect 2045 20754 2091 20800
rect 2045 20647 2091 20693
rect 2045 20540 2091 20586
rect 2045 20433 2091 20479
rect 2045 20326 2091 20372
rect 2269 21616 2315 21662
rect 2269 21508 2315 21554
rect 2269 21400 2315 21446
rect 2269 21292 2315 21338
rect 2269 21184 2315 21230
rect 2269 21076 2315 21122
rect 2269 20968 2315 21014
rect 2269 20861 2315 20907
rect 2269 20754 2315 20800
rect 2269 20647 2315 20693
rect 2269 20540 2315 20586
rect 2269 20433 2315 20479
rect 2269 20326 2315 20372
rect 2665 21616 2711 21662
rect 2665 21508 2711 21554
rect 2665 21400 2711 21446
rect 2665 21292 2711 21338
rect 2665 21184 2711 21230
rect 2665 21076 2711 21122
rect 2665 20968 2711 21014
rect 2665 20861 2711 20907
rect 2665 20754 2711 20800
rect 2665 20647 2711 20693
rect 2665 20540 2711 20586
rect 2665 20433 2711 20479
rect 2665 20326 2711 20372
rect 2889 21616 2935 21662
rect 2889 21508 2935 21554
rect 2889 21400 2935 21446
rect 2889 21292 2935 21338
rect 2889 21184 2935 21230
rect 2889 21076 2935 21122
rect 2889 20968 2935 21014
rect 2889 20861 2935 20907
rect 2889 20754 2935 20800
rect 2889 20647 2935 20693
rect 2889 20540 2935 20586
rect 2889 20433 2935 20479
rect 2889 20326 2935 20372
rect 3283 21616 3329 21662
rect 3283 21508 3329 21554
rect 3283 21400 3329 21446
rect 3283 21292 3329 21338
rect 3283 21184 3329 21230
rect 3283 21076 3329 21122
rect 3283 20968 3329 21014
rect 3283 20861 3329 20907
rect 3283 20754 3329 20800
rect 3283 20647 3329 20693
rect 3283 20540 3329 20586
rect 3283 20433 3329 20479
rect 3283 20326 3329 20372
rect 3507 21616 3553 21662
rect 3507 21508 3553 21554
rect 3507 21400 3553 21446
rect 3507 21292 3553 21338
rect 3507 21184 3553 21230
rect 3507 21076 3553 21122
rect 3507 20968 3553 21014
rect 3507 20861 3553 20907
rect 3507 20754 3553 20800
rect 3507 20647 3553 20693
rect 3507 20540 3553 20586
rect 3507 20433 3553 20479
rect 3507 20326 3553 20372
rect 3903 21616 3949 21662
rect 3903 21508 3949 21554
rect 3903 21400 3949 21446
rect 3903 21292 3949 21338
rect 3903 21184 3949 21230
rect 3903 21076 3949 21122
rect 3903 20968 3949 21014
rect 3903 20861 3949 20907
rect 3903 20754 3949 20800
rect 3903 20647 3949 20693
rect 3903 20540 3949 20586
rect 3903 20433 3949 20479
rect 3903 20326 3949 20372
rect 4127 21616 4173 21662
rect 4127 21508 4173 21554
rect 4127 21400 4173 21446
rect 4127 21292 4173 21338
rect 4127 21184 4173 21230
rect 4127 21076 4173 21122
rect 4127 20968 4173 21014
rect 4127 20861 4173 20907
rect 4127 20754 4173 20800
rect 4127 20647 4173 20693
rect 4127 20540 4173 20586
rect 4127 20433 4173 20479
rect 4127 20326 4173 20372
rect 4522 21616 4568 21662
rect 4522 21508 4568 21554
rect 4522 21400 4568 21446
rect 4522 21292 4568 21338
rect 4522 21184 4568 21230
rect 4522 21076 4568 21122
rect 4522 20968 4568 21014
rect 4522 20861 4568 20907
rect 4522 20754 4568 20800
rect 4522 20647 4568 20693
rect 4522 20540 4568 20586
rect 4522 20433 4568 20479
rect 4522 20326 4568 20372
rect 4746 21616 4792 21662
rect 4746 21508 4792 21554
rect 4746 21400 4792 21446
rect 4746 21292 4792 21338
rect 4746 21184 4792 21230
rect 4746 21076 4792 21122
rect 4746 20968 4792 21014
rect 4746 20861 4792 20907
rect 4746 20754 4792 20800
rect 4746 20647 4792 20693
rect 4746 20540 4792 20586
rect 4746 20433 4792 20479
rect 4746 20326 4792 20372
rect 5142 21616 5188 21662
rect 5142 21508 5188 21554
rect 5142 21400 5188 21446
rect 5142 21292 5188 21338
rect 5142 21184 5188 21230
rect 5142 21076 5188 21122
rect 5142 20968 5188 21014
rect 5142 20861 5188 20907
rect 5142 20754 5188 20800
rect 5142 20647 5188 20693
rect 5142 20540 5188 20586
rect 5142 20433 5188 20479
rect 5142 20326 5188 20372
rect 5366 21616 5412 21662
rect 5366 21508 5412 21554
rect 5366 21400 5412 21446
rect 5366 21292 5412 21338
rect 5366 21184 5412 21230
rect 5366 21076 5412 21122
rect 5366 20968 5412 21014
rect 5366 20861 5412 20907
rect 5366 20754 5412 20800
rect 5366 20647 5412 20693
rect 5366 20540 5412 20586
rect 5366 20433 5412 20479
rect 5366 20326 5412 20372
rect 780 17177 826 17223
rect 1004 17177 1050 17223
rect 1228 17177 1274 17223
rect 1452 17177 1498 17223
rect 1676 17177 1722 17223
rect 2019 17177 2065 17223
rect 2243 17177 2289 17223
rect 2467 17177 2513 17223
rect 2691 17177 2737 17223
rect 2915 17177 2961 17223
rect 3257 17177 3303 17223
rect 3481 17177 3527 17223
rect 3705 17177 3751 17223
rect 3929 17177 3975 17223
rect 4153 17177 4199 17223
rect 4496 17177 4542 17223
rect 4720 17177 4766 17223
rect 4944 17177 4990 17223
rect 5168 17177 5214 17223
rect 5392 17177 5438 17223
rect 948 15545 994 15591
rect 1211 15545 1257 15591
rect 300 9911 346 12607
rect 524 9911 570 12607
rect 748 12560 794 12606
rect 748 12456 794 12502
rect 748 12352 794 12398
rect 748 12248 794 12294
rect 748 12144 794 12190
rect 748 12040 794 12086
rect 748 11936 794 11982
rect 748 11832 794 11878
rect 748 11728 794 11774
rect 748 11624 794 11670
rect 748 11519 794 11565
rect 748 11414 794 11460
rect 748 11309 794 11355
rect 748 11204 794 11250
rect 748 11099 794 11145
rect 748 10994 794 11040
rect 748 10889 794 10935
rect 748 10784 794 10830
rect 748 10679 794 10725
rect 748 10574 794 10620
rect 748 10469 794 10515
rect 748 10364 794 10410
rect 972 12560 1018 12606
rect 972 12456 1018 12502
rect 972 12352 1018 12398
rect 972 12248 1018 12294
rect 972 12144 1018 12190
rect 972 12040 1018 12086
rect 972 11936 1018 11982
rect 972 11832 1018 11878
rect 972 11728 1018 11774
rect 972 11624 1018 11670
rect 972 11519 1018 11565
rect 972 11414 1018 11460
rect 972 11309 1018 11355
rect 972 11204 1018 11250
rect 972 11099 1018 11145
rect 972 10994 1018 11040
rect 972 10889 1018 10935
rect 972 10784 1018 10830
rect 972 10679 1018 10725
rect 972 10574 1018 10620
rect 972 10469 1018 10515
rect 972 10364 1018 10410
rect 1196 12560 1242 12606
rect 1196 12456 1242 12502
rect 1196 12352 1242 12398
rect 1196 12248 1242 12294
rect 1196 12144 1242 12190
rect 1196 12040 1242 12086
rect 1196 11936 1242 11982
rect 1196 11832 1242 11878
rect 1196 11728 1242 11774
rect 1196 11624 1242 11670
rect 1196 11519 1242 11565
rect 1196 11414 1242 11460
rect 1196 11309 1242 11355
rect 1196 11204 1242 11250
rect 1196 11099 1242 11145
rect 1196 10994 1242 11040
rect 1196 10889 1242 10935
rect 1196 10784 1242 10830
rect 1196 10679 1242 10725
rect 1196 10574 1242 10620
rect 1196 10469 1242 10515
rect 1196 10364 1242 10410
rect 1420 12560 1466 12606
rect 1420 12456 1466 12502
rect 1420 12352 1466 12398
rect 1420 12248 1466 12294
rect 1420 12144 1466 12190
rect 1420 12040 1466 12086
rect 1420 11936 1466 11982
rect 1420 11832 1466 11878
rect 1420 11728 1466 11774
rect 1420 11624 1466 11670
rect 1420 11519 1466 11565
rect 1420 11414 1466 11460
rect 1420 11309 1466 11355
rect 1420 11204 1466 11250
rect 1420 11099 1466 11145
rect 1420 10994 1466 11040
rect 1420 10889 1466 10935
rect 1420 10784 1466 10830
rect 1420 10679 1466 10725
rect 1420 10574 1466 10620
rect 1420 10469 1466 10515
rect 1420 10364 1466 10410
rect 1644 12560 1690 12606
rect 1644 12456 1690 12502
rect 1644 12352 1690 12398
rect 1644 12248 1690 12294
rect 1644 12144 1690 12190
rect 1644 12040 1690 12086
rect 1644 11936 1690 11982
rect 1644 11832 1690 11878
rect 1644 11728 1690 11774
rect 1644 11624 1690 11670
rect 1644 11519 1690 11565
rect 1644 11414 1690 11460
rect 1644 11309 1690 11355
rect 1644 11204 1690 11250
rect 1644 11099 1690 11145
rect 1644 10994 1690 11040
rect 1644 10889 1690 10935
rect 1644 10784 1690 10830
rect 1644 10679 1690 10725
rect 1644 10574 1690 10620
rect 1644 10469 1690 10515
rect 1644 10364 1690 10410
rect 1868 12560 1914 12606
rect 1868 12456 1914 12502
rect 1868 12352 1914 12398
rect 1868 12248 1914 12294
rect 1868 12144 1914 12190
rect 1868 12040 1914 12086
rect 1868 11936 1914 11982
rect 1868 11832 1914 11878
rect 1868 11728 1914 11774
rect 1868 11624 1914 11670
rect 1868 11519 1914 11565
rect 1868 11414 1914 11460
rect 1868 11309 1914 11355
rect 1868 11204 1914 11250
rect 1868 11099 1914 11145
rect 1868 10994 1914 11040
rect 1868 10889 1914 10935
rect 1868 10784 1914 10830
rect 1868 10679 1914 10725
rect 1868 10574 1914 10620
rect 1868 10469 1914 10515
rect 1868 10364 1914 10410
rect 2481 9938 2527 9984
rect 1629 9852 1675 9898
rect 911 9752 957 9798
rect 911 9632 957 9678
rect 1135 9752 1181 9798
rect 1629 9732 1675 9778
rect 1853 9852 1899 9898
rect 1853 9732 1899 9778
rect 2481 9810 2527 9856
rect 1135 9632 1181 9678
rect 2481 9683 2527 9729
rect 2481 9556 2527 9602
rect 2705 9938 2751 9984
rect 2705 9810 2751 9856
rect 2705 9683 2751 9729
rect 2705 9556 2751 9602
rect 801 8111 847 8157
rect 801 7991 847 8037
rect 1025 8111 1071 8157
rect 1025 7991 1071 8037
rect 1249 8111 1295 8157
rect 1249 7991 1295 8037
rect 1629 8090 1675 8136
rect 1629 7970 1675 8016
rect 1853 8090 1899 8136
rect 1853 7970 1899 8016
rect 2077 8090 2123 8136
rect 2077 7970 2123 8016
rect 5562 208 5608 536
<< mvpdiffc >>
rect 692 28542 738 28588
rect 692 28360 738 28406
rect 692 28179 738 28225
rect 692 27997 738 28043
rect 918 28542 964 28588
rect 918 28360 964 28406
rect 918 28179 964 28225
rect 918 27997 964 28043
rect 1228 28542 1274 28588
rect 1228 28360 1274 28406
rect 1228 28179 1274 28225
rect 1228 27997 1274 28043
rect 1538 28542 1584 28588
rect 1538 28360 1584 28406
rect 1538 28179 1584 28225
rect 1538 27997 1584 28043
rect 1764 28542 1810 28588
rect 1931 28542 1977 28588
rect 1764 28360 1810 28406
rect 1931 28360 1977 28406
rect 1764 28179 1810 28225
rect 1931 28179 1977 28225
rect 1764 27997 1810 28043
rect 1931 27997 1977 28043
rect 2157 28542 2203 28588
rect 2157 28360 2203 28406
rect 2157 28179 2203 28225
rect 2157 27997 2203 28043
rect 2467 28542 2513 28588
rect 2467 28360 2513 28406
rect 2467 28179 2513 28225
rect 2467 27997 2513 28043
rect 2777 28542 2823 28588
rect 2777 28360 2823 28406
rect 2777 28179 2823 28225
rect 2777 27997 2823 28043
rect 3003 28542 3049 28588
rect 3169 28542 3215 28588
rect 3003 28360 3049 28406
rect 3169 28360 3215 28406
rect 3003 28179 3049 28225
rect 3169 28179 3215 28225
rect 3003 27997 3049 28043
rect 3169 27997 3215 28043
rect 3395 28542 3441 28588
rect 3395 28360 3441 28406
rect 3395 28179 3441 28225
rect 3395 27997 3441 28043
rect 3705 28542 3751 28588
rect 3705 28360 3751 28406
rect 3705 28179 3751 28225
rect 3705 27997 3751 28043
rect 4015 28542 4061 28588
rect 4015 28360 4061 28406
rect 4015 28179 4061 28225
rect 4015 27997 4061 28043
rect 4241 28542 4287 28588
rect 4408 28542 4454 28588
rect 4241 28360 4287 28406
rect 4408 28360 4454 28406
rect 4241 28179 4287 28225
rect 4408 28179 4454 28225
rect 4241 27997 4287 28043
rect 4408 27997 4454 28043
rect 4634 28542 4680 28588
rect 4634 28360 4680 28406
rect 4634 28179 4680 28225
rect 4634 27997 4680 28043
rect 4944 28542 4990 28588
rect 4944 28360 4990 28406
rect 4944 28179 4990 28225
rect 4944 27997 4990 28043
rect 5219 28542 5265 28588
rect 5219 28360 5265 28406
rect 5219 28179 5265 28225
rect 5219 27997 5265 28043
rect 5480 28542 5526 28588
rect 5480 28360 5526 28406
rect 5480 28179 5526 28225
rect 5480 27997 5526 28043
rect 692 27766 738 27812
rect 692 27585 738 27631
rect 692 27404 738 27450
rect 692 27222 738 27268
rect 918 27766 964 27812
rect 918 27585 964 27631
rect 918 27404 964 27450
rect 918 27222 964 27268
rect 1228 27766 1274 27812
rect 1228 27585 1274 27631
rect 1228 27404 1274 27450
rect 1228 27222 1274 27268
rect 1538 27766 1584 27812
rect 1538 27585 1584 27631
rect 1538 27404 1584 27450
rect 1538 27222 1584 27268
rect 1764 27766 1810 27812
rect 1931 27766 1977 27812
rect 1764 27585 1810 27631
rect 1931 27585 1977 27631
rect 1764 27404 1810 27450
rect 1931 27404 1977 27450
rect 1764 27222 1810 27268
rect 1931 27222 1977 27268
rect 2157 27766 2203 27812
rect 2157 27585 2203 27631
rect 2157 27404 2203 27450
rect 2157 27222 2203 27268
rect 2467 27766 2513 27812
rect 2467 27585 2513 27631
rect 2467 27404 2513 27450
rect 2467 27222 2513 27268
rect 2777 27766 2823 27812
rect 2777 27585 2823 27631
rect 2777 27404 2823 27450
rect 2777 27222 2823 27268
rect 3003 27766 3049 27812
rect 3169 27766 3215 27812
rect 3003 27585 3049 27631
rect 3169 27585 3215 27631
rect 3003 27404 3049 27450
rect 3169 27404 3215 27450
rect 3003 27222 3049 27268
rect 3169 27222 3215 27268
rect 3395 27766 3441 27812
rect 3395 27585 3441 27631
rect 3395 27404 3441 27450
rect 3395 27222 3441 27268
rect 3705 27766 3751 27812
rect 3705 27585 3751 27631
rect 3705 27404 3751 27450
rect 3705 27222 3751 27268
rect 4015 27766 4061 27812
rect 4015 27585 4061 27631
rect 4015 27404 4061 27450
rect 4015 27222 4061 27268
rect 4241 27766 4287 27812
rect 4408 27766 4454 27812
rect 4241 27585 4287 27631
rect 4408 27585 4454 27631
rect 4241 27404 4287 27450
rect 4408 27404 4454 27450
rect 4241 27222 4287 27268
rect 4408 27222 4454 27268
rect 4634 27766 4680 27812
rect 4634 27585 4680 27631
rect 4634 27404 4680 27450
rect 4634 27222 4680 27268
rect 4944 27766 4990 27812
rect 4944 27585 4990 27631
rect 4944 27404 4990 27450
rect 4944 27222 4990 27268
rect 5219 27766 5265 27812
rect 5219 27585 5265 27631
rect 5219 27404 5265 27450
rect 5219 27222 5265 27268
rect 5480 27766 5526 27812
rect 5480 27585 5526 27631
rect 5480 27404 5526 27450
rect 5480 27222 5526 27268
rect 808 26898 854 26944
rect 808 26790 854 26836
rect 808 26682 854 26728
rect 808 26574 854 26620
rect 808 26466 854 26512
rect 808 26358 854 26404
rect 808 26250 854 26296
rect 808 26143 854 26189
rect 808 26036 854 26082
rect 808 25929 854 25975
rect 808 25822 854 25868
rect 808 25715 854 25761
rect 808 25608 854 25654
rect 1032 26898 1078 26944
rect 1032 26790 1078 26836
rect 1032 26682 1078 26728
rect 1032 26574 1078 26620
rect 1032 26466 1078 26512
rect 1032 26358 1078 26404
rect 1032 26250 1078 26296
rect 1032 26143 1078 26189
rect 1032 26036 1078 26082
rect 1032 25929 1078 25975
rect 1032 25822 1078 25868
rect 1032 25715 1078 25761
rect 1032 25608 1078 25654
rect 1424 26898 1470 26944
rect 1424 26790 1470 26836
rect 1424 26682 1470 26728
rect 1424 26574 1470 26620
rect 1424 26466 1470 26512
rect 1424 26358 1470 26404
rect 1424 26250 1470 26296
rect 1424 26143 1470 26189
rect 1424 26036 1470 26082
rect 1424 25929 1470 25975
rect 1424 25822 1470 25868
rect 1424 25715 1470 25761
rect 1424 25608 1470 25654
rect 1648 26898 1694 26944
rect 1648 26790 1694 26836
rect 1648 26682 1694 26728
rect 1648 26574 1694 26620
rect 1648 26466 1694 26512
rect 1648 26358 1694 26404
rect 1648 26250 1694 26296
rect 1648 26143 1694 26189
rect 1648 26036 1694 26082
rect 1648 25929 1694 25975
rect 1648 25822 1694 25868
rect 1648 25715 1694 25761
rect 1648 25608 1694 25654
rect 2047 26898 2093 26944
rect 2047 26790 2093 26836
rect 2047 26682 2093 26728
rect 2047 26574 2093 26620
rect 2047 26466 2093 26512
rect 2047 26358 2093 26404
rect 2047 26250 2093 26296
rect 2047 26143 2093 26189
rect 2047 26036 2093 26082
rect 2047 25929 2093 25975
rect 2047 25822 2093 25868
rect 2047 25715 2093 25761
rect 2047 25608 2093 25654
rect 2271 26898 2317 26944
rect 2271 26790 2317 26836
rect 2271 26682 2317 26728
rect 2271 26574 2317 26620
rect 2271 26466 2317 26512
rect 2271 26358 2317 26404
rect 2271 26250 2317 26296
rect 2271 26143 2317 26189
rect 2271 26036 2317 26082
rect 2271 25929 2317 25975
rect 2271 25822 2317 25868
rect 2271 25715 2317 25761
rect 2271 25608 2317 25654
rect 2663 26898 2709 26944
rect 2663 26790 2709 26836
rect 2663 26682 2709 26728
rect 2663 26574 2709 26620
rect 2663 26466 2709 26512
rect 2663 26358 2709 26404
rect 2663 26250 2709 26296
rect 2663 26143 2709 26189
rect 2663 26036 2709 26082
rect 2663 25929 2709 25975
rect 2663 25822 2709 25868
rect 2663 25715 2709 25761
rect 2663 25608 2709 25654
rect 2887 26898 2933 26944
rect 2887 26790 2933 26836
rect 2887 26682 2933 26728
rect 2887 26574 2933 26620
rect 2887 26466 2933 26512
rect 2887 26358 2933 26404
rect 2887 26250 2933 26296
rect 2887 26143 2933 26189
rect 2887 26036 2933 26082
rect 2887 25929 2933 25975
rect 2887 25822 2933 25868
rect 2887 25715 2933 25761
rect 2887 25608 2933 25654
rect 3285 26898 3331 26944
rect 3285 26790 3331 26836
rect 3285 26682 3331 26728
rect 3285 26574 3331 26620
rect 3285 26466 3331 26512
rect 3285 26358 3331 26404
rect 3285 26250 3331 26296
rect 3285 26143 3331 26189
rect 3285 26036 3331 26082
rect 3285 25929 3331 25975
rect 3285 25822 3331 25868
rect 3285 25715 3331 25761
rect 3285 25608 3331 25654
rect 3509 26898 3555 26944
rect 3509 26790 3555 26836
rect 3509 26682 3555 26728
rect 3509 26574 3555 26620
rect 3509 26466 3555 26512
rect 3509 26358 3555 26404
rect 3509 26250 3555 26296
rect 3509 26143 3555 26189
rect 3509 26036 3555 26082
rect 3509 25929 3555 25975
rect 3509 25822 3555 25868
rect 3509 25715 3555 25761
rect 3509 25608 3555 25654
rect 3901 26898 3947 26944
rect 3901 26790 3947 26836
rect 3901 26682 3947 26728
rect 3901 26574 3947 26620
rect 3901 26466 3947 26512
rect 3901 26358 3947 26404
rect 3901 26250 3947 26296
rect 3901 26143 3947 26189
rect 3901 26036 3947 26082
rect 3901 25929 3947 25975
rect 3901 25822 3947 25868
rect 3901 25715 3947 25761
rect 3901 25608 3947 25654
rect 4125 26898 4171 26944
rect 4125 26790 4171 26836
rect 4125 26682 4171 26728
rect 4125 26574 4171 26620
rect 4125 26466 4171 26512
rect 4125 26358 4171 26404
rect 4125 26250 4171 26296
rect 4125 26143 4171 26189
rect 4125 26036 4171 26082
rect 4125 25929 4171 25975
rect 4125 25822 4171 25868
rect 4125 25715 4171 25761
rect 4125 25608 4171 25654
rect 4524 26898 4570 26944
rect 4524 26790 4570 26836
rect 4524 26682 4570 26728
rect 4524 26574 4570 26620
rect 4524 26466 4570 26512
rect 4524 26358 4570 26404
rect 4524 26250 4570 26296
rect 4524 26143 4570 26189
rect 4524 26036 4570 26082
rect 4524 25929 4570 25975
rect 4524 25822 4570 25868
rect 4524 25715 4570 25761
rect 4524 25608 4570 25654
rect 4748 26898 4794 26944
rect 4748 26790 4794 26836
rect 4748 26682 4794 26728
rect 4748 26574 4794 26620
rect 4748 26466 4794 26512
rect 4748 26358 4794 26404
rect 4748 26250 4794 26296
rect 4748 26143 4794 26189
rect 4748 26036 4794 26082
rect 4748 25929 4794 25975
rect 4748 25822 4794 25868
rect 4748 25715 4794 25761
rect 4748 25608 4794 25654
rect 5140 26898 5186 26944
rect 5140 26790 5186 26836
rect 5140 26682 5186 26728
rect 5140 26574 5186 26620
rect 5140 26466 5186 26512
rect 5140 26358 5186 26404
rect 5140 26250 5186 26296
rect 5140 26143 5186 26189
rect 5140 26036 5186 26082
rect 5140 25929 5186 25975
rect 5140 25822 5186 25868
rect 5140 25715 5186 25761
rect 5140 25608 5186 25654
rect 5364 26898 5410 26944
rect 5364 26790 5410 26836
rect 5364 26682 5410 26728
rect 5364 26574 5410 26620
rect 5364 26466 5410 26512
rect 5364 26358 5410 26404
rect 5364 26250 5410 26296
rect 5364 26143 5410 26189
rect 5364 26036 5410 26082
rect 5364 25929 5410 25975
rect 5364 25822 5410 25868
rect 5364 25715 5410 25761
rect 5364 25608 5410 25654
rect 806 25311 852 25357
rect 806 25203 852 25249
rect 806 25095 852 25141
rect 806 24987 852 25033
rect 806 24879 852 24925
rect 806 24771 852 24817
rect 806 24663 852 24709
rect 806 24556 852 24602
rect 806 24449 852 24495
rect 806 24342 852 24388
rect 806 24235 852 24281
rect 806 24128 852 24174
rect 806 24021 852 24067
rect 1030 25311 1076 25357
rect 1030 25203 1076 25249
rect 1030 25095 1076 25141
rect 1030 24987 1076 25033
rect 1030 24879 1076 24925
rect 1030 24771 1076 24817
rect 1030 24663 1076 24709
rect 1426 25311 1472 25357
rect 1426 25203 1472 25249
rect 1426 25095 1472 25141
rect 1426 24987 1472 25033
rect 1426 24879 1472 24925
rect 1426 24771 1472 24817
rect 1030 24556 1076 24602
rect 1030 24449 1076 24495
rect 1426 24663 1472 24709
rect 1426 24556 1472 24602
rect 1426 24449 1472 24495
rect 1030 24342 1076 24388
rect 1030 24235 1076 24281
rect 1030 24128 1076 24174
rect 1030 24021 1076 24067
rect 1426 24342 1472 24388
rect 1426 24235 1472 24281
rect 1426 24128 1472 24174
rect 1426 24021 1472 24067
rect 1650 25311 1696 25357
rect 1650 25203 1696 25249
rect 1650 25095 1696 25141
rect 1650 24987 1696 25033
rect 1650 24879 1696 24925
rect 1650 24771 1696 24817
rect 1650 24663 1696 24709
rect 1650 24556 1696 24602
rect 1650 24449 1696 24495
rect 1650 24342 1696 24388
rect 1650 24235 1696 24281
rect 1650 24128 1696 24174
rect 1650 24021 1696 24067
rect 2045 25311 2091 25357
rect 2045 25203 2091 25249
rect 2045 25095 2091 25141
rect 2045 24987 2091 25033
rect 2045 24879 2091 24925
rect 2045 24771 2091 24817
rect 2045 24663 2091 24709
rect 2045 24556 2091 24602
rect 2045 24449 2091 24495
rect 2045 24342 2091 24388
rect 2045 24235 2091 24281
rect 2045 24128 2091 24174
rect 2045 24021 2091 24067
rect 2269 25311 2315 25357
rect 2269 25203 2315 25249
rect 2269 25095 2315 25141
rect 2269 24987 2315 25033
rect 2269 24879 2315 24925
rect 2269 24771 2315 24817
rect 2269 24663 2315 24709
rect 2665 25311 2711 25357
rect 2665 25203 2711 25249
rect 2665 25095 2711 25141
rect 2665 24987 2711 25033
rect 2665 24879 2711 24925
rect 2665 24771 2711 24817
rect 2269 24556 2315 24602
rect 2269 24449 2315 24495
rect 2665 24663 2711 24709
rect 2665 24556 2711 24602
rect 2665 24449 2711 24495
rect 2269 24342 2315 24388
rect 2269 24235 2315 24281
rect 2269 24128 2315 24174
rect 2269 24021 2315 24067
rect 2665 24342 2711 24388
rect 2665 24235 2711 24281
rect 2665 24128 2711 24174
rect 2665 24021 2711 24067
rect 2889 25311 2935 25357
rect 2889 25203 2935 25249
rect 2889 25095 2935 25141
rect 2889 24987 2935 25033
rect 2889 24879 2935 24925
rect 2889 24771 2935 24817
rect 2889 24663 2935 24709
rect 2889 24556 2935 24602
rect 2889 24449 2935 24495
rect 2889 24342 2935 24388
rect 2889 24235 2935 24281
rect 2889 24128 2935 24174
rect 2889 24021 2935 24067
rect 3283 25311 3329 25357
rect 3283 25203 3329 25249
rect 3283 25095 3329 25141
rect 3283 24987 3329 25033
rect 3283 24879 3329 24925
rect 3283 24771 3329 24817
rect 3283 24663 3329 24709
rect 3283 24556 3329 24602
rect 3283 24449 3329 24495
rect 3283 24342 3329 24388
rect 3283 24235 3329 24281
rect 3283 24128 3329 24174
rect 3283 24021 3329 24067
rect 3507 25311 3553 25357
rect 3507 25203 3553 25249
rect 3507 25095 3553 25141
rect 3507 24987 3553 25033
rect 3507 24879 3553 24925
rect 3507 24771 3553 24817
rect 3507 24663 3553 24709
rect 3903 25311 3949 25357
rect 3903 25203 3949 25249
rect 3903 25095 3949 25141
rect 3903 24987 3949 25033
rect 3903 24879 3949 24925
rect 3903 24771 3949 24817
rect 3507 24556 3553 24602
rect 3507 24449 3553 24495
rect 3903 24663 3949 24709
rect 3903 24556 3949 24602
rect 3903 24449 3949 24495
rect 3507 24342 3553 24388
rect 3507 24235 3553 24281
rect 3507 24128 3553 24174
rect 3507 24021 3553 24067
rect 3903 24342 3949 24388
rect 3903 24235 3949 24281
rect 3903 24128 3949 24174
rect 3903 24021 3949 24067
rect 4127 25311 4173 25357
rect 4127 25203 4173 25249
rect 4127 25095 4173 25141
rect 4127 24987 4173 25033
rect 4127 24879 4173 24925
rect 4127 24771 4173 24817
rect 4127 24663 4173 24709
rect 4127 24556 4173 24602
rect 4127 24449 4173 24495
rect 4127 24342 4173 24388
rect 4127 24235 4173 24281
rect 4127 24128 4173 24174
rect 4127 24021 4173 24067
rect 4522 25311 4568 25357
rect 4522 25203 4568 25249
rect 4522 25095 4568 25141
rect 4522 24987 4568 25033
rect 4522 24879 4568 24925
rect 4522 24771 4568 24817
rect 4522 24663 4568 24709
rect 4522 24556 4568 24602
rect 4522 24449 4568 24495
rect 4522 24342 4568 24388
rect 4522 24235 4568 24281
rect 4522 24128 4568 24174
rect 4522 24021 4568 24067
rect 4746 25311 4792 25357
rect 4746 25203 4792 25249
rect 4746 25095 4792 25141
rect 4746 24987 4792 25033
rect 4746 24879 4792 24925
rect 4746 24771 4792 24817
rect 4746 24663 4792 24709
rect 5142 25311 5188 25357
rect 5142 25203 5188 25249
rect 5142 25095 5188 25141
rect 5142 24987 5188 25033
rect 5142 24879 5188 24925
rect 5142 24771 5188 24817
rect 4746 24556 4792 24602
rect 4746 24449 4792 24495
rect 5142 24663 5188 24709
rect 5142 24556 5188 24602
rect 5142 24449 5188 24495
rect 4746 24342 4792 24388
rect 4746 24235 4792 24281
rect 4746 24128 4792 24174
rect 4746 24021 4792 24067
rect 5142 24342 5188 24388
rect 5142 24235 5188 24281
rect 5142 24128 5188 24174
rect 5142 24021 5188 24067
rect 5366 25311 5412 25357
rect 5366 25203 5412 25249
rect 5366 25095 5412 25141
rect 5366 24987 5412 25033
rect 5366 24879 5412 24925
rect 5366 24771 5412 24817
rect 5366 24663 5412 24709
rect 5366 24556 5412 24602
rect 5366 24449 5412 24495
rect 5366 24342 5412 24388
rect 5366 24235 5412 24281
rect 5366 24128 5412 24174
rect 5366 24021 5412 24067
rect 806 19761 852 19807
rect 806 19653 852 19699
rect 806 19545 852 19591
rect 806 19437 852 19483
rect 806 19329 852 19375
rect 806 19221 852 19267
rect 806 19113 852 19159
rect 806 19006 852 19052
rect 806 18899 852 18945
rect 806 18792 852 18838
rect 806 18685 852 18731
rect 806 18578 852 18624
rect 806 18471 852 18517
rect 1030 19761 1076 19807
rect 1030 19653 1076 19699
rect 1030 19545 1076 19591
rect 1030 19437 1076 19483
rect 1030 19329 1076 19375
rect 1030 19221 1076 19267
rect 1030 19113 1076 19159
rect 1030 19006 1076 19052
rect 1030 18899 1076 18945
rect 1030 18792 1076 18838
rect 1030 18685 1076 18731
rect 1030 18578 1076 18624
rect 1030 18471 1076 18517
rect 1426 19761 1472 19807
rect 1426 19653 1472 19699
rect 1426 19545 1472 19591
rect 1426 19437 1472 19483
rect 1426 19329 1472 19375
rect 1426 19221 1472 19267
rect 1426 19113 1472 19159
rect 1426 19006 1472 19052
rect 1426 18899 1472 18945
rect 1426 18792 1472 18838
rect 1426 18685 1472 18731
rect 1426 18578 1472 18624
rect 1426 18471 1472 18517
rect 1650 19761 1696 19807
rect 1650 19653 1696 19699
rect 1650 19545 1696 19591
rect 1650 19437 1696 19483
rect 1650 19329 1696 19375
rect 1650 19221 1696 19267
rect 1650 19113 1696 19159
rect 1650 19006 1696 19052
rect 1650 18899 1696 18945
rect 1650 18792 1696 18838
rect 1650 18685 1696 18731
rect 1650 18578 1696 18624
rect 1650 18471 1696 18517
rect 2045 19761 2091 19807
rect 2045 19653 2091 19699
rect 2045 19545 2091 19591
rect 2045 19437 2091 19483
rect 2045 19329 2091 19375
rect 2045 19221 2091 19267
rect 2045 19113 2091 19159
rect 2045 19006 2091 19052
rect 2045 18899 2091 18945
rect 2045 18792 2091 18838
rect 2045 18685 2091 18731
rect 2045 18578 2091 18624
rect 2045 18471 2091 18517
rect 2269 19761 2315 19807
rect 2269 19653 2315 19699
rect 2269 19545 2315 19591
rect 2269 19437 2315 19483
rect 2269 19329 2315 19375
rect 2269 19221 2315 19267
rect 2269 19113 2315 19159
rect 2269 19006 2315 19052
rect 2269 18899 2315 18945
rect 2269 18792 2315 18838
rect 2269 18685 2315 18731
rect 2269 18578 2315 18624
rect 2269 18471 2315 18517
rect 2665 19761 2711 19807
rect 2665 19653 2711 19699
rect 2665 19545 2711 19591
rect 2665 19437 2711 19483
rect 2665 19329 2711 19375
rect 2665 19221 2711 19267
rect 2665 19113 2711 19159
rect 2665 19006 2711 19052
rect 2665 18899 2711 18945
rect 2665 18792 2711 18838
rect 2665 18685 2711 18731
rect 2665 18578 2711 18624
rect 2665 18471 2711 18517
rect 2889 19761 2935 19807
rect 2889 19653 2935 19699
rect 2889 19545 2935 19591
rect 2889 19437 2935 19483
rect 2889 19329 2935 19375
rect 2889 19221 2935 19267
rect 2889 19113 2935 19159
rect 2889 19006 2935 19052
rect 2889 18899 2935 18945
rect 2889 18792 2935 18838
rect 2889 18685 2935 18731
rect 2889 18578 2935 18624
rect 2889 18471 2935 18517
rect 3283 19761 3329 19807
rect 3283 19653 3329 19699
rect 3283 19545 3329 19591
rect 3283 19437 3329 19483
rect 3283 19329 3329 19375
rect 3283 19221 3329 19267
rect 3283 19113 3329 19159
rect 3283 19006 3329 19052
rect 3283 18899 3329 18945
rect 3283 18792 3329 18838
rect 3283 18685 3329 18731
rect 3283 18578 3329 18624
rect 3283 18471 3329 18517
rect 3507 19761 3553 19807
rect 3507 19653 3553 19699
rect 3507 19545 3553 19591
rect 3507 19437 3553 19483
rect 3507 19329 3553 19375
rect 3507 19221 3553 19267
rect 3507 19113 3553 19159
rect 3507 19006 3553 19052
rect 3507 18899 3553 18945
rect 3507 18792 3553 18838
rect 3507 18685 3553 18731
rect 3507 18578 3553 18624
rect 3507 18471 3553 18517
rect 3903 19761 3949 19807
rect 3903 19653 3949 19699
rect 3903 19545 3949 19591
rect 3903 19437 3949 19483
rect 3903 19329 3949 19375
rect 3903 19221 3949 19267
rect 3903 19113 3949 19159
rect 3903 19006 3949 19052
rect 3903 18899 3949 18945
rect 3903 18792 3949 18838
rect 3903 18685 3949 18731
rect 3903 18578 3949 18624
rect 3903 18471 3949 18517
rect 4127 19761 4173 19807
rect 4127 19653 4173 19699
rect 4127 19545 4173 19591
rect 4127 19437 4173 19483
rect 4127 19329 4173 19375
rect 4127 19221 4173 19267
rect 4127 19113 4173 19159
rect 4127 19006 4173 19052
rect 4127 18899 4173 18945
rect 4127 18792 4173 18838
rect 4127 18685 4173 18731
rect 4127 18578 4173 18624
rect 4127 18471 4173 18517
rect 4522 19761 4568 19807
rect 4522 19653 4568 19699
rect 4522 19545 4568 19591
rect 4522 19437 4568 19483
rect 4522 19329 4568 19375
rect 4522 19221 4568 19267
rect 4522 19113 4568 19159
rect 4522 19006 4568 19052
rect 4522 18899 4568 18945
rect 4522 18792 4568 18838
rect 4522 18685 4568 18731
rect 4522 18578 4568 18624
rect 4522 18471 4568 18517
rect 4746 19761 4792 19807
rect 4746 19653 4792 19699
rect 4746 19545 4792 19591
rect 4746 19437 4792 19483
rect 4746 19329 4792 19375
rect 4746 19221 4792 19267
rect 4746 19113 4792 19159
rect 4746 19006 4792 19052
rect 4746 18899 4792 18945
rect 4746 18792 4792 18838
rect 4746 18685 4792 18731
rect 4746 18578 4792 18624
rect 4746 18471 4792 18517
rect 5142 19761 5188 19807
rect 5142 19653 5188 19699
rect 5142 19545 5188 19591
rect 5142 19437 5188 19483
rect 5142 19329 5188 19375
rect 5142 19221 5188 19267
rect 5142 19113 5188 19159
rect 5142 19006 5188 19052
rect 5142 18899 5188 18945
rect 5142 18792 5188 18838
rect 5142 18685 5188 18731
rect 5142 18578 5188 18624
rect 5142 18471 5188 18517
rect 5366 19761 5412 19807
rect 5366 19653 5412 19699
rect 5366 19545 5412 19591
rect 5366 19437 5412 19483
rect 5366 19329 5412 19375
rect 5366 19221 5412 19267
rect 5366 19113 5412 19159
rect 5366 19006 5412 19052
rect 5366 18899 5412 18945
rect 5366 18792 5412 18838
rect 5366 18685 5412 18731
rect 5366 18578 5412 18624
rect 5366 18471 5412 18517
rect 725 17674 771 17720
rect 975 17674 1021 17720
rect 1228 17674 1274 17720
rect 1481 17674 1527 17720
rect 1731 17674 1777 17720
rect 1964 17674 2010 17720
rect 2214 17674 2260 17720
rect 2467 17674 2513 17720
rect 2720 17674 2766 17720
rect 2970 17674 3016 17720
rect 3202 17674 3248 17720
rect 3452 17674 3498 17720
rect 3705 17674 3751 17720
rect 3958 17674 4004 17720
rect 4208 17674 4254 17720
rect 4441 17674 4487 17720
rect 4691 17674 4737 17720
rect 4944 17674 4990 17720
rect 5197 17674 5243 17720
rect 5447 17674 5493 17720
rect 300 13069 346 15765
rect 524 13069 570 15765
rect 1644 15265 1690 15311
rect 853 15026 899 15072
rect 1117 15026 1163 15072
rect 1350 15026 1396 15072
rect 1644 15161 1690 15207
rect 1644 15057 1690 15103
rect 1644 14953 1690 14999
rect 1644 14849 1690 14895
rect 1644 14745 1690 14791
rect 1644 14641 1690 14687
rect 1644 14537 1690 14583
rect 1644 14433 1690 14479
rect 748 14359 794 14405
rect 748 14252 794 14298
rect 748 14145 794 14191
rect 748 14038 794 14084
rect 748 13931 794 13977
rect 748 13824 794 13870
rect 748 13717 794 13763
rect 748 13609 794 13655
rect 748 13501 794 13547
rect 748 13393 794 13439
rect 748 13285 794 13331
rect 748 13177 794 13223
rect 748 13069 794 13115
rect 972 14359 1018 14405
rect 972 14252 1018 14298
rect 972 14145 1018 14191
rect 972 14038 1018 14084
rect 972 13931 1018 13977
rect 972 13824 1018 13870
rect 972 13717 1018 13763
rect 972 13609 1018 13655
rect 972 13501 1018 13547
rect 972 13393 1018 13439
rect 972 13285 1018 13331
rect 972 13177 1018 13223
rect 972 13069 1018 13115
rect 1196 14359 1242 14405
rect 1196 14252 1242 14298
rect 1196 14145 1242 14191
rect 1196 14038 1242 14084
rect 1196 13931 1242 13977
rect 1196 13824 1242 13870
rect 1196 13717 1242 13763
rect 1196 13609 1242 13655
rect 1196 13501 1242 13547
rect 1196 13393 1242 13439
rect 1196 13285 1242 13331
rect 1196 13177 1242 13223
rect 1196 13069 1242 13115
rect 1420 14359 1466 14405
rect 1420 14252 1466 14298
rect 1420 14145 1466 14191
rect 1420 14038 1466 14084
rect 1420 13931 1466 13977
rect 1420 13824 1466 13870
rect 1420 13717 1466 13763
rect 1420 13609 1466 13655
rect 1420 13501 1466 13547
rect 1420 13393 1466 13439
rect 1420 13285 1466 13331
rect 1420 13177 1466 13223
rect 1420 13069 1466 13115
rect 1644 14329 1690 14375
rect 1644 14224 1690 14270
rect 1644 14119 1690 14165
rect 1644 14014 1690 14060
rect 1644 13909 1690 13955
rect 1644 13804 1690 13850
rect 1644 13699 1690 13745
rect 1644 13594 1690 13640
rect 1644 13489 1690 13535
rect 1644 13384 1690 13430
rect 1644 13279 1690 13325
rect 1644 13174 1690 13220
rect 1644 13069 1690 13115
rect 1868 15265 1914 15311
rect 1868 15161 1914 15207
rect 1868 15057 1914 15103
rect 1868 14953 1914 14999
rect 1868 14849 1914 14895
rect 1868 14745 1914 14791
rect 1868 14641 1914 14687
rect 1868 14537 1914 14583
rect 1868 14433 1914 14479
rect 1868 14329 1914 14375
rect 1868 14224 1914 14270
rect 1868 14119 1914 14165
rect 1868 14014 1914 14060
rect 1868 13909 1914 13955
rect 1868 13804 1914 13850
rect 1868 13699 1914 13745
rect 1868 13594 1914 13640
rect 1868 13489 1914 13535
rect 1868 13384 1914 13430
rect 1868 13279 1914 13325
rect 1868 13174 1914 13220
rect 1868 13069 1914 13115
rect 1629 9381 1675 9427
rect 801 9188 847 9234
rect 801 9032 847 9078
rect 1025 9188 1071 9234
rect 1025 9032 1071 9078
rect 1249 9188 1295 9234
rect 1629 9225 1675 9271
rect 1853 9381 1899 9427
rect 1853 9225 1899 9271
rect 2077 9381 2123 9427
rect 2077 9225 2123 9271
rect 2481 9206 2527 9252
rect 1249 9032 1295 9078
rect 2481 9099 2527 9145
rect 2481 8992 2527 9038
rect 2481 8885 2527 8931
rect 2481 8778 2527 8824
rect 1629 8666 1675 8712
rect 801 8584 847 8630
rect 801 8464 847 8510
rect 1025 8584 1071 8630
rect 1025 8464 1071 8510
rect 1249 8584 1295 8630
rect 1629 8546 1675 8592
rect 1853 8666 1899 8712
rect 1853 8546 1899 8592
rect 2077 8666 2123 8712
rect 2077 8546 2123 8592
rect 2481 8671 2527 8717
rect 2481 8564 2527 8610
rect 1249 8464 1295 8510
rect 2481 8456 2527 8502
rect 2481 8348 2527 8394
rect 2481 8240 2527 8286
rect 2481 8132 2527 8178
rect 2481 8024 2527 8070
rect 2481 7916 2527 7962
rect 2705 9206 2751 9252
rect 2705 9099 2751 9145
rect 2705 8992 2751 9038
rect 2705 8885 2751 8931
rect 2705 8778 2751 8824
rect 2705 8671 2751 8717
rect 2705 8564 2751 8610
rect 2705 8456 2751 8502
rect 2705 8348 2751 8394
rect 2705 8240 2751 8286
rect 2705 8132 2751 8178
rect 2705 8024 2751 8070
rect 2705 7916 2751 7962
<< mvpsubdiff >>
rect 1171 22020 1331 22080
rect 1171 21974 1228 22020
rect 1274 21974 1331 22020
rect 1171 21914 1331 21974
rect 2410 22020 2570 22080
rect 2410 21974 2467 22020
rect 2513 21974 2570 22020
rect 2410 21914 2570 21974
rect 3648 22020 3808 22080
rect 3648 21974 3705 22020
rect 3751 21974 3808 22020
rect 3648 21914 3808 21974
rect 4887 22020 5047 22080
rect 4887 21974 4944 22020
rect 4990 21974 5047 22020
rect 4887 21914 5047 21974
rect 5507 22020 5667 22080
rect 5507 21974 5564 22020
rect 5610 21974 5667 22020
rect 5507 21914 5667 21974
rect 502 17252 586 17271
rect 502 17112 521 17252
rect 567 17112 586 17252
rect 1829 17252 1913 17271
rect 502 17093 586 17112
rect 1829 17112 1848 17252
rect 1894 17112 1913 17252
rect 3068 17252 3152 17271
rect 1829 17093 1913 17112
rect 3068 17112 3087 17252
rect 3133 17112 3152 17252
rect 4306 17252 4390 17271
rect 3068 17093 3152 17112
rect 4306 17112 4325 17252
rect 4371 17112 4390 17252
rect 5545 17252 5629 17271
rect 4306 17093 4390 17112
rect 5545 17112 5564 17252
rect 5610 17112 5629 17252
rect 5545 17093 5629 17112
rect 631 16856 5587 16915
rect 631 16810 754 16856
rect 800 16810 912 16856
rect 958 16810 1070 16856
rect 1116 16810 1228 16856
rect 1274 16810 1386 16856
rect 1432 16810 1544 16856
rect 1590 16810 1702 16856
rect 1748 16810 1993 16856
rect 2039 16810 2151 16856
rect 2197 16810 2309 16856
rect 2355 16810 2467 16856
rect 2513 16810 2625 16856
rect 2671 16810 2783 16856
rect 2829 16810 2941 16856
rect 2987 16810 3231 16856
rect 3277 16810 3389 16856
rect 3435 16810 3547 16856
rect 3593 16810 3705 16856
rect 3751 16810 3863 16856
rect 3909 16810 4021 16856
rect 4067 16810 4179 16856
rect 4225 16810 4470 16856
rect 4516 16810 4628 16856
rect 4674 16810 4786 16856
rect 4832 16810 4944 16856
rect 4990 16810 5102 16856
rect 5148 16810 5260 16856
rect 5306 16810 5418 16856
rect 5464 16810 5587 16856
rect 631 16750 5587 16810
rect 2309 15509 2469 15568
rect 2309 15463 2366 15509
rect 2412 15463 2469 15509
rect 2309 15345 2469 15463
rect 2309 15299 2366 15345
rect 2412 15299 2469 15345
rect 2309 15182 2469 15299
rect 2309 15136 2366 15182
rect 2412 15136 2469 15182
rect 2309 15019 2469 15136
rect 2309 14973 2366 15019
rect 2412 14973 2469 15019
rect 2309 14856 2469 14973
rect 2309 14810 2366 14856
rect 2412 14810 2469 14856
rect 2309 14693 2469 14810
rect 2309 14647 2366 14693
rect 2412 14647 2469 14693
rect 2309 14529 2469 14647
rect 2309 14483 2366 14529
rect 2412 14483 2469 14529
rect 2309 14366 2469 14483
rect 2309 14320 2366 14366
rect 2412 14320 2469 14366
rect 2309 14203 2469 14320
rect 2309 14157 2366 14203
rect 2412 14157 2469 14203
rect 2309 14040 2469 14157
rect 2309 13994 2366 14040
rect 2412 13994 2469 14040
rect 2309 13876 2469 13994
rect 2309 13830 2366 13876
rect 2412 13830 2469 13876
rect 2309 13713 2469 13830
rect 2309 13667 2366 13713
rect 2412 13667 2469 13713
rect 2309 13550 2469 13667
rect 2309 13504 2366 13550
rect 2412 13504 2469 13550
rect 2309 13387 2469 13504
rect 2309 13341 2366 13387
rect 2412 13341 2469 13387
rect 2309 13223 2469 13341
rect 2309 13177 2366 13223
rect 2412 13177 2469 13223
rect 2309 13060 2469 13177
rect 2309 13014 2366 13060
rect 2412 13014 2469 13060
rect 2309 12897 2469 13014
rect 2309 12851 2366 12897
rect 2412 12851 2469 12897
rect 2309 12733 2469 12851
rect 2309 12687 2366 12733
rect 2412 12687 2469 12733
rect 2309 12630 2469 12687
rect 2151 12571 2469 12630
rect 2151 12525 2208 12571
rect 2254 12570 2469 12571
rect 2254 12525 2366 12570
rect 2151 12524 2366 12525
rect 2412 12524 2469 12570
rect 2151 12407 2469 12524
rect 2151 12361 2208 12407
rect 2254 12361 2366 12407
rect 2412 12361 2469 12407
rect 2151 12244 2469 12361
rect 2151 12198 2208 12244
rect 2254 12198 2366 12244
rect 2412 12198 2469 12244
rect 2151 12081 2469 12198
rect 2151 12035 2208 12081
rect 2254 12080 2469 12081
rect 2254 12035 2366 12080
rect 2151 12034 2366 12035
rect 2412 12034 2469 12080
rect 2151 11918 2469 12034
rect 2151 11872 2208 11918
rect 2254 11917 2469 11918
rect 2254 11872 2366 11917
rect 2151 11871 2366 11872
rect 2412 11871 2469 11917
rect 2151 11754 2469 11871
rect 2151 11708 2208 11754
rect 2254 11708 2366 11754
rect 2412 11708 2469 11754
rect 2151 11591 2469 11708
rect 2151 11545 2208 11591
rect 2254 11545 2366 11591
rect 2412 11545 2469 11591
rect 2151 11428 2469 11545
rect 2151 11382 2208 11428
rect 2254 11427 2469 11428
rect 2254 11382 2366 11427
rect 2151 11381 2366 11382
rect 2412 11381 2469 11427
rect 2151 11264 2469 11381
rect 2151 11218 2208 11264
rect 2254 11218 2366 11264
rect 2412 11218 2469 11264
rect 2151 11101 2469 11218
rect 2151 11055 2208 11101
rect 2254 11055 2366 11101
rect 2412 11055 2469 11101
rect 2151 10938 2469 11055
rect 2151 10892 2208 10938
rect 2254 10892 2366 10938
rect 2412 10892 2469 10938
rect 2151 10775 2469 10892
rect 2151 10729 2208 10775
rect 2254 10729 2366 10775
rect 2412 10729 2469 10775
rect 2151 10611 2469 10729
rect 2151 10565 2208 10611
rect 2254 10565 2366 10611
rect 2412 10565 2469 10611
rect 2151 10507 2469 10565
rect 243 9526 403 9586
rect 243 9480 300 9526
rect 346 9480 403 9526
rect 243 9420 403 9480
rect 314 8131 398 8150
rect 314 7991 333 8131
rect 379 7991 398 8131
rect 314 7972 398 7991
<< mvnsubdiff >>
rect 601 28925 5618 28982
rect 601 28879 760 28925
rect 806 28879 918 28925
rect 964 28879 1076 28925
rect 1122 28879 1380 28925
rect 1426 28879 1538 28925
rect 1584 28879 1696 28925
rect 1742 28879 1999 28925
rect 2045 28879 2157 28925
rect 2203 28879 2315 28925
rect 2361 28879 2619 28925
rect 2665 28879 2777 28925
rect 2823 28879 2935 28925
rect 2981 28879 3237 28925
rect 3283 28879 3395 28925
rect 3441 28879 3553 28925
rect 3599 28879 3857 28925
rect 3903 28879 4015 28925
rect 4061 28879 4173 28925
rect 4219 28879 4476 28925
rect 4522 28879 4634 28925
rect 4680 28879 4792 28925
rect 4838 28879 5096 28925
rect 5142 28879 5254 28925
rect 5300 28879 5412 28925
rect 5458 28879 5618 28925
rect 601 28822 5618 28879
rect 1209 24657 1293 24676
rect 1209 24423 1228 24657
rect 1274 24423 1293 24657
rect 1209 24404 1293 24423
rect 2448 24657 2532 24676
rect 2448 24423 2467 24657
rect 2513 24423 2532 24657
rect 2448 24404 2532 24423
rect 3686 24657 3770 24676
rect 3686 24423 3705 24657
rect 3751 24423 3770 24657
rect 3686 24404 3770 24423
rect 4925 24657 5009 24676
rect 4925 24423 4944 24657
rect 4990 24423 5009 24657
rect 4925 24404 5009 24423
rect 631 18175 5587 18232
rect 631 18129 754 18175
rect 800 18129 912 18175
rect 958 18129 1070 18175
rect 1116 18129 1228 18175
rect 1274 18129 1386 18175
rect 1432 18129 1544 18175
rect 1590 18129 1702 18175
rect 1748 18129 1993 18175
rect 2039 18129 2151 18175
rect 2197 18129 2309 18175
rect 2355 18129 2467 18175
rect 2513 18129 2625 18175
rect 2671 18129 2783 18175
rect 2829 18129 2941 18175
rect 2987 18129 3231 18175
rect 3277 18129 3389 18175
rect 3435 18129 3547 18175
rect 3593 18129 3705 18175
rect 3751 18129 3863 18175
rect 3909 18129 4021 18175
rect 4067 18129 4179 18175
rect 4225 18129 4470 18175
rect 4516 18129 4628 18175
rect 4674 18129 4786 18175
rect 4832 18129 4944 18175
rect 4990 18129 5102 18175
rect 5148 18129 5260 18175
rect 5306 18129 5418 18175
rect 5464 18129 5587 18175
rect 631 18072 5587 18129
rect 1646 15562 1918 15581
rect 1646 15516 1665 15562
rect 1899 15516 1918 15562
rect 1646 15497 1918 15516
rect 245 8978 401 9035
rect 245 8932 300 8978
rect 346 8932 401 8978
rect 245 8814 401 8932
rect 245 8768 300 8814
rect 346 8768 401 8814
rect 245 8711 401 8768
<< mvpsubdiffcont >>
rect 1228 21974 1274 22020
rect 2467 21974 2513 22020
rect 3705 21974 3751 22020
rect 4944 21974 4990 22020
rect 5564 21974 5610 22020
rect 521 17112 567 17252
rect 1848 17112 1894 17252
rect 3087 17112 3133 17252
rect 4325 17112 4371 17252
rect 5564 17112 5610 17252
rect 754 16810 800 16856
rect 912 16810 958 16856
rect 1070 16810 1116 16856
rect 1228 16810 1274 16856
rect 1386 16810 1432 16856
rect 1544 16810 1590 16856
rect 1702 16810 1748 16856
rect 1993 16810 2039 16856
rect 2151 16810 2197 16856
rect 2309 16810 2355 16856
rect 2467 16810 2513 16856
rect 2625 16810 2671 16856
rect 2783 16810 2829 16856
rect 2941 16810 2987 16856
rect 3231 16810 3277 16856
rect 3389 16810 3435 16856
rect 3547 16810 3593 16856
rect 3705 16810 3751 16856
rect 3863 16810 3909 16856
rect 4021 16810 4067 16856
rect 4179 16810 4225 16856
rect 4470 16810 4516 16856
rect 4628 16810 4674 16856
rect 4786 16810 4832 16856
rect 4944 16810 4990 16856
rect 5102 16810 5148 16856
rect 5260 16810 5306 16856
rect 5418 16810 5464 16856
rect 2366 15463 2412 15509
rect 2366 15299 2412 15345
rect 2366 15136 2412 15182
rect 2366 14973 2412 15019
rect 2366 14810 2412 14856
rect 2366 14647 2412 14693
rect 2366 14483 2412 14529
rect 2366 14320 2412 14366
rect 2366 14157 2412 14203
rect 2366 13994 2412 14040
rect 2366 13830 2412 13876
rect 2366 13667 2412 13713
rect 2366 13504 2412 13550
rect 2366 13341 2412 13387
rect 2366 13177 2412 13223
rect 2366 13014 2412 13060
rect 2366 12851 2412 12897
rect 2366 12687 2412 12733
rect 2208 12525 2254 12571
rect 2366 12524 2412 12570
rect 2208 12361 2254 12407
rect 2366 12361 2412 12407
rect 2208 12198 2254 12244
rect 2366 12198 2412 12244
rect 2208 12035 2254 12081
rect 2366 12034 2412 12080
rect 2208 11872 2254 11918
rect 2366 11871 2412 11917
rect 2208 11708 2254 11754
rect 2366 11708 2412 11754
rect 2208 11545 2254 11591
rect 2366 11545 2412 11591
rect 2208 11382 2254 11428
rect 2366 11381 2412 11427
rect 2208 11218 2254 11264
rect 2366 11218 2412 11264
rect 2208 11055 2254 11101
rect 2366 11055 2412 11101
rect 2208 10892 2254 10938
rect 2366 10892 2412 10938
rect 2208 10729 2254 10775
rect 2366 10729 2412 10775
rect 2208 10565 2254 10611
rect 2366 10565 2412 10611
rect 300 9480 346 9526
rect 333 7991 379 8131
<< mvnsubdiffcont >>
rect 760 28879 806 28925
rect 918 28879 964 28925
rect 1076 28879 1122 28925
rect 1380 28879 1426 28925
rect 1538 28879 1584 28925
rect 1696 28879 1742 28925
rect 1999 28879 2045 28925
rect 2157 28879 2203 28925
rect 2315 28879 2361 28925
rect 2619 28879 2665 28925
rect 2777 28879 2823 28925
rect 2935 28879 2981 28925
rect 3237 28879 3283 28925
rect 3395 28879 3441 28925
rect 3553 28879 3599 28925
rect 3857 28879 3903 28925
rect 4015 28879 4061 28925
rect 4173 28879 4219 28925
rect 4476 28879 4522 28925
rect 4634 28879 4680 28925
rect 4792 28879 4838 28925
rect 5096 28879 5142 28925
rect 5254 28879 5300 28925
rect 5412 28879 5458 28925
rect 1228 24423 1274 24657
rect 2467 24423 2513 24657
rect 3705 24423 3751 24657
rect 4944 24423 4990 24657
rect 754 18129 800 18175
rect 912 18129 958 18175
rect 1070 18129 1116 18175
rect 1228 18129 1274 18175
rect 1386 18129 1432 18175
rect 1544 18129 1590 18175
rect 1702 18129 1748 18175
rect 1993 18129 2039 18175
rect 2151 18129 2197 18175
rect 2309 18129 2355 18175
rect 2467 18129 2513 18175
rect 2625 18129 2671 18175
rect 2783 18129 2829 18175
rect 2941 18129 2987 18175
rect 3231 18129 3277 18175
rect 3389 18129 3435 18175
rect 3547 18129 3593 18175
rect 3705 18129 3751 18175
rect 3863 18129 3909 18175
rect 4021 18129 4067 18175
rect 4179 18129 4225 18175
rect 4470 18129 4516 18175
rect 4628 18129 4674 18175
rect 4786 18129 4832 18175
rect 4944 18129 4990 18175
rect 5102 18129 5148 18175
rect 5260 18129 5306 18175
rect 5418 18129 5464 18175
rect 1665 15516 1899 15562
rect 300 8932 346 8978
rect 300 8768 346 8814
<< polysilicon >>
rect 769 28633 889 28706
rect 993 28633 1113 28706
rect 1389 28633 1509 28706
rect 1613 28633 1733 28706
rect 2008 28633 2128 28706
rect 2232 28633 2352 28706
rect 2628 28633 2748 28706
rect 2852 28633 2972 28706
rect 3246 28633 3366 28706
rect 3470 28633 3590 28706
rect 3866 28633 3986 28706
rect 4090 28633 4210 28706
rect 4485 28633 4605 28706
rect 4709 28633 4829 28706
rect 5069 28633 5189 28706
rect 5294 28633 5414 28706
rect 769 27858 889 27951
rect 993 27858 1113 27951
rect 1389 27858 1509 27951
rect 1613 27858 1733 27951
rect 2008 27858 2128 27951
rect 2232 27858 2352 27951
rect 2628 27858 2748 27951
rect 2852 27858 2972 27951
rect 3246 27858 3366 27951
rect 3470 27858 3590 27951
rect 3866 27858 3986 27951
rect 4090 27858 4210 27951
rect 4485 27858 4605 27951
rect 4709 27858 4829 27951
rect 5069 27858 5189 27951
rect 5294 27858 5414 27951
rect 769 27112 889 27176
rect 993 27112 1113 27176
rect 769 27093 1113 27112
rect 769 27047 847 27093
rect 1081 27047 1113 27093
rect 769 27028 1113 27047
rect 1389 27112 1509 27176
rect 1613 27112 1733 27176
rect 1389 27093 1733 27112
rect 1389 27047 1421 27093
rect 1655 27047 1733 27093
rect 1389 27028 1733 27047
rect 2008 27112 2128 27176
rect 2232 27112 2352 27176
rect 2008 27093 2352 27112
rect 2008 27047 2086 27093
rect 2320 27047 2352 27093
rect 2008 27028 2352 27047
rect 2628 27112 2748 27176
rect 2852 27112 2972 27176
rect 2628 27093 2972 27112
rect 2628 27047 2660 27093
rect 2894 27047 2972 27093
rect 2628 27028 2972 27047
rect 3246 27112 3366 27176
rect 3470 27112 3590 27176
rect 3246 27093 3590 27112
rect 3246 27047 3324 27093
rect 3558 27047 3590 27093
rect 3246 27028 3590 27047
rect 3866 27112 3986 27176
rect 4090 27112 4210 27176
rect 3866 27093 4210 27112
rect 3866 27047 3898 27093
rect 4132 27047 4210 27093
rect 3866 27028 4210 27047
rect 4485 27112 4605 27176
rect 4709 27112 4829 27176
rect 4485 27093 4829 27112
rect 4485 27047 4563 27093
rect 4797 27047 4829 27093
rect 4485 27028 4829 27047
rect 5069 27108 5189 27176
rect 5294 27108 5414 27176
rect 5069 27089 5414 27108
rect 5069 27043 5122 27089
rect 5356 27043 5414 27089
rect 883 26957 1003 27028
rect 1499 26957 1619 27028
rect 2122 26957 2242 27028
rect 2738 26957 2858 27028
rect 3360 26957 3480 27028
rect 3976 26957 4096 27028
rect 4599 26957 4719 27028
rect 5069 27024 5414 27043
rect 5215 26957 5335 27024
rect 883 25524 1003 25595
rect 1499 25524 1619 25595
rect 2122 25524 2242 25595
rect 2738 25524 2858 25595
rect 3360 25524 3480 25595
rect 3976 25524 4096 25595
rect 4599 25524 4719 25595
rect 5215 25524 5335 25595
rect 881 25370 1001 25444
rect 1501 25370 1621 25444
rect 2120 25370 2240 25444
rect 2740 25370 2860 25444
rect 3358 25370 3478 25444
rect 3978 25370 4098 25444
rect 4597 25370 4717 25444
rect 5217 25370 5337 25444
rect 881 23924 1001 24008
rect 881 23878 912 23924
rect 958 23878 1001 23924
rect 881 23859 1001 23878
rect 1501 23924 1621 24008
rect 1501 23878 1544 23924
rect 1590 23878 1621 23924
rect 1501 23859 1621 23878
rect 2120 23924 2240 24008
rect 2120 23878 2151 23924
rect 2197 23878 2240 23924
rect 2120 23859 2240 23878
rect 2740 23924 2860 24008
rect 2740 23878 2783 23924
rect 2829 23878 2860 23924
rect 2740 23859 2860 23878
rect 3358 23924 3478 24008
rect 3358 23878 3389 23924
rect 3435 23878 3478 23924
rect 3358 23859 3478 23878
rect 3978 23924 4098 24008
rect 3978 23878 4021 23924
rect 4067 23878 4098 23924
rect 3978 23859 4098 23878
rect 4597 23924 4717 24008
rect 4597 23878 4628 23924
rect 4674 23878 4717 23924
rect 4597 23859 4717 23878
rect 5217 23924 5337 24008
rect 5217 23878 5260 23924
rect 5306 23878 5337 23924
rect 5217 23859 5337 23878
rect 881 23679 1001 23753
rect 1501 23679 1621 23753
rect 2120 23679 2240 23753
rect 2740 23679 2860 23753
rect 3358 23679 3478 23753
rect 3978 23679 4098 23753
rect 4597 23679 4717 23753
rect 5217 23679 5337 23753
rect 881 22245 1001 22317
rect 882 21749 1001 22245
rect 1501 22245 1621 22317
rect 2120 22245 2240 22317
rect 881 21675 1001 21749
rect 1501 21749 1620 22245
rect 2121 21749 2240 22245
rect 2740 22245 2860 22317
rect 3358 22245 3478 22317
rect 1501 21675 1621 21749
rect 2120 21675 2240 21749
rect 2740 21749 2859 22245
rect 3359 21749 3478 22245
rect 3978 22245 4098 22317
rect 4597 22245 4717 22317
rect 2740 21675 2860 21749
rect 3358 21675 3478 21749
rect 3978 21749 4097 22245
rect 4598 21749 4717 22245
rect 3978 21675 4098 21749
rect 4597 21675 4717 21749
rect 5217 21675 5337 22317
rect 881 20229 1001 20313
rect 881 20183 918 20229
rect 964 20183 1001 20229
rect 881 20164 1001 20183
rect 1501 20229 1621 20313
rect 1501 20183 1538 20229
rect 1584 20183 1621 20229
rect 1501 20164 1621 20183
rect 2120 20229 2240 20313
rect 2120 20183 2157 20229
rect 2203 20183 2240 20229
rect 2120 20164 2240 20183
rect 2740 20229 2860 20313
rect 2740 20183 2777 20229
rect 2823 20183 2860 20229
rect 2740 20164 2860 20183
rect 3358 20229 3478 20313
rect 3358 20183 3395 20229
rect 3441 20183 3478 20229
rect 3358 20164 3478 20183
rect 3978 20229 4098 20313
rect 3978 20183 4015 20229
rect 4061 20183 4098 20229
rect 3978 20164 4098 20183
rect 4597 20229 4717 20313
rect 4597 20183 4634 20229
rect 4680 20183 4717 20229
rect 4597 20164 4717 20183
rect 5217 20229 5337 20313
rect 5217 20183 5254 20229
rect 5300 20183 5337 20229
rect 5217 20164 5337 20183
rect 881 19952 1001 19971
rect 881 19906 918 19952
rect 964 19906 1001 19952
rect 881 19820 1001 19906
rect 1501 19952 1621 19971
rect 1501 19906 1538 19952
rect 1584 19906 1621 19952
rect 1501 19820 1621 19906
rect 2120 19952 2240 19971
rect 2120 19906 2157 19952
rect 2203 19906 2240 19952
rect 2120 19820 2240 19906
rect 2740 19952 2860 19971
rect 2740 19906 2777 19952
rect 2823 19906 2860 19952
rect 2740 19820 2860 19906
rect 3358 19952 3478 19971
rect 3358 19906 3395 19952
rect 3441 19906 3478 19952
rect 3358 19820 3478 19906
rect 3978 19952 4098 19971
rect 3978 19906 4015 19952
rect 4061 19906 4098 19952
rect 3978 19820 4098 19906
rect 4597 19952 4717 19971
rect 4597 19906 4634 19952
rect 4680 19906 4717 19952
rect 4597 19820 4717 19906
rect 5217 19952 5337 19971
rect 5217 19906 5254 19952
rect 5300 19906 5337 19952
rect 5217 19820 5337 19906
rect 881 18387 1001 18458
rect 1501 18387 1621 18458
rect 2120 18387 2240 18458
rect 2740 18387 2860 18458
rect 3358 18387 3478 18458
rect 3978 18387 4098 18458
rect 4597 18387 4717 18458
rect 5217 18387 5337 18458
rect 812 17985 1184 18004
rect 812 17939 975 17985
rect 1021 17939 1184 17985
rect 812 17905 1184 17939
rect 812 17845 932 17905
rect 1064 17845 1184 17905
rect 1318 17985 1690 18004
rect 1318 17939 1481 17985
rect 1527 17939 1690 17985
rect 1318 17905 1690 17939
rect 1318 17845 1438 17905
rect 1570 17845 1690 17905
rect 2051 17985 2423 18004
rect 2051 17939 2214 17985
rect 2260 17939 2423 17985
rect 2051 17905 2423 17939
rect 2051 17845 2171 17905
rect 2303 17845 2423 17905
rect 2557 17985 2929 18004
rect 2557 17939 2720 17985
rect 2766 17939 2929 17985
rect 2557 17905 2929 17939
rect 2557 17845 2677 17905
rect 2809 17845 2929 17905
rect 3289 17985 3661 18004
rect 3289 17939 3452 17985
rect 3498 17939 3661 17985
rect 3289 17905 3661 17939
rect 3289 17845 3409 17905
rect 3541 17845 3661 17905
rect 3795 17985 4167 18004
rect 3795 17939 3958 17985
rect 4004 17939 4167 17985
rect 3795 17905 4167 17939
rect 3795 17845 3915 17905
rect 4047 17845 4167 17905
rect 4528 17985 4900 18004
rect 4528 17939 4691 17985
rect 4737 17939 4900 17985
rect 4528 17905 4900 17939
rect 4528 17845 4648 17905
rect 4780 17845 4900 17905
rect 5034 17985 5405 18004
rect 5034 17939 5197 17985
rect 5243 17939 5405 17985
rect 5034 17905 5405 17939
rect 5034 17845 5154 17905
rect 5285 17845 5405 17905
rect 812 17361 932 17548
rect 1064 17421 1184 17548
rect 855 17330 932 17361
rect 1079 17372 1184 17421
rect 1318 17421 1438 17548
rect 1318 17372 1423 17421
rect 855 17257 975 17330
rect 1079 17257 1199 17372
rect 1303 17257 1423 17372
rect 1570 17361 1690 17548
rect 2051 17361 2171 17548
rect 2303 17421 2423 17548
rect 1570 17330 1647 17361
rect 1527 17257 1647 17330
rect 2094 17330 2171 17361
rect 2318 17372 2423 17421
rect 2557 17421 2677 17548
rect 2557 17372 2662 17421
rect 2094 17257 2214 17330
rect 2318 17257 2438 17372
rect 2542 17257 2662 17372
rect 2809 17361 2929 17548
rect 3289 17361 3409 17548
rect 3541 17421 3661 17548
rect 2809 17330 2886 17361
rect 2766 17257 2886 17330
rect 3332 17330 3409 17361
rect 3556 17372 3661 17421
rect 3795 17421 3915 17548
rect 3795 17372 3900 17421
rect 855 17070 975 17143
rect 1079 17070 1199 17143
rect 1303 17070 1423 17143
rect 1527 17070 1647 17143
rect 3332 17257 3452 17330
rect 3556 17257 3676 17372
rect 3780 17257 3900 17372
rect 4047 17361 4167 17548
rect 4528 17361 4648 17548
rect 4780 17421 4900 17548
rect 4047 17330 4124 17361
rect 4004 17257 4124 17330
rect 4571 17330 4648 17361
rect 4795 17372 4900 17421
rect 5034 17395 5154 17548
rect 5285 17396 5405 17548
rect 2094 17070 2214 17143
rect 2318 17070 2438 17143
rect 2542 17070 2662 17143
rect 2766 17070 2886 17143
rect 4571 17257 4691 17330
rect 4795 17257 4915 17372
rect 5019 17358 5154 17395
rect 5243 17362 5405 17396
rect 5019 17257 5139 17358
rect 5243 17257 5363 17362
rect 3332 17070 3452 17143
rect 3556 17070 3676 17143
rect 3780 17070 3900 17143
rect 4004 17070 4124 17143
rect 4571 17070 4691 17143
rect 4795 17070 4915 17143
rect 5019 17070 5139 17143
rect 5243 17070 5363 17143
rect 375 15822 494 15850
rect 375 15778 495 15822
rect 1043 15704 1163 15777
rect 1043 15414 1163 15476
rect 916 15407 1163 15414
rect 916 15368 1321 15407
rect 916 15322 990 15368
rect 1036 15322 1321 15368
rect 1719 15324 1839 15368
rect 916 15277 1321 15322
rect 928 15267 1321 15277
rect 928 15197 1048 15267
rect 1201 15197 1321 15267
rect 928 14828 1048 14900
rect 1201 14828 1321 14900
rect 1034 14702 1228 14748
rect 1034 14656 1108 14702
rect 1154 14656 1228 14702
rect 1034 14538 1228 14656
rect 823 14478 1391 14538
rect 823 14418 943 14478
rect 1271 14418 1391 14478
rect 375 12620 495 13056
rect 823 12982 943 13056
rect 1271 12982 1391 13056
rect 1719 12905 1839 13056
rect 1574 12904 1839 12905
rect 1443 12859 1839 12904
rect 1443 12813 1516 12859
rect 1562 12813 1839 12859
rect 1443 12768 1839 12813
rect 1574 12767 1839 12768
rect 823 12619 943 12692
rect 1271 12619 1391 12692
rect 1719 12619 1839 12767
rect 823 10291 943 10351
rect 1271 10291 1391 10351
rect 823 10265 1391 10291
rect 1719 10278 1839 10351
rect 823 10219 976 10265
rect 1022 10219 1391 10265
rect 823 10200 1391 10219
rect 1704 10052 1824 10071
rect 1704 10006 1741 10052
rect 1787 10006 1824 10052
rect 1704 9911 1824 10006
rect 2556 9997 2676 10041
rect 375 9825 495 9898
rect 339 9780 531 9825
rect 986 9811 1106 9883
rect 339 9734 412 9780
rect 458 9734 531 9780
rect 339 9689 531 9734
rect 1704 9636 1824 9719
rect 986 9361 1106 9619
rect 1704 9576 2048 9636
rect 1704 9440 1824 9576
rect 1928 9440 2048 9576
rect 876 9307 1220 9361
rect 876 9247 996 9307
rect 1100 9247 1220 9307
rect 2556 9265 2676 9543
rect 1704 9140 1824 9212
rect 1928 9140 2048 9212
rect 1371 9027 1563 9072
rect 876 8932 996 9019
rect 1100 8947 1220 9019
rect 1371 8981 1444 9027
rect 1490 8996 1563 9027
rect 1490 8981 2048 8996
rect 1371 8936 2048 8981
rect 1927 8935 2048 8936
rect 802 8887 996 8932
rect 802 8841 875 8887
rect 921 8856 996 8887
rect 921 8841 1824 8856
rect 802 8796 1824 8841
rect 876 8795 1824 8796
rect 1704 8725 1824 8795
rect 1928 8725 2048 8935
rect 876 8643 996 8687
rect 1100 8643 1220 8687
rect 599 8341 793 8380
rect 876 8341 996 8451
rect 1100 8379 1220 8451
rect 1704 8380 1824 8533
rect 1928 8460 2048 8533
rect 599 8334 996 8341
rect 599 8288 673 8334
rect 719 8288 996 8334
rect 599 8281 996 8288
rect 599 8243 793 8281
rect 611 8242 793 8243
rect 876 8170 996 8281
rect 1044 8334 1236 8379
rect 1044 8288 1117 8334
rect 1163 8288 1236 8334
rect 1704 8319 2048 8380
rect 1044 8243 1236 8288
rect 1425 8269 1509 8278
rect 1425 8259 1824 8269
rect 1100 8170 1220 8243
rect 1425 8213 1444 8259
rect 1490 8213 1824 8259
rect 1425 8209 1824 8213
rect 1425 8194 1509 8209
rect 1704 8149 1824 8209
rect 1928 8149 2048 8319
rect 876 7934 996 7978
rect 1100 7934 1220 7978
rect 1704 7913 1824 7957
rect 1928 7913 2048 7957
rect 2556 7820 2676 7903
rect 2556 7774 2593 7820
rect 2639 7774 2676 7820
rect 2556 7755 2676 7774
<< polycontact >>
rect 847 27047 1081 27093
rect 1421 27047 1655 27093
rect 2086 27047 2320 27093
rect 2660 27047 2894 27093
rect 3324 27047 3558 27093
rect 3898 27047 4132 27093
rect 4563 27047 4797 27093
rect 5122 27043 5356 27089
rect 912 23878 958 23924
rect 1544 23878 1590 23924
rect 2151 23878 2197 23924
rect 2783 23878 2829 23924
rect 3389 23878 3435 23924
rect 4021 23878 4067 23924
rect 4628 23878 4674 23924
rect 5260 23878 5306 23924
rect 918 20183 964 20229
rect 1538 20183 1584 20229
rect 2157 20183 2203 20229
rect 2777 20183 2823 20229
rect 3395 20183 3441 20229
rect 4015 20183 4061 20229
rect 4634 20183 4680 20229
rect 5254 20183 5300 20229
rect 918 19906 964 19952
rect 1538 19906 1584 19952
rect 2157 19906 2203 19952
rect 2777 19906 2823 19952
rect 3395 19906 3441 19952
rect 4015 19906 4061 19952
rect 4634 19906 4680 19952
rect 5254 19906 5300 19952
rect 975 17939 1021 17985
rect 1481 17939 1527 17985
rect 2214 17939 2260 17985
rect 2720 17939 2766 17985
rect 3452 17939 3498 17985
rect 3958 17939 4004 17985
rect 4691 17939 4737 17985
rect 5197 17939 5243 17985
rect 990 15322 1036 15368
rect 1108 14656 1154 14702
rect 1516 12813 1562 12859
rect 976 10219 1022 10265
rect 1741 10006 1787 10052
rect 412 9734 458 9780
rect 1444 8981 1490 9027
rect 875 8841 921 8887
rect 673 8288 719 8334
rect 1117 8288 1163 8334
rect 1444 8213 1490 8259
rect 2593 7774 2639 7820
<< metal1 >>
rect 631 28963 5587 28987
rect 631 28925 918 28963
rect 970 28925 1532 28963
rect 1584 28925 2157 28963
rect 2209 28925 2771 28963
rect 2823 28925 3395 28963
rect 3447 28925 4009 28963
rect 4061 28925 4634 28963
rect 4686 28925 5248 28963
rect 5300 28925 5587 28963
rect 631 28879 760 28925
rect 806 28879 918 28925
rect 970 28911 1076 28925
rect 964 28879 1076 28911
rect 1122 28879 1380 28925
rect 1426 28911 1532 28925
rect 1426 28879 1538 28911
rect 1584 28879 1696 28925
rect 1742 28879 1999 28925
rect 2045 28879 2157 28925
rect 2209 28911 2315 28925
rect 2203 28879 2315 28911
rect 2361 28879 2619 28925
rect 2665 28911 2771 28925
rect 2665 28879 2777 28911
rect 2823 28879 2935 28925
rect 2981 28879 3237 28925
rect 3283 28879 3395 28925
rect 3447 28911 3553 28925
rect 3441 28879 3553 28911
rect 3599 28879 3857 28925
rect 3903 28911 4009 28925
rect 3903 28879 4015 28911
rect 4061 28879 4173 28925
rect 4219 28879 4476 28925
rect 4522 28879 4634 28925
rect 4686 28911 4792 28925
rect 4680 28879 4792 28911
rect 4838 28879 5096 28925
rect 5142 28911 5248 28925
rect 5142 28879 5254 28911
rect 5300 28879 5412 28925
rect 5458 28879 5587 28925
rect 631 28777 5587 28879
rect 631 28725 918 28777
rect 970 28725 1532 28777
rect 1584 28725 2157 28777
rect 2209 28725 2771 28777
rect 2823 28725 3395 28777
rect 3447 28725 4009 28777
rect 4061 28725 4634 28777
rect 4686 28725 5248 28777
rect 5300 28725 5587 28777
rect 631 28704 5587 28725
rect 631 28588 779 28704
rect 631 28542 692 28588
rect 738 28542 779 28588
rect 631 28406 779 28542
rect 631 28360 692 28406
rect 738 28360 779 28406
rect 631 28225 779 28360
rect 631 28179 692 28225
rect 738 28179 779 28225
rect 631 28043 779 28179
rect 631 27997 692 28043
rect 738 27997 779 28043
rect 631 27812 779 27997
rect 884 28588 999 28624
rect 884 28542 918 28588
rect 964 28542 999 28588
rect 884 28406 999 28542
rect 884 28393 918 28406
rect 964 28393 999 28406
rect 884 28237 914 28393
rect 966 28237 999 28393
rect 884 28225 999 28237
rect 884 28179 918 28225
rect 964 28179 999 28225
rect 884 28043 999 28179
rect 884 27997 918 28043
rect 964 27997 999 28043
rect 884 27960 999 27997
rect 1104 28588 1398 28704
rect 1104 28542 1228 28588
rect 1274 28542 1398 28588
rect 1104 28406 1398 28542
rect 1104 28360 1228 28406
rect 1274 28360 1398 28406
rect 1104 28225 1398 28360
rect 1104 28179 1228 28225
rect 1274 28179 1398 28225
rect 1104 28043 1398 28179
rect 1104 27997 1228 28043
rect 1274 27997 1398 28043
rect 631 27766 692 27812
rect 738 27766 779 27812
rect 631 27631 779 27766
rect 631 27585 692 27631
rect 738 27585 779 27631
rect 631 27450 779 27585
rect 631 27404 692 27450
rect 738 27404 779 27450
rect 631 27268 779 27404
rect 631 27222 692 27268
rect 738 27222 779 27268
rect 631 27185 779 27222
rect 884 27812 999 27849
rect 884 27766 918 27812
rect 964 27766 999 27812
rect 884 27631 999 27766
rect 884 27618 918 27631
rect 964 27618 999 27631
rect 884 27462 914 27618
rect 966 27462 999 27618
rect 884 27450 999 27462
rect 884 27404 918 27450
rect 964 27404 999 27450
rect 884 27268 999 27404
rect 884 27222 918 27268
rect 964 27222 999 27268
rect 884 27185 999 27222
rect 1104 27812 1398 27997
rect 1503 28588 1618 28624
rect 1503 28542 1538 28588
rect 1584 28542 1618 28588
rect 1503 28406 1618 28542
rect 1503 28393 1538 28406
rect 1584 28393 1618 28406
rect 1503 28237 1536 28393
rect 1588 28237 1618 28393
rect 1503 28225 1618 28237
rect 1503 28179 1538 28225
rect 1584 28179 1618 28225
rect 1503 28043 1618 28179
rect 1503 27997 1538 28043
rect 1584 27997 1618 28043
rect 1503 27960 1618 27997
rect 1723 28588 2018 28704
rect 1723 28542 1764 28588
rect 1810 28542 1931 28588
rect 1977 28542 2018 28588
rect 1723 28406 2018 28542
rect 1723 28360 1764 28406
rect 1810 28360 1931 28406
rect 1977 28360 2018 28406
rect 1723 28225 2018 28360
rect 1723 28179 1764 28225
rect 1810 28179 1931 28225
rect 1977 28179 2018 28225
rect 1723 28043 2018 28179
rect 1723 27997 1764 28043
rect 1810 27997 1931 28043
rect 1977 27997 2018 28043
rect 1104 27766 1228 27812
rect 1274 27766 1398 27812
rect 1104 27631 1398 27766
rect 1104 27585 1228 27631
rect 1274 27585 1398 27631
rect 1104 27450 1398 27585
rect 1104 27404 1228 27450
rect 1274 27404 1398 27450
rect 1104 27268 1398 27404
rect 1104 27222 1228 27268
rect 1274 27222 1398 27268
rect 1104 27185 1398 27222
rect 1503 27812 1618 27849
rect 1503 27766 1538 27812
rect 1584 27766 1618 27812
rect 1503 27631 1618 27766
rect 1503 27618 1538 27631
rect 1584 27618 1618 27631
rect 1503 27462 1536 27618
rect 1588 27462 1618 27618
rect 1503 27450 1618 27462
rect 1503 27404 1538 27450
rect 1584 27404 1618 27450
rect 1503 27268 1618 27404
rect 1503 27222 1538 27268
rect 1584 27222 1618 27268
rect 1503 27185 1618 27222
rect 1723 27812 2018 27997
rect 2123 28588 2238 28624
rect 2123 28542 2157 28588
rect 2203 28542 2238 28588
rect 2123 28406 2238 28542
rect 2123 28393 2157 28406
rect 2203 28393 2238 28406
rect 2123 28237 2153 28393
rect 2205 28237 2238 28393
rect 2123 28225 2238 28237
rect 2123 28179 2157 28225
rect 2203 28179 2238 28225
rect 2123 28043 2238 28179
rect 2123 27997 2157 28043
rect 2203 27997 2238 28043
rect 2123 27960 2238 27997
rect 2343 28588 2637 28704
rect 2343 28542 2467 28588
rect 2513 28542 2637 28588
rect 2343 28406 2637 28542
rect 2343 28360 2467 28406
rect 2513 28360 2637 28406
rect 2343 28225 2637 28360
rect 2343 28179 2467 28225
rect 2513 28179 2637 28225
rect 2343 28043 2637 28179
rect 2343 27997 2467 28043
rect 2513 27997 2637 28043
rect 1723 27766 1764 27812
rect 1810 27766 1931 27812
rect 1977 27766 2018 27812
rect 1723 27631 2018 27766
rect 1723 27585 1764 27631
rect 1810 27585 1931 27631
rect 1977 27585 2018 27631
rect 1723 27450 2018 27585
rect 1723 27404 1764 27450
rect 1810 27404 1931 27450
rect 1977 27404 2018 27450
rect 1723 27268 2018 27404
rect 1723 27222 1764 27268
rect 1810 27222 1931 27268
rect 1977 27222 2018 27268
rect 1723 27185 2018 27222
rect 2123 27812 2238 27849
rect 2123 27766 2157 27812
rect 2203 27766 2238 27812
rect 2123 27631 2238 27766
rect 2123 27618 2157 27631
rect 2203 27618 2238 27631
rect 2123 27462 2153 27618
rect 2205 27462 2238 27618
rect 2123 27450 2238 27462
rect 2123 27404 2157 27450
rect 2203 27404 2238 27450
rect 2123 27268 2238 27404
rect 2123 27222 2157 27268
rect 2203 27222 2238 27268
rect 2123 27185 2238 27222
rect 2343 27812 2637 27997
rect 2742 28588 2857 28624
rect 2742 28542 2777 28588
rect 2823 28542 2857 28588
rect 2742 28406 2857 28542
rect 2742 28393 2777 28406
rect 2823 28393 2857 28406
rect 2742 28237 2775 28393
rect 2827 28237 2857 28393
rect 2742 28225 2857 28237
rect 2742 28179 2777 28225
rect 2823 28179 2857 28225
rect 2742 28043 2857 28179
rect 2742 27997 2777 28043
rect 2823 27997 2857 28043
rect 2742 27960 2857 27997
rect 2962 28588 3256 28704
rect 2962 28542 3003 28588
rect 3049 28542 3169 28588
rect 3215 28542 3256 28588
rect 2962 28406 3256 28542
rect 2962 28360 3003 28406
rect 3049 28360 3169 28406
rect 3215 28360 3256 28406
rect 2962 28225 3256 28360
rect 2962 28179 3003 28225
rect 3049 28179 3169 28225
rect 3215 28179 3256 28225
rect 2962 28043 3256 28179
rect 2962 27997 3003 28043
rect 3049 27997 3169 28043
rect 3215 27997 3256 28043
rect 2343 27766 2467 27812
rect 2513 27766 2637 27812
rect 2343 27631 2637 27766
rect 2343 27585 2467 27631
rect 2513 27585 2637 27631
rect 2343 27450 2637 27585
rect 2343 27404 2467 27450
rect 2513 27404 2637 27450
rect 2343 27268 2637 27404
rect 2343 27222 2467 27268
rect 2513 27222 2637 27268
rect 2343 27185 2637 27222
rect 2742 27812 2857 27849
rect 2742 27766 2777 27812
rect 2823 27766 2857 27812
rect 2742 27631 2857 27766
rect 2742 27618 2777 27631
rect 2823 27618 2857 27631
rect 2742 27462 2775 27618
rect 2827 27462 2857 27618
rect 2742 27450 2857 27462
rect 2742 27404 2777 27450
rect 2823 27404 2857 27450
rect 2742 27268 2857 27404
rect 2742 27222 2777 27268
rect 2823 27222 2857 27268
rect 2742 27185 2857 27222
rect 2962 27812 3256 27997
rect 3361 28588 3476 28624
rect 3361 28542 3395 28588
rect 3441 28542 3476 28588
rect 3361 28406 3476 28542
rect 3361 28393 3395 28406
rect 3441 28393 3476 28406
rect 3361 28237 3391 28393
rect 3443 28237 3476 28393
rect 3361 28225 3476 28237
rect 3361 28179 3395 28225
rect 3441 28179 3476 28225
rect 3361 28043 3476 28179
rect 3361 27997 3395 28043
rect 3441 27997 3476 28043
rect 3361 27960 3476 27997
rect 3581 28588 3875 28704
rect 3581 28542 3705 28588
rect 3751 28542 3875 28588
rect 3581 28406 3875 28542
rect 3581 28360 3705 28406
rect 3751 28360 3875 28406
rect 3581 28225 3875 28360
rect 3581 28179 3705 28225
rect 3751 28179 3875 28225
rect 3581 28043 3875 28179
rect 3581 27997 3705 28043
rect 3751 27997 3875 28043
rect 2962 27766 3003 27812
rect 3049 27766 3169 27812
rect 3215 27766 3256 27812
rect 2962 27631 3256 27766
rect 2962 27585 3003 27631
rect 3049 27585 3169 27631
rect 3215 27585 3256 27631
rect 2962 27450 3256 27585
rect 2962 27404 3003 27450
rect 3049 27404 3169 27450
rect 3215 27404 3256 27450
rect 2962 27268 3256 27404
rect 2962 27222 3003 27268
rect 3049 27222 3169 27268
rect 3215 27222 3256 27268
rect 2962 27185 3256 27222
rect 3361 27812 3476 27849
rect 3361 27766 3395 27812
rect 3441 27766 3476 27812
rect 3361 27631 3476 27766
rect 3361 27618 3395 27631
rect 3441 27618 3476 27631
rect 3361 27462 3391 27618
rect 3443 27462 3476 27618
rect 3361 27450 3476 27462
rect 3361 27404 3395 27450
rect 3441 27404 3476 27450
rect 3361 27268 3476 27404
rect 3361 27222 3395 27268
rect 3441 27222 3476 27268
rect 3361 27185 3476 27222
rect 3581 27812 3875 27997
rect 3980 28588 4095 28624
rect 3980 28542 4015 28588
rect 4061 28542 4095 28588
rect 3980 28406 4095 28542
rect 3980 28393 4015 28406
rect 4061 28393 4095 28406
rect 3980 28237 4013 28393
rect 4065 28237 4095 28393
rect 3980 28225 4095 28237
rect 3980 28179 4015 28225
rect 4061 28179 4095 28225
rect 3980 28043 4095 28179
rect 3980 27997 4015 28043
rect 4061 27997 4095 28043
rect 3980 27960 4095 27997
rect 4200 28588 4495 28704
rect 4200 28542 4241 28588
rect 4287 28542 4408 28588
rect 4454 28542 4495 28588
rect 4200 28406 4495 28542
rect 4200 28360 4241 28406
rect 4287 28360 4408 28406
rect 4454 28360 4495 28406
rect 4200 28225 4495 28360
rect 4200 28179 4241 28225
rect 4287 28179 4408 28225
rect 4454 28179 4495 28225
rect 4200 28043 4495 28179
rect 4200 27997 4241 28043
rect 4287 27997 4408 28043
rect 4454 27997 4495 28043
rect 3581 27766 3705 27812
rect 3751 27766 3875 27812
rect 3581 27631 3875 27766
rect 3581 27585 3705 27631
rect 3751 27585 3875 27631
rect 3581 27450 3875 27585
rect 3581 27404 3705 27450
rect 3751 27404 3875 27450
rect 3581 27268 3875 27404
rect 3581 27222 3705 27268
rect 3751 27222 3875 27268
rect 3581 27185 3875 27222
rect 3980 27812 4095 27849
rect 3980 27766 4015 27812
rect 4061 27766 4095 27812
rect 3980 27631 4095 27766
rect 3980 27618 4015 27631
rect 4061 27618 4095 27631
rect 3980 27462 4013 27618
rect 4065 27462 4095 27618
rect 3980 27450 4095 27462
rect 3980 27404 4015 27450
rect 4061 27404 4095 27450
rect 3980 27268 4095 27404
rect 3980 27222 4015 27268
rect 4061 27222 4095 27268
rect 3980 27185 4095 27222
rect 4200 27812 4495 27997
rect 4600 28588 4715 28624
rect 4600 28542 4634 28588
rect 4680 28542 4715 28588
rect 4600 28406 4715 28542
rect 4600 28393 4634 28406
rect 4680 28393 4715 28406
rect 4600 28237 4630 28393
rect 4682 28237 4715 28393
rect 4600 28225 4715 28237
rect 4600 28179 4634 28225
rect 4680 28179 4715 28225
rect 4600 28043 4715 28179
rect 4600 27997 4634 28043
rect 4680 27997 4715 28043
rect 4600 27960 4715 27997
rect 4820 28588 5025 28704
rect 4820 28542 4944 28588
rect 4990 28542 5025 28588
rect 4820 28406 5025 28542
rect 4820 28360 4944 28406
rect 4990 28360 5025 28406
rect 4820 28225 5025 28360
rect 4820 28179 4944 28225
rect 4990 28179 5025 28225
rect 4820 28043 5025 28179
rect 4820 27997 4944 28043
rect 4990 27997 5025 28043
rect 4200 27766 4241 27812
rect 4287 27766 4408 27812
rect 4454 27766 4495 27812
rect 4200 27631 4495 27766
rect 4200 27585 4241 27631
rect 4287 27585 4408 27631
rect 4454 27585 4495 27631
rect 4200 27450 4495 27585
rect 4200 27404 4241 27450
rect 4287 27404 4408 27450
rect 4454 27404 4495 27450
rect 4200 27268 4495 27404
rect 4200 27222 4241 27268
rect 4287 27222 4408 27268
rect 4454 27222 4495 27268
rect 4200 27185 4495 27222
rect 4600 27812 4715 27849
rect 4600 27766 4634 27812
rect 4680 27766 4715 27812
rect 4600 27631 4715 27766
rect 4600 27618 4634 27631
rect 4680 27618 4715 27631
rect 4600 27462 4630 27618
rect 4682 27462 4715 27618
rect 4600 27450 4715 27462
rect 4600 27404 4634 27450
rect 4680 27404 4715 27450
rect 4600 27268 4715 27404
rect 4600 27222 4634 27268
rect 4680 27222 4715 27268
rect 4600 27185 4715 27222
rect 4820 27812 5025 27997
rect 5184 28588 5300 28624
rect 5184 28542 5219 28588
rect 5265 28542 5300 28588
rect 5184 28406 5300 28542
rect 5184 28360 5219 28406
rect 5265 28393 5300 28406
rect 5184 28341 5226 28360
rect 5278 28341 5300 28393
rect 5184 28225 5300 28341
rect 5184 28179 5219 28225
rect 5265 28207 5300 28225
rect 5184 28155 5226 28179
rect 5278 28155 5300 28207
rect 5184 28043 5300 28155
rect 5184 27997 5219 28043
rect 5265 27997 5300 28043
rect 5184 27960 5300 27997
rect 5445 28588 5587 28704
rect 5445 28542 5480 28588
rect 5526 28542 5587 28588
rect 5445 28406 5587 28542
rect 5445 28360 5480 28406
rect 5526 28360 5587 28406
rect 5445 28225 5587 28360
rect 5445 28179 5480 28225
rect 5526 28179 5587 28225
rect 5445 28043 5587 28179
rect 5445 27997 5480 28043
rect 5526 27997 5587 28043
rect 4820 27766 4944 27812
rect 4990 27766 5025 27812
rect 4820 27631 5025 27766
rect 4820 27585 4944 27631
rect 4990 27585 5025 27631
rect 4820 27450 5025 27585
rect 4820 27404 4944 27450
rect 4990 27404 5025 27450
rect 4820 27268 5025 27404
rect 4820 27222 4944 27268
rect 4990 27222 5025 27268
rect 4820 27185 5025 27222
rect 5184 27812 5300 27849
rect 5184 27766 5219 27812
rect 5265 27766 5300 27812
rect 5184 27631 5300 27766
rect 5184 27618 5219 27631
rect 5265 27618 5300 27631
rect 5184 27462 5216 27618
rect 5268 27462 5300 27618
rect 5184 27450 5300 27462
rect 5184 27404 5219 27450
rect 5265 27404 5300 27450
rect 5184 27268 5300 27404
rect 5184 27222 5219 27268
rect 5265 27222 5300 27268
rect 5184 27185 5300 27222
rect 5445 27812 5587 27997
rect 5445 27766 5480 27812
rect 5526 27766 5587 27812
rect 5445 27631 5587 27766
rect 5445 27585 5480 27631
rect 5526 27585 5587 27631
rect 5445 27450 5587 27585
rect 5445 27404 5480 27450
rect 5526 27404 5587 27450
rect 5445 27268 5587 27404
rect 5445 27222 5480 27268
rect 5526 27222 5587 27268
rect 5445 27185 5587 27222
rect 487 27093 5519 27105
rect 487 27041 499 27093
rect 551 27047 847 27093
rect 1081 27047 1421 27093
rect 1655 27047 2086 27093
rect 2320 27047 2660 27093
rect 2894 27047 3324 27093
rect 3558 27047 3898 27093
rect 4132 27047 4563 27093
rect 4797 27089 5519 27093
rect 4797 27047 5122 27089
rect 551 27043 5122 27047
rect 5356 27043 5519 27089
rect 551 27041 5519 27043
rect 487 27031 5519 27041
rect 487 27029 563 27031
rect 808 26944 854 26957
rect 808 26836 854 26898
rect 808 26728 854 26790
rect 808 26620 854 26682
rect 808 26512 854 26574
rect 808 26410 854 26466
rect 687 26404 854 26410
rect 687 26398 808 26404
rect 687 26242 699 26398
rect 751 26358 808 26398
rect 751 26296 854 26358
rect 751 26250 808 26296
rect 751 26242 854 26250
rect 687 26230 854 26242
rect 808 26189 854 26230
rect 808 26082 854 26143
rect 808 25975 854 26036
rect 808 25868 854 25929
rect 808 25761 854 25822
rect 808 25654 854 25715
rect 808 25595 854 25608
rect 1032 26944 1078 26957
rect 1032 26836 1078 26898
rect 1032 26728 1078 26790
rect 1032 26620 1078 26682
rect 1032 26512 1078 26574
rect 1032 26410 1078 26466
rect 1424 26944 1470 26957
rect 1424 26836 1470 26898
rect 1424 26728 1470 26790
rect 1424 26620 1470 26682
rect 1424 26512 1470 26574
rect 1424 26410 1470 26466
rect 1032 26404 1193 26410
rect 1078 26398 1193 26404
rect 1078 26358 1129 26398
rect 1032 26296 1129 26358
rect 1078 26250 1129 26296
rect 1032 26242 1129 26250
rect 1181 26242 1193 26398
rect 1032 26230 1193 26242
rect 1309 26404 1470 26410
rect 1309 26398 1424 26404
rect 1309 26242 1321 26398
rect 1373 26358 1424 26398
rect 1373 26296 1470 26358
rect 1373 26250 1424 26296
rect 1373 26242 1470 26250
rect 1309 26230 1470 26242
rect 1032 26189 1078 26230
rect 1032 26082 1078 26143
rect 1032 25975 1078 26036
rect 1032 25868 1078 25929
rect 1032 25761 1078 25822
rect 1032 25654 1078 25715
rect 1032 25595 1078 25608
rect 1424 26189 1470 26230
rect 1424 26082 1470 26143
rect 1424 25975 1470 26036
rect 1424 25868 1470 25929
rect 1424 25761 1470 25822
rect 1424 25654 1470 25715
rect 1424 25595 1470 25608
rect 1648 26944 1694 26957
rect 1648 26836 1694 26898
rect 1648 26728 1694 26790
rect 1648 26620 1694 26682
rect 1648 26512 1694 26574
rect 1648 26410 1694 26466
rect 2047 26944 2093 26957
rect 2047 26836 2093 26898
rect 2047 26728 2093 26790
rect 2047 26620 2093 26682
rect 2047 26512 2093 26574
rect 2047 26410 2093 26466
rect 1648 26404 1815 26410
rect 1694 26398 1815 26404
rect 1694 26358 1751 26398
rect 1648 26296 1751 26358
rect 1694 26250 1751 26296
rect 1648 26242 1751 26250
rect 1803 26242 1815 26398
rect 1648 26230 1815 26242
rect 1926 26404 2093 26410
rect 1926 26398 2047 26404
rect 1926 26242 1938 26398
rect 1990 26358 2047 26398
rect 1990 26296 2093 26358
rect 1990 26250 2047 26296
rect 1990 26242 2093 26250
rect 1926 26230 2093 26242
rect 1648 26189 1694 26230
rect 1648 26082 1694 26143
rect 1648 25975 1694 26036
rect 1648 25868 1694 25929
rect 1648 25761 1694 25822
rect 1648 25654 1694 25715
rect 1648 25595 1694 25608
rect 2047 26189 2093 26230
rect 2047 26082 2093 26143
rect 2047 25975 2093 26036
rect 2047 25868 2093 25929
rect 2047 25761 2093 25822
rect 2047 25654 2093 25715
rect 2047 25595 2093 25608
rect 2271 26944 2317 26957
rect 2271 26836 2317 26898
rect 2271 26728 2317 26790
rect 2271 26620 2317 26682
rect 2271 26512 2317 26574
rect 2271 26410 2317 26466
rect 2663 26944 2709 26957
rect 2663 26836 2709 26898
rect 2663 26728 2709 26790
rect 2663 26620 2709 26682
rect 2663 26512 2709 26574
rect 2663 26410 2709 26466
rect 2271 26404 2432 26410
rect 2317 26398 2432 26404
rect 2317 26358 2368 26398
rect 2271 26296 2368 26358
rect 2317 26250 2368 26296
rect 2271 26242 2368 26250
rect 2420 26242 2432 26398
rect 2271 26230 2432 26242
rect 2548 26404 2709 26410
rect 2548 26398 2663 26404
rect 2548 26242 2560 26398
rect 2612 26358 2663 26398
rect 2612 26296 2709 26358
rect 2612 26250 2663 26296
rect 2612 26242 2709 26250
rect 2548 26230 2709 26242
rect 2271 26189 2317 26230
rect 2271 26082 2317 26143
rect 2271 25975 2317 26036
rect 2271 25868 2317 25929
rect 2271 25761 2317 25822
rect 2271 25654 2317 25715
rect 2271 25595 2317 25608
rect 2663 26189 2709 26230
rect 2663 26082 2709 26143
rect 2663 25975 2709 26036
rect 2663 25868 2709 25929
rect 2663 25761 2709 25822
rect 2663 25654 2709 25715
rect 2663 25595 2709 25608
rect 2887 26944 2933 26957
rect 2887 26836 2933 26898
rect 2887 26728 2933 26790
rect 2887 26620 2933 26682
rect 2887 26512 2933 26574
rect 2887 26410 2933 26466
rect 3285 26944 3331 26957
rect 3285 26836 3331 26898
rect 3285 26728 3331 26790
rect 3285 26620 3331 26682
rect 3285 26512 3331 26574
rect 3285 26410 3331 26466
rect 2887 26404 3054 26410
rect 2933 26398 3054 26404
rect 2933 26358 2990 26398
rect 2887 26296 2990 26358
rect 2933 26250 2990 26296
rect 2887 26242 2990 26250
rect 3042 26242 3054 26398
rect 2887 26230 3054 26242
rect 3164 26404 3331 26410
rect 3164 26398 3285 26404
rect 3164 26242 3176 26398
rect 3228 26358 3285 26398
rect 3228 26296 3331 26358
rect 3228 26250 3285 26296
rect 3228 26242 3331 26250
rect 3164 26230 3331 26242
rect 2887 26189 2933 26230
rect 2887 26082 2933 26143
rect 2887 25975 2933 26036
rect 2887 25868 2933 25929
rect 2887 25761 2933 25822
rect 2887 25654 2933 25715
rect 2887 25595 2933 25608
rect 3285 26189 3331 26230
rect 3285 26082 3331 26143
rect 3285 25975 3331 26036
rect 3285 25868 3331 25929
rect 3285 25761 3331 25822
rect 3285 25654 3331 25715
rect 3285 25595 3331 25608
rect 3509 26944 3555 26957
rect 3509 26836 3555 26898
rect 3509 26728 3555 26790
rect 3509 26620 3555 26682
rect 3509 26512 3555 26574
rect 3509 26410 3555 26466
rect 3901 26944 3947 26957
rect 3901 26836 3947 26898
rect 3901 26728 3947 26790
rect 3901 26620 3947 26682
rect 3901 26512 3947 26574
rect 3901 26410 3947 26466
rect 3509 26404 3670 26410
rect 3555 26398 3670 26404
rect 3555 26358 3606 26398
rect 3509 26296 3606 26358
rect 3555 26250 3606 26296
rect 3509 26242 3606 26250
rect 3658 26242 3670 26398
rect 3509 26230 3670 26242
rect 3786 26404 3947 26410
rect 3786 26398 3901 26404
rect 3786 26242 3798 26398
rect 3850 26358 3901 26398
rect 3850 26296 3947 26358
rect 3850 26250 3901 26296
rect 3850 26242 3947 26250
rect 3786 26230 3947 26242
rect 3509 26189 3555 26230
rect 3509 26082 3555 26143
rect 3509 25975 3555 26036
rect 3509 25868 3555 25929
rect 3509 25761 3555 25822
rect 3509 25654 3555 25715
rect 3509 25595 3555 25608
rect 3901 26189 3947 26230
rect 3901 26082 3947 26143
rect 3901 25975 3947 26036
rect 3901 25868 3947 25929
rect 3901 25761 3947 25822
rect 3901 25654 3947 25715
rect 3901 25595 3947 25608
rect 4125 26944 4171 26957
rect 4125 26836 4171 26898
rect 4125 26728 4171 26790
rect 4125 26620 4171 26682
rect 4125 26512 4171 26574
rect 4125 26410 4171 26466
rect 4524 26944 4570 26957
rect 4524 26836 4570 26898
rect 4524 26728 4570 26790
rect 4524 26620 4570 26682
rect 4524 26512 4570 26574
rect 4524 26410 4570 26466
rect 4125 26404 4292 26410
rect 4171 26398 4292 26404
rect 4171 26358 4228 26398
rect 4125 26296 4228 26358
rect 4171 26250 4228 26296
rect 4125 26242 4228 26250
rect 4280 26242 4292 26398
rect 4125 26230 4292 26242
rect 4403 26404 4570 26410
rect 4403 26398 4524 26404
rect 4403 26242 4415 26398
rect 4467 26358 4524 26398
rect 4467 26296 4570 26358
rect 4467 26250 4524 26296
rect 4467 26242 4570 26250
rect 4403 26230 4570 26242
rect 4125 26189 4171 26230
rect 4125 26082 4171 26143
rect 4125 25975 4171 26036
rect 4125 25868 4171 25929
rect 4125 25761 4171 25822
rect 4125 25654 4171 25715
rect 4125 25595 4171 25608
rect 4524 26189 4570 26230
rect 4524 26082 4570 26143
rect 4524 25975 4570 26036
rect 4524 25868 4570 25929
rect 4524 25761 4570 25822
rect 4524 25654 4570 25715
rect 4524 25595 4570 25608
rect 4748 26944 4794 26957
rect 4748 26836 4794 26898
rect 4748 26728 4794 26790
rect 4748 26620 4794 26682
rect 4748 26512 4794 26574
rect 4748 26410 4794 26466
rect 5140 26944 5186 26957
rect 5140 26836 5186 26898
rect 5140 26728 5186 26790
rect 5140 26620 5186 26682
rect 5140 26512 5186 26574
rect 5140 26410 5186 26466
rect 4748 26404 4909 26410
rect 4794 26398 4909 26404
rect 4794 26358 4845 26398
rect 4748 26296 4845 26358
rect 4794 26250 4845 26296
rect 4748 26242 4845 26250
rect 4897 26242 4909 26398
rect 4748 26230 4909 26242
rect 5029 26404 5186 26410
rect 5029 26398 5140 26404
rect 5029 26242 5041 26398
rect 5093 26358 5140 26398
rect 5093 26296 5186 26358
rect 5093 26250 5140 26296
rect 5093 26242 5186 26250
rect 5029 26230 5186 26242
rect 4748 26189 4794 26230
rect 4748 26082 4794 26143
rect 4748 25975 4794 26036
rect 4748 25868 4794 25929
rect 4748 25761 4794 25822
rect 4748 25654 4794 25715
rect 4748 25595 4794 25608
rect 5140 26189 5186 26230
rect 5140 26082 5186 26143
rect 5140 25975 5186 26036
rect 5140 25868 5186 25929
rect 5140 25761 5186 25822
rect 5140 25654 5186 25715
rect 5140 25595 5186 25608
rect 5364 26944 5410 26957
rect 5364 26836 5410 26898
rect 5364 26728 5410 26790
rect 5364 26620 5410 26682
rect 5364 26512 5410 26574
rect 5364 26410 5410 26466
rect 5364 26404 5523 26410
rect 5410 26398 5523 26404
rect 5410 26358 5459 26398
rect 5364 26296 5459 26358
rect 5410 26250 5459 26296
rect 5364 26242 5459 26250
rect 5511 26242 5523 26398
rect 5364 26230 5523 26242
rect 5364 26189 5410 26230
rect 5364 26082 5410 26143
rect 5364 25975 5410 26036
rect 5364 25868 5410 25929
rect 5364 25761 5410 25822
rect 5364 25654 5410 25715
rect 5364 25595 5410 25608
rect 702 25357 852 25370
rect 702 25311 806 25357
rect 702 25249 852 25311
rect 702 25203 806 25249
rect 702 25141 852 25203
rect 702 25095 806 25141
rect 702 25033 852 25095
rect 702 24987 806 25033
rect 702 24925 852 24987
rect 702 24879 806 24925
rect 702 24817 852 24879
rect 702 24771 806 24817
rect 702 24709 852 24771
rect 702 24663 806 24709
rect 702 24602 852 24663
rect 702 24556 806 24602
rect 702 24495 852 24556
rect 702 24449 806 24495
rect 702 24388 852 24449
rect 702 24342 806 24388
rect 702 24281 852 24342
rect 702 24235 806 24281
rect 702 24174 852 24235
rect 702 24128 806 24174
rect 702 24067 852 24128
rect 702 24021 806 24067
rect 702 24008 852 24021
rect 1030 25358 1181 25370
rect 1030 25357 1117 25358
rect 1076 25311 1117 25357
rect 1030 25249 1117 25311
rect 1076 25203 1117 25249
rect 1030 25202 1117 25203
rect 1169 25202 1181 25358
rect 1030 25141 1181 25202
rect 1076 25095 1181 25141
rect 1030 25033 1181 25095
rect 1076 24987 1181 25033
rect 1030 24925 1181 24987
rect 1076 24879 1181 24925
rect 1030 24817 1181 24879
rect 1076 24805 1181 24817
rect 1321 25358 1472 25370
rect 1321 25202 1333 25358
rect 1385 25357 1472 25358
rect 1385 25311 1426 25357
rect 1385 25249 1472 25311
rect 1385 25203 1426 25249
rect 1385 25202 1472 25203
rect 1321 25141 1472 25202
rect 1321 25095 1426 25141
rect 1321 25033 1472 25095
rect 1321 24987 1426 25033
rect 1321 24925 1472 24987
rect 1321 24879 1426 24925
rect 1321 24817 1472 24879
rect 1321 24805 1426 24817
rect 1076 24771 1137 24805
rect 1030 24709 1137 24771
rect 1076 24663 1137 24709
rect 1365 24771 1426 24805
rect 1365 24709 1472 24771
rect 1030 24602 1137 24663
rect 1076 24556 1137 24602
rect 1030 24495 1137 24556
rect 1076 24449 1137 24495
rect 1030 24388 1137 24449
rect 1213 24684 1289 24696
rect 1213 24424 1225 24684
rect 1277 24424 1289 24684
rect 1213 24423 1228 24424
rect 1274 24423 1289 24424
rect 1213 24412 1289 24423
rect 1365 24663 1426 24709
rect 1365 24602 1472 24663
rect 1365 24556 1426 24602
rect 1365 24495 1472 24556
rect 1365 24449 1426 24495
rect 1076 24342 1137 24388
rect 1030 24285 1137 24342
rect 1365 24388 1472 24449
rect 1365 24342 1426 24388
rect 1365 24285 1472 24342
rect 1030 24281 1181 24285
rect 1076 24235 1181 24281
rect 1030 24174 1181 24235
rect 1076 24128 1181 24174
rect 1030 24067 1181 24128
rect 1076 24021 1181 24067
rect 1030 24008 1181 24021
rect 702 23679 772 24008
rect 851 23926 1032 23938
rect 851 23770 909 23926
rect 961 23770 1032 23926
rect 851 23755 1032 23770
rect 1110 23679 1181 24008
rect 702 23666 852 23679
rect 702 23620 806 23666
rect 702 23558 852 23620
rect 702 23512 806 23558
rect 702 23450 852 23512
rect 702 23404 806 23450
rect 702 23342 852 23404
rect 702 23296 806 23342
rect 702 23234 852 23296
rect 702 23188 806 23234
rect 702 23126 852 23188
rect 702 23080 806 23126
rect 702 23018 852 23080
rect 702 22972 806 23018
rect 702 22911 852 22972
rect 702 22865 806 22911
rect 702 22804 852 22865
rect 702 22758 806 22804
rect 702 22697 852 22758
rect 702 22651 806 22697
rect 702 22590 852 22651
rect 702 22544 806 22590
rect 702 22483 852 22544
rect 702 22437 806 22483
rect 702 22376 852 22437
rect 702 22330 806 22376
rect 702 22327 852 22330
rect 806 22247 852 22327
rect 1030 23666 1181 23679
rect 1076 23620 1181 23666
rect 1030 23558 1181 23620
rect 1076 23512 1181 23558
rect 1030 23450 1181 23512
rect 1076 23404 1181 23450
rect 1030 23342 1181 23404
rect 1076 23296 1181 23342
rect 1030 23234 1181 23296
rect 1076 23188 1181 23234
rect 1030 23126 1181 23188
rect 1076 23080 1181 23126
rect 1030 23018 1181 23080
rect 1076 22972 1181 23018
rect 1030 22911 1181 22972
rect 1076 22865 1181 22911
rect 1030 22804 1181 22865
rect 1076 22758 1181 22804
rect 1030 22697 1181 22758
rect 1076 22651 1181 22697
rect 1030 22590 1181 22651
rect 1076 22544 1181 22590
rect 1030 22483 1181 22544
rect 1076 22437 1181 22483
rect 1030 22376 1181 22437
rect 1076 22330 1181 22376
rect 1030 22317 1181 22330
rect 1321 24281 1472 24285
rect 1321 24235 1426 24281
rect 1321 24174 1472 24235
rect 1321 24128 1426 24174
rect 1321 24067 1472 24128
rect 1321 24021 1426 24067
rect 1321 24008 1472 24021
rect 1650 25357 1800 25370
rect 1696 25311 1800 25357
rect 1650 25249 1800 25311
rect 1696 25203 1800 25249
rect 1650 25141 1800 25203
rect 1696 25095 1800 25141
rect 1650 25033 1800 25095
rect 1696 24987 1800 25033
rect 1650 24925 1800 24987
rect 1696 24879 1800 24925
rect 1650 24817 1800 24879
rect 1696 24771 1800 24817
rect 1650 24709 1800 24771
rect 1696 24663 1800 24709
rect 1650 24602 1800 24663
rect 1696 24556 1800 24602
rect 1650 24495 1800 24556
rect 1696 24449 1800 24495
rect 1650 24388 1800 24449
rect 1696 24342 1800 24388
rect 1650 24281 1800 24342
rect 1696 24235 1800 24281
rect 1650 24174 1800 24235
rect 1696 24128 1800 24174
rect 1650 24067 1800 24128
rect 1696 24021 1800 24067
rect 1650 24008 1800 24021
rect 1321 23679 1392 24008
rect 1470 23926 1651 23938
rect 1470 23770 1541 23926
rect 1593 23770 1651 23926
rect 1470 23755 1651 23770
rect 1730 23679 1800 24008
rect 1321 23666 1472 23679
rect 1321 23620 1426 23666
rect 1321 23558 1472 23620
rect 1321 23512 1426 23558
rect 1321 23450 1472 23512
rect 1321 23404 1426 23450
rect 1321 23342 1472 23404
rect 1321 23296 1426 23342
rect 1321 23234 1472 23296
rect 1321 23188 1426 23234
rect 1321 23126 1472 23188
rect 1321 23080 1426 23126
rect 1321 23018 1472 23080
rect 1321 22972 1426 23018
rect 1321 22911 1472 22972
rect 1321 22865 1426 22911
rect 1321 22804 1472 22865
rect 1321 22758 1426 22804
rect 1321 22697 1472 22758
rect 1321 22651 1426 22697
rect 1321 22590 1472 22651
rect 1321 22544 1426 22590
rect 1321 22483 1472 22544
rect 1321 22437 1426 22483
rect 1321 22376 1472 22437
rect 1321 22330 1426 22376
rect 1321 22317 1472 22330
rect 1650 23666 1800 23679
rect 1696 23620 1800 23666
rect 1650 23558 1800 23620
rect 1696 23512 1800 23558
rect 1650 23450 1800 23512
rect 1696 23404 1800 23450
rect 1650 23342 1800 23404
rect 1696 23296 1800 23342
rect 1650 23234 1800 23296
rect 1696 23188 1800 23234
rect 1650 23126 1800 23188
rect 1696 23080 1800 23126
rect 1650 23018 1800 23080
rect 1696 22972 1800 23018
rect 1650 22911 1800 22972
rect 1696 22865 1800 22911
rect 1650 22804 1800 22865
rect 1696 22758 1800 22804
rect 1650 22697 1800 22758
rect 1696 22651 1800 22697
rect 1650 22590 1800 22651
rect 1696 22544 1800 22590
rect 1650 22483 1800 22544
rect 1696 22437 1800 22483
rect 1650 22376 1800 22437
rect 1696 22330 1800 22376
rect 1650 22327 1800 22330
rect 1941 25357 2091 25370
rect 1941 25311 2045 25357
rect 1941 25249 2091 25311
rect 1941 25203 2045 25249
rect 1941 25141 2091 25203
rect 1941 25095 2045 25141
rect 1941 25033 2091 25095
rect 1941 24987 2045 25033
rect 1941 24925 2091 24987
rect 1941 24879 2045 24925
rect 1941 24817 2091 24879
rect 1941 24771 2045 24817
rect 1941 24709 2091 24771
rect 1941 24663 2045 24709
rect 1941 24602 2091 24663
rect 1941 24556 2045 24602
rect 1941 24495 2091 24556
rect 1941 24449 2045 24495
rect 1941 24388 2091 24449
rect 1941 24342 2045 24388
rect 1941 24281 2091 24342
rect 1941 24235 2045 24281
rect 1941 24174 2091 24235
rect 1941 24128 2045 24174
rect 1941 24067 2091 24128
rect 1941 24021 2045 24067
rect 1941 24008 2091 24021
rect 2269 25358 2420 25370
rect 2269 25357 2356 25358
rect 2315 25311 2356 25357
rect 2269 25249 2356 25311
rect 2315 25203 2356 25249
rect 2269 25202 2356 25203
rect 2408 25202 2420 25358
rect 2269 25141 2420 25202
rect 2315 25095 2420 25141
rect 2269 25033 2420 25095
rect 2315 24987 2420 25033
rect 2269 24925 2420 24987
rect 2315 24879 2420 24925
rect 2269 24817 2420 24879
rect 2315 24805 2420 24817
rect 2560 25358 2711 25370
rect 2560 25202 2572 25358
rect 2624 25357 2711 25358
rect 2624 25311 2665 25357
rect 2624 25249 2711 25311
rect 2624 25203 2665 25249
rect 2624 25202 2711 25203
rect 2560 25141 2711 25202
rect 2560 25095 2665 25141
rect 2560 25033 2711 25095
rect 2560 24987 2665 25033
rect 2560 24925 2711 24987
rect 2560 24879 2665 24925
rect 2560 24817 2711 24879
rect 2560 24805 2665 24817
rect 2315 24771 2376 24805
rect 2269 24709 2376 24771
rect 2315 24663 2376 24709
rect 2604 24771 2665 24805
rect 2604 24709 2711 24771
rect 2269 24602 2376 24663
rect 2315 24556 2376 24602
rect 2269 24495 2376 24556
rect 2315 24449 2376 24495
rect 2269 24388 2376 24449
rect 2452 24684 2528 24696
rect 2452 24424 2464 24684
rect 2516 24424 2528 24684
rect 2452 24423 2467 24424
rect 2513 24423 2528 24424
rect 2452 24412 2528 24423
rect 2604 24663 2665 24709
rect 2604 24602 2711 24663
rect 2604 24556 2665 24602
rect 2604 24495 2711 24556
rect 2604 24449 2665 24495
rect 2315 24342 2376 24388
rect 2269 24285 2376 24342
rect 2604 24388 2711 24449
rect 2604 24342 2665 24388
rect 2604 24285 2711 24342
rect 2269 24281 2420 24285
rect 2315 24235 2420 24281
rect 2269 24174 2420 24235
rect 2315 24128 2420 24174
rect 2269 24067 2420 24128
rect 2315 24021 2420 24067
rect 2269 24008 2420 24021
rect 1941 23679 2011 24008
rect 2090 23926 2271 23938
rect 2090 23770 2148 23926
rect 2200 23770 2271 23926
rect 2090 23755 2271 23770
rect 2349 23679 2420 24008
rect 1941 23666 2091 23679
rect 1941 23620 2045 23666
rect 1941 23558 2091 23620
rect 1941 23512 2045 23558
rect 1941 23450 2091 23512
rect 1941 23404 2045 23450
rect 1941 23342 2091 23404
rect 1941 23296 2045 23342
rect 1941 23234 2091 23296
rect 1941 23188 2045 23234
rect 1941 23126 2091 23188
rect 1941 23080 2045 23126
rect 1941 23018 2091 23080
rect 1941 22972 2045 23018
rect 1941 22911 2091 22972
rect 1941 22865 2045 22911
rect 1941 22804 2091 22865
rect 1941 22758 2045 22804
rect 1941 22697 2091 22758
rect 1941 22651 2045 22697
rect 1941 22590 2091 22651
rect 1941 22544 2045 22590
rect 1941 22483 2091 22544
rect 1941 22437 2045 22483
rect 1941 22376 2091 22437
rect 1941 22330 2045 22376
rect 1941 22327 2091 22330
rect 1650 22247 1696 22327
rect 806 22225 1206 22247
rect 806 22173 1124 22225
rect 1176 22173 1206 22225
rect 806 22150 1206 22173
rect 1296 22225 1696 22247
rect 1296 22173 1326 22225
rect 1378 22173 1696 22225
rect 1296 22150 1696 22173
rect 2045 22247 2091 22327
rect 2269 23666 2420 23679
rect 2315 23620 2420 23666
rect 2269 23558 2420 23620
rect 2315 23512 2420 23558
rect 2269 23450 2420 23512
rect 2315 23404 2420 23450
rect 2269 23342 2420 23404
rect 2315 23296 2420 23342
rect 2269 23234 2420 23296
rect 2315 23188 2420 23234
rect 2269 23126 2420 23188
rect 2315 23080 2420 23126
rect 2269 23018 2420 23080
rect 2315 22972 2420 23018
rect 2269 22911 2420 22972
rect 2315 22865 2420 22911
rect 2269 22804 2420 22865
rect 2315 22758 2420 22804
rect 2269 22697 2420 22758
rect 2315 22651 2420 22697
rect 2269 22590 2420 22651
rect 2315 22544 2420 22590
rect 2269 22483 2420 22544
rect 2315 22437 2420 22483
rect 2269 22376 2420 22437
rect 2315 22330 2420 22376
rect 2269 22317 2420 22330
rect 2560 24281 2711 24285
rect 2560 24235 2665 24281
rect 2560 24174 2711 24235
rect 2560 24128 2665 24174
rect 2560 24067 2711 24128
rect 2560 24021 2665 24067
rect 2560 24008 2711 24021
rect 2889 25357 3039 25370
rect 2935 25311 3039 25357
rect 2889 25249 3039 25311
rect 2935 25203 3039 25249
rect 2889 25141 3039 25203
rect 2935 25095 3039 25141
rect 2889 25033 3039 25095
rect 2935 24987 3039 25033
rect 2889 24925 3039 24987
rect 2935 24879 3039 24925
rect 2889 24817 3039 24879
rect 2935 24771 3039 24817
rect 2889 24709 3039 24771
rect 2935 24663 3039 24709
rect 2889 24602 3039 24663
rect 2935 24556 3039 24602
rect 2889 24495 3039 24556
rect 2935 24449 3039 24495
rect 2889 24388 3039 24449
rect 2935 24342 3039 24388
rect 2889 24281 3039 24342
rect 2935 24235 3039 24281
rect 2889 24174 3039 24235
rect 2935 24128 3039 24174
rect 2889 24067 3039 24128
rect 2935 24021 3039 24067
rect 2889 24008 3039 24021
rect 2560 23679 2631 24008
rect 2709 23926 2890 23938
rect 2709 23770 2780 23926
rect 2832 23770 2890 23926
rect 2709 23755 2890 23770
rect 2969 23679 3039 24008
rect 2560 23666 2711 23679
rect 2560 23620 2665 23666
rect 2560 23558 2711 23620
rect 2560 23512 2665 23558
rect 2560 23450 2711 23512
rect 2560 23404 2665 23450
rect 2560 23342 2711 23404
rect 2560 23296 2665 23342
rect 2560 23234 2711 23296
rect 2560 23188 2665 23234
rect 2560 23126 2711 23188
rect 2560 23080 2665 23126
rect 2560 23018 2711 23080
rect 2560 22972 2665 23018
rect 2560 22911 2711 22972
rect 2560 22865 2665 22911
rect 2560 22804 2711 22865
rect 2560 22758 2665 22804
rect 2560 22697 2711 22758
rect 2560 22651 2665 22697
rect 2560 22590 2711 22651
rect 2560 22544 2665 22590
rect 2560 22483 2711 22544
rect 2560 22437 2665 22483
rect 2560 22376 2711 22437
rect 2560 22330 2665 22376
rect 2560 22317 2711 22330
rect 2889 23666 3039 23679
rect 2935 23620 3039 23666
rect 2889 23558 3039 23620
rect 2935 23512 3039 23558
rect 2889 23450 3039 23512
rect 2935 23404 3039 23450
rect 2889 23342 3039 23404
rect 2935 23296 3039 23342
rect 2889 23234 3039 23296
rect 2935 23188 3039 23234
rect 2889 23126 3039 23188
rect 2935 23080 3039 23126
rect 2889 23018 3039 23080
rect 2935 22972 3039 23018
rect 2889 22911 3039 22972
rect 2935 22865 3039 22911
rect 2889 22804 3039 22865
rect 2935 22758 3039 22804
rect 2889 22697 3039 22758
rect 2935 22651 3039 22697
rect 2889 22590 3039 22651
rect 2935 22544 3039 22590
rect 2889 22483 3039 22544
rect 2935 22437 3039 22483
rect 2889 22376 3039 22437
rect 2935 22330 3039 22376
rect 2889 22327 3039 22330
rect 3179 25357 3329 25370
rect 3179 25311 3283 25357
rect 3179 25249 3329 25311
rect 3179 25203 3283 25249
rect 3179 25141 3329 25203
rect 3179 25095 3283 25141
rect 3179 25033 3329 25095
rect 3179 24987 3283 25033
rect 3179 24925 3329 24987
rect 3179 24879 3283 24925
rect 3179 24817 3329 24879
rect 3179 24771 3283 24817
rect 3179 24709 3329 24771
rect 3179 24663 3283 24709
rect 3179 24602 3329 24663
rect 3179 24556 3283 24602
rect 3179 24495 3329 24556
rect 3179 24449 3283 24495
rect 3179 24388 3329 24449
rect 3179 24342 3283 24388
rect 3179 24281 3329 24342
rect 3179 24235 3283 24281
rect 3179 24174 3329 24235
rect 3179 24128 3283 24174
rect 3179 24067 3329 24128
rect 3179 24021 3283 24067
rect 3179 24008 3329 24021
rect 3507 25358 3658 25370
rect 3507 25357 3594 25358
rect 3553 25311 3594 25357
rect 3507 25249 3594 25311
rect 3553 25203 3594 25249
rect 3507 25202 3594 25203
rect 3646 25202 3658 25358
rect 3507 25141 3658 25202
rect 3553 25095 3658 25141
rect 3507 25033 3658 25095
rect 3553 24987 3658 25033
rect 3507 24925 3658 24987
rect 3553 24879 3658 24925
rect 3507 24817 3658 24879
rect 3553 24805 3658 24817
rect 3798 25358 3949 25370
rect 3798 25202 3810 25358
rect 3862 25357 3949 25358
rect 3862 25311 3903 25357
rect 3862 25249 3949 25311
rect 3862 25203 3903 25249
rect 3862 25202 3949 25203
rect 3798 25141 3949 25202
rect 3798 25095 3903 25141
rect 3798 25033 3949 25095
rect 3798 24987 3903 25033
rect 3798 24925 3949 24987
rect 3798 24879 3903 24925
rect 3798 24817 3949 24879
rect 3798 24805 3903 24817
rect 3553 24771 3614 24805
rect 3507 24709 3614 24771
rect 3553 24663 3614 24709
rect 3842 24771 3903 24805
rect 3842 24709 3949 24771
rect 3507 24602 3614 24663
rect 3553 24556 3614 24602
rect 3507 24495 3614 24556
rect 3553 24449 3614 24495
rect 3507 24388 3614 24449
rect 3690 24684 3766 24696
rect 3690 24424 3702 24684
rect 3754 24424 3766 24684
rect 3690 24423 3705 24424
rect 3751 24423 3766 24424
rect 3690 24412 3766 24423
rect 3842 24663 3903 24709
rect 3842 24602 3949 24663
rect 3842 24556 3903 24602
rect 3842 24495 3949 24556
rect 3842 24449 3903 24495
rect 3553 24342 3614 24388
rect 3507 24285 3614 24342
rect 3842 24388 3949 24449
rect 3842 24342 3903 24388
rect 3842 24285 3949 24342
rect 3507 24281 3658 24285
rect 3553 24235 3658 24281
rect 3507 24174 3658 24235
rect 3553 24128 3658 24174
rect 3507 24067 3658 24128
rect 3553 24021 3658 24067
rect 3507 24008 3658 24021
rect 3179 23679 3249 24008
rect 3328 23926 3509 23938
rect 3328 23770 3386 23926
rect 3438 23770 3509 23926
rect 3328 23755 3509 23770
rect 3587 23679 3658 24008
rect 3179 23666 3329 23679
rect 3179 23620 3283 23666
rect 3179 23558 3329 23620
rect 3179 23512 3283 23558
rect 3179 23450 3329 23512
rect 3179 23404 3283 23450
rect 3179 23342 3329 23404
rect 3179 23296 3283 23342
rect 3179 23234 3329 23296
rect 3179 23188 3283 23234
rect 3179 23126 3329 23188
rect 3179 23080 3283 23126
rect 3179 23018 3329 23080
rect 3179 22972 3283 23018
rect 3179 22911 3329 22972
rect 3179 22865 3283 22911
rect 3179 22804 3329 22865
rect 3179 22758 3283 22804
rect 3179 22697 3329 22758
rect 3179 22651 3283 22697
rect 3179 22590 3329 22651
rect 3179 22544 3283 22590
rect 3179 22483 3329 22544
rect 3179 22437 3283 22483
rect 3179 22376 3329 22437
rect 3179 22330 3283 22376
rect 3179 22327 3329 22330
rect 2889 22247 2935 22327
rect 2045 22225 2445 22247
rect 2045 22173 2363 22225
rect 2415 22173 2445 22225
rect 2045 22150 2445 22173
rect 2535 22225 2935 22247
rect 2535 22173 2565 22225
rect 2617 22173 2935 22225
rect 2535 22150 2935 22173
rect 3283 22247 3329 22327
rect 3507 23666 3658 23679
rect 3553 23620 3658 23666
rect 3507 23558 3658 23620
rect 3553 23512 3658 23558
rect 3507 23450 3658 23512
rect 3553 23404 3658 23450
rect 3507 23342 3658 23404
rect 3553 23296 3658 23342
rect 3507 23234 3658 23296
rect 3553 23188 3658 23234
rect 3507 23126 3658 23188
rect 3553 23080 3658 23126
rect 3507 23018 3658 23080
rect 3553 22972 3658 23018
rect 3507 22911 3658 22972
rect 3553 22865 3658 22911
rect 3507 22804 3658 22865
rect 3553 22758 3658 22804
rect 3507 22697 3658 22758
rect 3553 22651 3658 22697
rect 3507 22590 3658 22651
rect 3553 22544 3658 22590
rect 3507 22483 3658 22544
rect 3553 22437 3658 22483
rect 3507 22376 3658 22437
rect 3553 22330 3658 22376
rect 3507 22317 3658 22330
rect 3798 24281 3949 24285
rect 3798 24235 3903 24281
rect 3798 24174 3949 24235
rect 3798 24128 3903 24174
rect 3798 24067 3949 24128
rect 3798 24021 3903 24067
rect 3798 24008 3949 24021
rect 4127 25357 4277 25370
rect 4173 25311 4277 25357
rect 4127 25249 4277 25311
rect 4173 25203 4277 25249
rect 4127 25141 4277 25203
rect 4173 25095 4277 25141
rect 4127 25033 4277 25095
rect 4173 24987 4277 25033
rect 4127 24925 4277 24987
rect 4173 24879 4277 24925
rect 4127 24817 4277 24879
rect 4173 24771 4277 24817
rect 4127 24709 4277 24771
rect 4173 24663 4277 24709
rect 4127 24602 4277 24663
rect 4173 24556 4277 24602
rect 4127 24495 4277 24556
rect 4173 24449 4277 24495
rect 4127 24388 4277 24449
rect 4173 24342 4277 24388
rect 4127 24281 4277 24342
rect 4173 24235 4277 24281
rect 4127 24174 4277 24235
rect 4173 24128 4277 24174
rect 4127 24067 4277 24128
rect 4173 24021 4277 24067
rect 4127 24008 4277 24021
rect 3798 23679 3869 24008
rect 3947 23926 4128 23938
rect 3947 23770 4018 23926
rect 4070 23770 4128 23926
rect 3947 23755 4128 23770
rect 4207 23679 4277 24008
rect 3798 23666 3949 23679
rect 3798 23620 3903 23666
rect 3798 23558 3949 23620
rect 3798 23512 3903 23558
rect 3798 23450 3949 23512
rect 3798 23404 3903 23450
rect 3798 23342 3949 23404
rect 3798 23296 3903 23342
rect 3798 23234 3949 23296
rect 3798 23188 3903 23234
rect 3798 23126 3949 23188
rect 3798 23080 3903 23126
rect 3798 23018 3949 23080
rect 3798 22972 3903 23018
rect 3798 22911 3949 22972
rect 3798 22865 3903 22911
rect 3798 22804 3949 22865
rect 3798 22758 3903 22804
rect 3798 22697 3949 22758
rect 3798 22651 3903 22697
rect 3798 22590 3949 22651
rect 3798 22544 3903 22590
rect 3798 22483 3949 22544
rect 3798 22437 3903 22483
rect 3798 22376 3949 22437
rect 3798 22330 3903 22376
rect 3798 22317 3949 22330
rect 4127 23666 4277 23679
rect 4173 23620 4277 23666
rect 4127 23558 4277 23620
rect 4173 23512 4277 23558
rect 4127 23450 4277 23512
rect 4173 23404 4277 23450
rect 4127 23342 4277 23404
rect 4173 23296 4277 23342
rect 4127 23234 4277 23296
rect 4173 23188 4277 23234
rect 4127 23126 4277 23188
rect 4173 23080 4277 23126
rect 4127 23018 4277 23080
rect 4173 22972 4277 23018
rect 4127 22911 4277 22972
rect 4173 22865 4277 22911
rect 4127 22804 4277 22865
rect 4173 22758 4277 22804
rect 4127 22697 4277 22758
rect 4173 22651 4277 22697
rect 4127 22590 4277 22651
rect 4173 22544 4277 22590
rect 4127 22483 4277 22544
rect 4173 22437 4277 22483
rect 4127 22376 4277 22437
rect 4173 22330 4277 22376
rect 4127 22327 4277 22330
rect 4418 25357 4568 25370
rect 4418 25311 4522 25357
rect 4418 25249 4568 25311
rect 4418 25203 4522 25249
rect 4418 25141 4568 25203
rect 4418 25095 4522 25141
rect 4418 25033 4568 25095
rect 4418 24987 4522 25033
rect 4418 24925 4568 24987
rect 4418 24879 4522 24925
rect 4418 24817 4568 24879
rect 4418 24771 4522 24817
rect 4418 24709 4568 24771
rect 4418 24663 4522 24709
rect 4418 24602 4568 24663
rect 4418 24556 4522 24602
rect 4418 24495 4568 24556
rect 4418 24449 4522 24495
rect 4418 24388 4568 24449
rect 4418 24342 4522 24388
rect 4418 24281 4568 24342
rect 4418 24235 4522 24281
rect 4418 24174 4568 24235
rect 4418 24128 4522 24174
rect 4418 24067 4568 24128
rect 4418 24021 4522 24067
rect 4418 24008 4568 24021
rect 4746 25358 4897 25370
rect 4746 25357 4833 25358
rect 4792 25311 4833 25357
rect 4746 25249 4833 25311
rect 4792 25203 4833 25249
rect 4746 25202 4833 25203
rect 4885 25202 4897 25358
rect 4746 25141 4897 25202
rect 4792 25095 4897 25141
rect 4746 25033 4897 25095
rect 4792 24987 4897 25033
rect 4746 24925 4897 24987
rect 4792 24879 4897 24925
rect 4746 24817 4897 24879
rect 4792 24805 4897 24817
rect 5041 25358 5188 25370
rect 5041 25202 5053 25358
rect 5105 25357 5188 25358
rect 5105 25311 5142 25357
rect 5105 25249 5188 25311
rect 5105 25203 5142 25249
rect 5105 25202 5188 25203
rect 5041 25141 5188 25202
rect 5041 25095 5142 25141
rect 5041 25033 5188 25095
rect 5041 24987 5142 25033
rect 5041 24925 5188 24987
rect 5041 24879 5142 24925
rect 5041 24817 5188 24879
rect 5041 24805 5142 24817
rect 4792 24771 4853 24805
rect 4746 24709 4853 24771
rect 4792 24663 4853 24709
rect 5081 24771 5142 24805
rect 5081 24709 5188 24771
rect 4746 24602 4853 24663
rect 4792 24556 4853 24602
rect 4746 24495 4853 24556
rect 4792 24449 4853 24495
rect 4746 24388 4853 24449
rect 4929 24684 5005 24696
rect 4929 24424 4941 24684
rect 4993 24424 5005 24684
rect 4929 24423 4944 24424
rect 4990 24423 5005 24424
rect 4929 24412 5005 24423
rect 5081 24663 5142 24709
rect 5081 24602 5188 24663
rect 5081 24556 5142 24602
rect 5081 24495 5188 24556
rect 5081 24449 5142 24495
rect 4792 24342 4853 24388
rect 4746 24285 4853 24342
rect 5081 24388 5188 24449
rect 5081 24342 5142 24388
rect 5081 24285 5188 24342
rect 4746 24281 4897 24285
rect 4792 24235 4897 24281
rect 4746 24174 4897 24235
rect 4792 24128 4897 24174
rect 4746 24067 4897 24128
rect 4792 24021 4897 24067
rect 4746 24008 4897 24021
rect 4418 23679 4488 24008
rect 4567 23926 4748 23938
rect 4567 23770 4625 23926
rect 4677 23770 4748 23926
rect 4567 23755 4748 23770
rect 4826 23679 4897 24008
rect 4418 23666 4568 23679
rect 4418 23620 4522 23666
rect 4418 23558 4568 23620
rect 4418 23512 4522 23558
rect 4418 23450 4568 23512
rect 4418 23404 4522 23450
rect 4418 23342 4568 23404
rect 4418 23296 4522 23342
rect 4418 23234 4568 23296
rect 4418 23188 4522 23234
rect 4418 23126 4568 23188
rect 4418 23080 4522 23126
rect 4418 23018 4568 23080
rect 4418 22972 4522 23018
rect 4418 22911 4568 22972
rect 4418 22865 4522 22911
rect 4418 22804 4568 22865
rect 4418 22758 4522 22804
rect 4418 22697 4568 22758
rect 4418 22651 4522 22697
rect 4418 22590 4568 22651
rect 4418 22544 4522 22590
rect 4418 22483 4568 22544
rect 4418 22437 4522 22483
rect 4418 22376 4568 22437
rect 4418 22330 4522 22376
rect 4418 22327 4568 22330
rect 4127 22247 4173 22327
rect 3283 22225 3683 22247
rect 3283 22173 3601 22225
rect 3653 22173 3683 22225
rect 3283 22150 3683 22173
rect 3773 22225 4173 22247
rect 3773 22173 3803 22225
rect 3855 22173 4173 22225
rect 3773 22150 4173 22173
rect 4522 22247 4568 22327
rect 4746 23666 4897 23679
rect 4792 23620 4897 23666
rect 4746 23558 4897 23620
rect 4792 23512 4897 23558
rect 4746 23450 4897 23512
rect 4792 23404 4897 23450
rect 4746 23342 4897 23404
rect 4792 23296 4897 23342
rect 4746 23234 4897 23296
rect 4792 23188 4897 23234
rect 4746 23126 4897 23188
rect 4792 23080 4897 23126
rect 4746 23018 4897 23080
rect 4792 22972 4897 23018
rect 4746 22911 4897 22972
rect 4792 22865 4897 22911
rect 4746 22804 4897 22865
rect 4792 22758 4897 22804
rect 4746 22697 4897 22758
rect 4792 22651 4897 22697
rect 4746 22590 4897 22651
rect 4792 22544 4897 22590
rect 4746 22483 4897 22544
rect 4792 22437 4897 22483
rect 4746 22376 4897 22437
rect 4792 22330 4897 22376
rect 4746 22317 4897 22330
rect 5041 24281 5188 24285
rect 5041 24235 5142 24281
rect 5041 24174 5188 24235
rect 5041 24128 5142 24174
rect 5041 24067 5188 24128
rect 5041 24021 5142 24067
rect 5041 24008 5188 24021
rect 5366 25362 5412 25370
rect 5366 25357 5517 25362
rect 5412 25311 5517 25357
rect 5366 25249 5517 25311
rect 5412 25203 5517 25249
rect 5366 25141 5517 25203
rect 5412 25095 5517 25141
rect 5366 25033 5517 25095
rect 5412 24987 5517 25033
rect 5366 24925 5517 24987
rect 5412 24879 5517 24925
rect 5366 24817 5517 24879
rect 5412 24771 5517 24817
rect 5366 24709 5517 24771
rect 5412 24663 5517 24709
rect 5366 24602 5517 24663
rect 5412 24556 5517 24602
rect 5366 24495 5517 24556
rect 5412 24449 5517 24495
rect 5366 24388 5517 24449
rect 5412 24342 5517 24388
rect 5366 24281 5517 24342
rect 5412 24235 5517 24281
rect 5366 24174 5517 24235
rect 5412 24128 5517 24174
rect 5366 24067 5517 24128
rect 5412 24021 5517 24067
rect 5366 24008 5517 24021
rect 5041 23679 5129 24008
rect 5186 23926 5368 23938
rect 5186 23770 5257 23926
rect 5309 23770 5368 23926
rect 5186 23755 5368 23770
rect 5425 23679 5517 24008
rect 5041 23666 5188 23679
rect 5041 23620 5142 23666
rect 5041 23558 5188 23620
rect 5041 23512 5142 23558
rect 5041 23450 5188 23512
rect 5041 23404 5142 23450
rect 5041 23342 5188 23404
rect 5041 23296 5142 23342
rect 5041 23234 5188 23296
rect 5041 23188 5142 23234
rect 5041 23126 5188 23188
rect 5041 23080 5142 23126
rect 5041 23018 5188 23080
rect 5041 22972 5142 23018
rect 5041 22911 5188 22972
rect 5041 22865 5142 22911
rect 5041 22804 5188 22865
rect 5041 22758 5142 22804
rect 5041 22697 5188 22758
rect 5041 22651 5142 22697
rect 5041 22590 5188 22651
rect 5041 22544 5142 22590
rect 5041 22483 5188 22544
rect 5041 22437 5142 22483
rect 5041 22376 5188 22437
rect 5041 22330 5142 22376
rect 5041 22327 5188 22330
rect 5142 22317 5188 22327
rect 5366 23666 5517 23679
rect 5412 23620 5517 23666
rect 5366 23558 5517 23620
rect 5412 23512 5517 23558
rect 5366 23450 5517 23512
rect 5412 23404 5517 23450
rect 5366 23342 5517 23404
rect 5412 23296 5517 23342
rect 5366 23234 5517 23296
rect 5412 23188 5517 23234
rect 5366 23126 5517 23188
rect 5412 23080 5517 23126
rect 5366 23018 5517 23080
rect 5412 22972 5517 23018
rect 5366 22911 5517 22972
rect 5412 22865 5517 22911
rect 5366 22804 5517 22865
rect 5412 22758 5517 22804
rect 5366 22697 5517 22758
rect 5412 22651 5517 22697
rect 5366 22590 5517 22651
rect 5412 22544 5517 22590
rect 5366 22483 5517 22544
rect 5412 22437 5517 22483
rect 5366 22376 5517 22437
rect 5412 22330 5517 22376
rect 5366 22327 5517 22330
rect 5366 22247 5412 22327
rect 4522 22225 4922 22247
rect 4522 22173 4840 22225
rect 4892 22173 4922 22225
rect 4522 22150 4922 22173
rect 5012 22225 5412 22247
rect 5012 22173 5042 22225
rect 5094 22173 5412 22225
rect 5012 22150 5412 22173
rect 1180 22066 1322 22071
rect 2419 22066 2561 22071
rect 3657 22066 3799 22071
rect 4896 22066 5038 22071
rect 5516 22066 5658 22071
rect 631 22027 5658 22066
rect 631 21975 831 22027
rect 883 22020 1619 22027
rect 883 21975 1228 22020
rect 631 21974 1228 21975
rect 1274 21975 1619 22020
rect 1671 21975 2070 22027
rect 2122 22020 2858 22027
rect 2122 21975 2467 22020
rect 1274 21974 2467 21975
rect 2513 21975 2858 22020
rect 2910 21975 3308 22027
rect 3360 22020 4096 22027
rect 3360 21975 3705 22020
rect 2513 21974 3705 21975
rect 3751 21975 4096 22020
rect 4148 21975 4547 22027
rect 4599 22020 5314 22027
rect 4599 21975 4944 22020
rect 3751 21974 4944 21975
rect 4990 21975 5314 22020
rect 5366 22020 5658 22027
rect 5366 21975 5564 22020
rect 4990 21974 5564 21975
rect 5610 21974 5658 22020
rect 631 21932 5658 21974
rect 1180 21923 1322 21932
rect 2419 21923 2561 21932
rect 3657 21923 3799 21932
rect 4896 21923 5038 21932
rect 5516 21923 5658 21932
rect 686 21819 1203 21844
rect 686 21767 699 21819
rect 751 21767 1203 21819
rect 686 21747 1203 21767
rect 1110 21675 1203 21747
rect 806 21667 852 21675
rect 702 21662 852 21667
rect 702 21616 806 21662
rect 702 21554 852 21616
rect 702 21508 806 21554
rect 702 21446 852 21508
rect 702 21400 806 21446
rect 702 21338 852 21400
rect 702 21292 806 21338
rect 702 21230 852 21292
rect 702 21184 806 21230
rect 702 21122 852 21184
rect 702 21076 806 21122
rect 702 21014 852 21076
rect 702 20968 806 21014
rect 702 20907 852 20968
rect 702 20861 806 20907
rect 702 20800 852 20861
rect 702 20754 806 20800
rect 702 20693 852 20754
rect 702 20647 806 20693
rect 702 20586 852 20647
rect 702 20540 806 20586
rect 702 20479 852 20540
rect 702 20433 806 20479
rect 702 20372 852 20433
rect 702 20326 806 20372
rect 702 20313 852 20326
rect 1030 21662 1203 21675
rect 1076 21616 1203 21662
rect 1030 21554 1203 21616
rect 1076 21508 1203 21554
rect 1030 21446 1203 21508
rect 1076 21400 1203 21446
rect 1030 21338 1203 21400
rect 1076 21292 1203 21338
rect 1030 21230 1203 21292
rect 1076 21184 1203 21230
rect 1030 21122 1203 21184
rect 1076 21076 1203 21122
rect 1030 21014 1203 21076
rect 1076 20968 1203 21014
rect 1030 20907 1203 20968
rect 1076 20861 1203 20907
rect 1030 20800 1203 20861
rect 1076 20754 1203 20800
rect 1030 20693 1203 20754
rect 1076 20647 1203 20693
rect 1030 20586 1203 20647
rect 1076 20540 1203 20586
rect 1030 20479 1203 20540
rect 1076 20433 1203 20479
rect 1030 20372 1203 20433
rect 1076 20326 1203 20372
rect 1030 20313 1203 20326
rect 702 19820 772 20313
rect 851 20229 1032 20243
rect 851 20219 918 20229
rect 964 20219 1032 20229
rect 851 20167 913 20219
rect 965 20167 1032 20219
rect 851 20108 1032 20167
rect 851 19955 1032 20028
rect 851 19903 915 19955
rect 967 19903 1032 19955
rect 851 19892 1032 19903
rect 903 19891 979 19892
rect 1110 19820 1203 20313
rect 702 19807 852 19820
rect 702 19761 806 19807
rect 702 19699 852 19761
rect 702 19653 806 19699
rect 702 19591 852 19653
rect 702 19545 806 19591
rect 702 19483 852 19545
rect 702 19437 806 19483
rect 702 19375 852 19437
rect 702 19329 806 19375
rect 702 19267 852 19329
rect 702 19221 806 19267
rect 702 19159 852 19221
rect 702 19113 806 19159
rect 702 19052 852 19113
rect 702 19006 806 19052
rect 702 18945 852 19006
rect 702 18899 806 18945
rect 702 18838 852 18899
rect 702 18792 806 18838
rect 702 18731 852 18792
rect 702 18685 806 18731
rect 702 18624 852 18685
rect 702 18578 806 18624
rect 702 18517 852 18578
rect 702 18471 806 18517
rect 702 18470 852 18471
rect 1030 19807 1203 19820
rect 1076 19761 1203 19807
rect 1030 19699 1203 19761
rect 1076 19653 1203 19699
rect 1030 19591 1203 19653
rect 1076 19545 1203 19591
rect 1030 19483 1203 19545
rect 1076 19437 1203 19483
rect 1030 19375 1203 19437
rect 1076 19329 1203 19375
rect 1030 19267 1203 19329
rect 1076 19221 1203 19267
rect 1030 19159 1203 19221
rect 1076 19113 1203 19159
rect 1030 19052 1203 19113
rect 1076 19006 1203 19052
rect 1030 18945 1203 19006
rect 1076 18899 1203 18945
rect 1030 18838 1203 18899
rect 1076 18792 1203 18838
rect 1030 18731 1203 18792
rect 1076 18685 1203 18731
rect 1030 18624 1203 18685
rect 1076 18578 1203 18624
rect 1030 18517 1203 18578
rect 1076 18471 1203 18517
rect 702 18378 887 18470
rect 1030 18468 1203 18471
rect 1299 21819 1816 21844
rect 1299 21767 1751 21819
rect 1803 21767 1816 21819
rect 1299 21747 1816 21767
rect 1925 21819 2442 21844
rect 1925 21767 1938 21819
rect 1990 21767 2442 21819
rect 1925 21747 2442 21767
rect 1299 21675 1392 21747
rect 2349 21675 2442 21747
rect 1299 21662 1472 21675
rect 1299 21616 1426 21662
rect 1299 21554 1472 21616
rect 1299 21508 1426 21554
rect 1299 21446 1472 21508
rect 1299 21400 1426 21446
rect 1299 21338 1472 21400
rect 1299 21292 1426 21338
rect 1299 21230 1472 21292
rect 1299 21184 1426 21230
rect 1299 21122 1472 21184
rect 1299 21076 1426 21122
rect 1299 21014 1472 21076
rect 1299 20968 1426 21014
rect 1299 20907 1472 20968
rect 1299 20861 1426 20907
rect 1299 20800 1472 20861
rect 1299 20754 1426 20800
rect 1299 20693 1472 20754
rect 1299 20647 1426 20693
rect 1299 20586 1472 20647
rect 1299 20540 1426 20586
rect 1299 20479 1472 20540
rect 1299 20433 1426 20479
rect 1299 20372 1472 20433
rect 1299 20326 1426 20372
rect 1299 20313 1472 20326
rect 1650 21667 1696 21675
rect 2045 21667 2091 21675
rect 1650 21662 1800 21667
rect 1696 21616 1800 21662
rect 1650 21554 1800 21616
rect 1696 21508 1800 21554
rect 1650 21446 1800 21508
rect 1696 21400 1800 21446
rect 1650 21338 1800 21400
rect 1696 21292 1800 21338
rect 1650 21230 1800 21292
rect 1696 21184 1800 21230
rect 1650 21122 1800 21184
rect 1696 21076 1800 21122
rect 1650 21014 1800 21076
rect 1696 20968 1800 21014
rect 1650 20907 1800 20968
rect 1696 20861 1800 20907
rect 1650 20800 1800 20861
rect 1696 20754 1800 20800
rect 1650 20693 1800 20754
rect 1696 20647 1800 20693
rect 1650 20586 1800 20647
rect 1696 20540 1800 20586
rect 1650 20479 1800 20540
rect 1696 20433 1800 20479
rect 1650 20372 1800 20433
rect 1696 20326 1800 20372
rect 1650 20313 1800 20326
rect 1299 19820 1392 20313
rect 1470 20229 1651 20243
rect 1470 20219 1538 20229
rect 1584 20219 1651 20229
rect 1470 20167 1537 20219
rect 1589 20167 1651 20219
rect 1470 20108 1651 20167
rect 1470 19955 1651 20028
rect 1470 19903 1535 19955
rect 1587 19903 1651 19955
rect 1470 19892 1651 19903
rect 1523 19891 1599 19892
rect 1730 19820 1800 20313
rect 1299 19807 1472 19820
rect 1299 19761 1426 19807
rect 1299 19699 1472 19761
rect 1299 19653 1426 19699
rect 1299 19591 1472 19653
rect 1299 19545 1426 19591
rect 1299 19483 1472 19545
rect 1299 19437 1426 19483
rect 1299 19375 1472 19437
rect 1299 19329 1426 19375
rect 1299 19267 1472 19329
rect 1299 19221 1426 19267
rect 1299 19159 1472 19221
rect 1299 19113 1426 19159
rect 1299 19052 1472 19113
rect 1299 19006 1426 19052
rect 1299 18945 1472 19006
rect 1299 18899 1426 18945
rect 1299 18838 1472 18899
rect 1299 18792 1426 18838
rect 1299 18731 1472 18792
rect 1299 18685 1426 18731
rect 1299 18624 1472 18685
rect 1299 18578 1426 18624
rect 1299 18517 1472 18578
rect 1299 18471 1426 18517
rect 1299 18468 1472 18471
rect 1650 19807 1800 19820
rect 1696 19761 1800 19807
rect 1650 19699 1800 19761
rect 1696 19653 1800 19699
rect 1650 19591 1800 19653
rect 1696 19545 1800 19591
rect 1650 19483 1800 19545
rect 1696 19437 1800 19483
rect 1650 19375 1800 19437
rect 1696 19329 1800 19375
rect 1650 19267 1800 19329
rect 1696 19221 1800 19267
rect 1650 19159 1800 19221
rect 1696 19113 1800 19159
rect 1650 19052 1800 19113
rect 1696 19006 1800 19052
rect 1650 18945 1800 19006
rect 1696 18899 1800 18945
rect 1650 18838 1800 18899
rect 1696 18792 1800 18838
rect 1650 18731 1800 18792
rect 1696 18685 1800 18731
rect 1650 18624 1800 18685
rect 1696 18578 1800 18624
rect 1650 18517 1800 18578
rect 1696 18471 1800 18517
rect 1650 18470 1800 18471
rect 1030 18458 1076 18468
rect 1426 18458 1472 18468
rect 702 18326 714 18378
rect 766 18326 887 18378
rect 702 18314 887 18326
rect 1615 18406 1800 18470
rect 1941 21662 2091 21667
rect 1941 21616 2045 21662
rect 1941 21554 2091 21616
rect 1941 21508 2045 21554
rect 1941 21446 2091 21508
rect 1941 21400 2045 21446
rect 1941 21338 2091 21400
rect 1941 21292 2045 21338
rect 1941 21230 2091 21292
rect 1941 21184 2045 21230
rect 1941 21122 2091 21184
rect 1941 21076 2045 21122
rect 1941 21014 2091 21076
rect 1941 20968 2045 21014
rect 1941 20907 2091 20968
rect 1941 20861 2045 20907
rect 1941 20800 2091 20861
rect 1941 20754 2045 20800
rect 1941 20693 2091 20754
rect 1941 20647 2045 20693
rect 1941 20586 2091 20647
rect 1941 20540 2045 20586
rect 1941 20479 2091 20540
rect 1941 20433 2045 20479
rect 1941 20372 2091 20433
rect 1941 20326 2045 20372
rect 1941 20313 2091 20326
rect 2269 21662 2442 21675
rect 2315 21616 2442 21662
rect 2269 21554 2442 21616
rect 2315 21508 2442 21554
rect 2269 21446 2442 21508
rect 2315 21400 2442 21446
rect 2269 21338 2442 21400
rect 2315 21292 2442 21338
rect 2269 21230 2442 21292
rect 2315 21184 2442 21230
rect 2269 21122 2442 21184
rect 2315 21076 2442 21122
rect 2269 21014 2442 21076
rect 2315 20968 2442 21014
rect 2269 20907 2442 20968
rect 2315 20861 2442 20907
rect 2269 20800 2442 20861
rect 2315 20754 2442 20800
rect 2269 20693 2442 20754
rect 2315 20647 2442 20693
rect 2269 20586 2442 20647
rect 2315 20540 2442 20586
rect 2269 20479 2442 20540
rect 2315 20433 2442 20479
rect 2269 20372 2442 20433
rect 2315 20326 2442 20372
rect 2269 20313 2442 20326
rect 1941 19820 2011 20313
rect 2090 20229 2271 20243
rect 2090 20219 2157 20229
rect 2203 20219 2271 20229
rect 2090 20167 2152 20219
rect 2204 20167 2271 20219
rect 2090 20108 2271 20167
rect 2090 19955 2271 20028
rect 2090 19903 2154 19955
rect 2206 19903 2271 19955
rect 2090 19892 2271 19903
rect 2142 19891 2218 19892
rect 2349 19820 2442 20313
rect 1941 19807 2091 19820
rect 1941 19761 2045 19807
rect 1941 19699 2091 19761
rect 1941 19653 2045 19699
rect 1941 19591 2091 19653
rect 1941 19545 2045 19591
rect 1941 19483 2091 19545
rect 1941 19437 2045 19483
rect 1941 19375 2091 19437
rect 1941 19329 2045 19375
rect 1941 19267 2091 19329
rect 1941 19221 2045 19267
rect 1941 19159 2091 19221
rect 1941 19113 2045 19159
rect 1941 19052 2091 19113
rect 1941 19006 2045 19052
rect 1941 18945 2091 19006
rect 1941 18899 2045 18945
rect 1941 18838 2091 18899
rect 1941 18792 2045 18838
rect 1941 18731 2091 18792
rect 1941 18685 2045 18731
rect 1941 18624 2091 18685
rect 1941 18578 2045 18624
rect 1941 18517 2091 18578
rect 1941 18471 2045 18517
rect 1941 18470 2091 18471
rect 2269 19807 2442 19820
rect 2315 19761 2442 19807
rect 2269 19699 2442 19761
rect 2315 19653 2442 19699
rect 2269 19591 2442 19653
rect 2315 19545 2442 19591
rect 2269 19483 2442 19545
rect 2315 19437 2442 19483
rect 2269 19375 2442 19437
rect 2315 19329 2442 19375
rect 2269 19267 2442 19329
rect 2315 19221 2442 19267
rect 2269 19159 2442 19221
rect 2315 19113 2442 19159
rect 2269 19052 2442 19113
rect 2315 19006 2442 19052
rect 2269 18945 2442 19006
rect 2315 18899 2442 18945
rect 2269 18838 2442 18899
rect 2315 18792 2442 18838
rect 2269 18731 2442 18792
rect 2315 18685 2442 18731
rect 2269 18624 2442 18685
rect 2315 18578 2442 18624
rect 2269 18517 2442 18578
rect 2315 18471 2442 18517
rect 1941 18406 2126 18470
rect 2269 18468 2442 18471
rect 2538 21819 3055 21844
rect 2538 21767 2990 21819
rect 3042 21767 3055 21819
rect 2538 21747 3055 21767
rect 3163 21819 3680 21844
rect 3163 21767 3176 21819
rect 3228 21767 3680 21819
rect 3163 21747 3680 21767
rect 2538 21675 2631 21747
rect 3587 21675 3680 21747
rect 2538 21662 2711 21675
rect 2538 21616 2665 21662
rect 2538 21554 2711 21616
rect 2538 21508 2665 21554
rect 2538 21446 2711 21508
rect 2538 21400 2665 21446
rect 2538 21338 2711 21400
rect 2538 21292 2665 21338
rect 2538 21230 2711 21292
rect 2538 21184 2665 21230
rect 2538 21122 2711 21184
rect 2538 21076 2665 21122
rect 2538 21014 2711 21076
rect 2538 20968 2665 21014
rect 2538 20907 2711 20968
rect 2538 20861 2665 20907
rect 2538 20800 2711 20861
rect 2538 20754 2665 20800
rect 2538 20693 2711 20754
rect 2538 20647 2665 20693
rect 2538 20586 2711 20647
rect 2538 20540 2665 20586
rect 2538 20479 2711 20540
rect 2538 20433 2665 20479
rect 2538 20372 2711 20433
rect 2538 20326 2665 20372
rect 2538 20313 2711 20326
rect 2889 21667 2935 21675
rect 3283 21667 3329 21675
rect 2889 21662 3039 21667
rect 2935 21616 3039 21662
rect 2889 21554 3039 21616
rect 2935 21508 3039 21554
rect 2889 21446 3039 21508
rect 2935 21400 3039 21446
rect 2889 21338 3039 21400
rect 2935 21292 3039 21338
rect 2889 21230 3039 21292
rect 2935 21184 3039 21230
rect 2889 21122 3039 21184
rect 2935 21076 3039 21122
rect 2889 21014 3039 21076
rect 2935 20968 3039 21014
rect 2889 20907 3039 20968
rect 2935 20861 3039 20907
rect 2889 20800 3039 20861
rect 2935 20754 3039 20800
rect 2889 20693 3039 20754
rect 2935 20647 3039 20693
rect 2889 20586 3039 20647
rect 2935 20540 3039 20586
rect 2889 20479 3039 20540
rect 2935 20433 3039 20479
rect 2889 20372 3039 20433
rect 2935 20326 3039 20372
rect 2889 20313 3039 20326
rect 2538 19820 2631 20313
rect 2709 20229 2890 20243
rect 2709 20219 2777 20229
rect 2823 20219 2890 20229
rect 2709 20167 2776 20219
rect 2828 20167 2890 20219
rect 2709 20108 2890 20167
rect 2709 19955 2890 20028
rect 2709 19903 2774 19955
rect 2826 19903 2890 19955
rect 2709 19892 2890 19903
rect 2762 19891 2838 19892
rect 2969 19820 3039 20313
rect 2538 19807 2711 19820
rect 2538 19761 2665 19807
rect 2538 19699 2711 19761
rect 2538 19653 2665 19699
rect 2538 19591 2711 19653
rect 2538 19545 2665 19591
rect 2538 19483 2711 19545
rect 2538 19437 2665 19483
rect 2538 19375 2711 19437
rect 2538 19329 2665 19375
rect 2538 19267 2711 19329
rect 2538 19221 2665 19267
rect 2538 19159 2711 19221
rect 2538 19113 2665 19159
rect 2538 19052 2711 19113
rect 2538 19006 2665 19052
rect 2538 18945 2711 19006
rect 2538 18899 2665 18945
rect 2538 18838 2711 18899
rect 2538 18792 2665 18838
rect 2538 18731 2711 18792
rect 2538 18685 2665 18731
rect 2538 18624 2711 18685
rect 2538 18578 2665 18624
rect 2538 18517 2711 18578
rect 2538 18471 2665 18517
rect 2538 18468 2711 18471
rect 2889 19807 3039 19820
rect 2935 19761 3039 19807
rect 2889 19699 3039 19761
rect 2935 19653 3039 19699
rect 2889 19591 3039 19653
rect 2935 19545 3039 19591
rect 2889 19483 3039 19545
rect 2935 19437 3039 19483
rect 2889 19375 3039 19437
rect 2935 19329 3039 19375
rect 2889 19267 3039 19329
rect 2935 19221 3039 19267
rect 2889 19159 3039 19221
rect 2935 19113 3039 19159
rect 2889 19052 3039 19113
rect 2935 19006 3039 19052
rect 2889 18945 3039 19006
rect 2935 18899 3039 18945
rect 2889 18838 3039 18899
rect 2935 18792 3039 18838
rect 2889 18731 3039 18792
rect 2935 18685 3039 18731
rect 2889 18624 3039 18685
rect 2935 18578 3039 18624
rect 2889 18517 3039 18578
rect 2935 18471 3039 18517
rect 2889 18470 3039 18471
rect 2269 18458 2315 18468
rect 2665 18458 2711 18468
rect 1615 18386 2126 18406
rect 1615 18334 1747 18386
rect 1799 18334 1933 18386
rect 1985 18334 2126 18386
rect 1615 18314 2126 18334
rect 2854 18406 3039 18470
rect 3179 21662 3329 21667
rect 3179 21616 3283 21662
rect 3179 21554 3329 21616
rect 3179 21508 3283 21554
rect 3179 21446 3329 21508
rect 3179 21400 3283 21446
rect 3179 21338 3329 21400
rect 3179 21292 3283 21338
rect 3179 21230 3329 21292
rect 3179 21184 3283 21230
rect 3179 21122 3329 21184
rect 3179 21076 3283 21122
rect 3179 21014 3329 21076
rect 3179 20968 3283 21014
rect 3179 20907 3329 20968
rect 3179 20861 3283 20907
rect 3179 20800 3329 20861
rect 3179 20754 3283 20800
rect 3179 20693 3329 20754
rect 3179 20647 3283 20693
rect 3179 20586 3329 20647
rect 3179 20540 3283 20586
rect 3179 20479 3329 20540
rect 3179 20433 3283 20479
rect 3179 20372 3329 20433
rect 3179 20326 3283 20372
rect 3179 20313 3329 20326
rect 3507 21662 3680 21675
rect 3553 21616 3680 21662
rect 3507 21554 3680 21616
rect 3553 21508 3680 21554
rect 3507 21446 3680 21508
rect 3553 21400 3680 21446
rect 3507 21338 3680 21400
rect 3553 21292 3680 21338
rect 3507 21230 3680 21292
rect 3553 21184 3680 21230
rect 3507 21122 3680 21184
rect 3553 21076 3680 21122
rect 3507 21014 3680 21076
rect 3553 20968 3680 21014
rect 3507 20907 3680 20968
rect 3553 20861 3680 20907
rect 3507 20800 3680 20861
rect 3553 20754 3680 20800
rect 3507 20693 3680 20754
rect 3553 20647 3680 20693
rect 3507 20586 3680 20647
rect 3553 20540 3680 20586
rect 3507 20479 3680 20540
rect 3553 20433 3680 20479
rect 3507 20372 3680 20433
rect 3553 20326 3680 20372
rect 3507 20313 3680 20326
rect 3179 19820 3249 20313
rect 3328 20229 3509 20243
rect 3328 20219 3395 20229
rect 3441 20219 3509 20229
rect 3328 20167 3390 20219
rect 3442 20167 3509 20219
rect 3328 20108 3509 20167
rect 3328 19955 3509 20028
rect 3328 19903 3392 19955
rect 3444 19903 3509 19955
rect 3328 19892 3509 19903
rect 3380 19891 3456 19892
rect 3587 19820 3680 20313
rect 3179 19807 3329 19820
rect 3179 19761 3283 19807
rect 3179 19699 3329 19761
rect 3179 19653 3283 19699
rect 3179 19591 3329 19653
rect 3179 19545 3283 19591
rect 3179 19483 3329 19545
rect 3179 19437 3283 19483
rect 3179 19375 3329 19437
rect 3179 19329 3283 19375
rect 3179 19267 3329 19329
rect 3179 19221 3283 19267
rect 3179 19159 3329 19221
rect 3179 19113 3283 19159
rect 3179 19052 3329 19113
rect 3179 19006 3283 19052
rect 3179 18945 3329 19006
rect 3179 18899 3283 18945
rect 3179 18838 3329 18899
rect 3179 18792 3283 18838
rect 3179 18731 3329 18792
rect 3179 18685 3283 18731
rect 3179 18624 3329 18685
rect 3179 18578 3283 18624
rect 3179 18517 3329 18578
rect 3179 18471 3283 18517
rect 3179 18470 3329 18471
rect 3507 19807 3680 19820
rect 3553 19761 3680 19807
rect 3507 19699 3680 19761
rect 3553 19653 3680 19699
rect 3507 19591 3680 19653
rect 3553 19545 3680 19591
rect 3507 19483 3680 19545
rect 3553 19437 3680 19483
rect 3507 19375 3680 19437
rect 3553 19329 3680 19375
rect 3507 19267 3680 19329
rect 3553 19221 3680 19267
rect 3507 19159 3680 19221
rect 3553 19113 3680 19159
rect 3507 19052 3680 19113
rect 3553 19006 3680 19052
rect 3507 18945 3680 19006
rect 3553 18899 3680 18945
rect 3507 18838 3680 18899
rect 3553 18792 3680 18838
rect 3507 18731 3680 18792
rect 3553 18685 3680 18731
rect 3507 18624 3680 18685
rect 3553 18578 3680 18624
rect 3507 18517 3680 18578
rect 3553 18471 3680 18517
rect 3179 18406 3364 18470
rect 3507 18468 3680 18471
rect 3776 21819 4293 21844
rect 3776 21767 4228 21819
rect 4280 21767 4293 21819
rect 3776 21747 4293 21767
rect 4402 21819 4919 21844
rect 4402 21767 4415 21819
rect 4467 21767 4919 21819
rect 4402 21747 4919 21767
rect 3776 21675 3869 21747
rect 4826 21675 4919 21747
rect 3776 21662 3949 21675
rect 3776 21616 3903 21662
rect 3776 21554 3949 21616
rect 3776 21508 3903 21554
rect 3776 21446 3949 21508
rect 3776 21400 3903 21446
rect 3776 21338 3949 21400
rect 3776 21292 3903 21338
rect 3776 21230 3949 21292
rect 3776 21184 3903 21230
rect 3776 21122 3949 21184
rect 3776 21076 3903 21122
rect 3776 21014 3949 21076
rect 3776 20968 3903 21014
rect 3776 20907 3949 20968
rect 3776 20861 3903 20907
rect 3776 20800 3949 20861
rect 3776 20754 3903 20800
rect 3776 20693 3949 20754
rect 3776 20647 3903 20693
rect 3776 20586 3949 20647
rect 3776 20540 3903 20586
rect 3776 20479 3949 20540
rect 3776 20433 3903 20479
rect 3776 20372 3949 20433
rect 3776 20326 3903 20372
rect 3776 20313 3949 20326
rect 4127 21667 4173 21675
rect 4522 21667 4568 21675
rect 4127 21662 4277 21667
rect 4173 21616 4277 21662
rect 4127 21554 4277 21616
rect 4173 21508 4277 21554
rect 4127 21446 4277 21508
rect 4173 21400 4277 21446
rect 4127 21338 4277 21400
rect 4173 21292 4277 21338
rect 4127 21230 4277 21292
rect 4173 21184 4277 21230
rect 4127 21122 4277 21184
rect 4173 21076 4277 21122
rect 4127 21014 4277 21076
rect 4173 20968 4277 21014
rect 4127 20907 4277 20968
rect 4173 20861 4277 20907
rect 4127 20800 4277 20861
rect 4173 20754 4277 20800
rect 4127 20693 4277 20754
rect 4173 20647 4277 20693
rect 4127 20586 4277 20647
rect 4173 20540 4277 20586
rect 4127 20479 4277 20540
rect 4173 20433 4277 20479
rect 4127 20372 4277 20433
rect 4173 20326 4277 20372
rect 4127 20313 4277 20326
rect 3776 19820 3869 20313
rect 3947 20229 4128 20243
rect 3947 20219 4015 20229
rect 4061 20219 4128 20229
rect 3947 20167 4014 20219
rect 4066 20167 4128 20219
rect 3947 20108 4128 20167
rect 3947 19955 4128 20028
rect 3947 19903 4012 19955
rect 4064 19903 4128 19955
rect 3947 19892 4128 19903
rect 4000 19891 4076 19892
rect 4207 19820 4277 20313
rect 3776 19807 3949 19820
rect 3776 19761 3903 19807
rect 3776 19699 3949 19761
rect 3776 19653 3903 19699
rect 3776 19591 3949 19653
rect 3776 19545 3903 19591
rect 3776 19483 3949 19545
rect 3776 19437 3903 19483
rect 3776 19375 3949 19437
rect 3776 19329 3903 19375
rect 3776 19267 3949 19329
rect 3776 19221 3903 19267
rect 3776 19159 3949 19221
rect 3776 19113 3903 19159
rect 3776 19052 3949 19113
rect 3776 19006 3903 19052
rect 3776 18945 3949 19006
rect 3776 18899 3903 18945
rect 3776 18838 3949 18899
rect 3776 18792 3903 18838
rect 3776 18731 3949 18792
rect 3776 18685 3903 18731
rect 3776 18624 3949 18685
rect 3776 18578 3903 18624
rect 3776 18517 3949 18578
rect 3776 18471 3903 18517
rect 3776 18468 3949 18471
rect 4127 19807 4277 19820
rect 4173 19761 4277 19807
rect 4127 19699 4277 19761
rect 4173 19653 4277 19699
rect 4127 19591 4277 19653
rect 4173 19545 4277 19591
rect 4127 19483 4277 19545
rect 4173 19437 4277 19483
rect 4127 19375 4277 19437
rect 4173 19329 4277 19375
rect 4127 19267 4277 19329
rect 4173 19221 4277 19267
rect 4127 19159 4277 19221
rect 4173 19113 4277 19159
rect 4127 19052 4277 19113
rect 4173 19006 4277 19052
rect 4127 18945 4277 19006
rect 4173 18899 4277 18945
rect 4127 18838 4277 18899
rect 4173 18792 4277 18838
rect 4127 18731 4277 18792
rect 4173 18685 4277 18731
rect 4127 18624 4277 18685
rect 4173 18578 4277 18624
rect 4127 18517 4277 18578
rect 4173 18471 4277 18517
rect 4127 18470 4277 18471
rect 3507 18458 3553 18468
rect 3903 18458 3949 18468
rect 2854 18386 3364 18406
rect 2854 18334 2985 18386
rect 3037 18334 3171 18386
rect 3223 18334 3364 18386
rect 2854 18314 3364 18334
rect 4092 18406 4277 18470
rect 4418 21662 4568 21667
rect 4418 21616 4522 21662
rect 4418 21554 4568 21616
rect 4418 21508 4522 21554
rect 4418 21446 4568 21508
rect 4418 21400 4522 21446
rect 4418 21338 4568 21400
rect 4418 21292 4522 21338
rect 4418 21230 4568 21292
rect 4418 21184 4522 21230
rect 4418 21122 4568 21184
rect 4418 21076 4522 21122
rect 4418 21014 4568 21076
rect 4418 20968 4522 21014
rect 4418 20907 4568 20968
rect 4418 20861 4522 20907
rect 4418 20800 4568 20861
rect 4418 20754 4522 20800
rect 4418 20693 4568 20754
rect 4418 20647 4522 20693
rect 4418 20586 4568 20647
rect 4418 20540 4522 20586
rect 4418 20479 4568 20540
rect 4418 20433 4522 20479
rect 4418 20372 4568 20433
rect 4418 20326 4522 20372
rect 4418 20313 4568 20326
rect 4746 21662 4919 21675
rect 4792 21616 4919 21662
rect 4746 21554 4919 21616
rect 4792 21508 4919 21554
rect 4746 21446 4919 21508
rect 4792 21400 4919 21446
rect 4746 21338 4919 21400
rect 4792 21292 4919 21338
rect 4746 21230 4919 21292
rect 4792 21184 4919 21230
rect 4746 21122 4919 21184
rect 4792 21076 4919 21122
rect 4746 21014 4919 21076
rect 4792 20968 4919 21014
rect 4746 20907 4919 20968
rect 4792 20861 4919 20907
rect 4746 20800 4919 20861
rect 4792 20754 4919 20800
rect 4746 20693 4919 20754
rect 4792 20647 4919 20693
rect 4746 20586 4919 20647
rect 4792 20540 4919 20586
rect 4746 20479 4919 20540
rect 4792 20433 4919 20479
rect 4746 20372 4919 20433
rect 4792 20326 4919 20372
rect 4746 20313 4919 20326
rect 4418 19820 4488 20313
rect 4567 20229 4748 20243
rect 4567 20219 4634 20229
rect 4680 20219 4748 20229
rect 4567 20167 4629 20219
rect 4681 20167 4748 20219
rect 4567 20108 4748 20167
rect 4567 19955 4748 20028
rect 4567 19903 4631 19955
rect 4683 19903 4748 19955
rect 4567 19892 4748 19903
rect 4619 19891 4695 19892
rect 4826 19820 4919 20313
rect 4418 19807 4568 19820
rect 4418 19761 4522 19807
rect 4418 19699 4568 19761
rect 4418 19653 4522 19699
rect 4418 19591 4568 19653
rect 4418 19545 4522 19591
rect 4418 19483 4568 19545
rect 4418 19437 4522 19483
rect 4418 19375 4568 19437
rect 4418 19329 4522 19375
rect 4418 19267 4568 19329
rect 4418 19221 4522 19267
rect 4418 19159 4568 19221
rect 4418 19113 4522 19159
rect 4418 19052 4568 19113
rect 4418 19006 4522 19052
rect 4418 18945 4568 19006
rect 4418 18899 4522 18945
rect 4418 18838 4568 18899
rect 4418 18792 4522 18838
rect 4418 18731 4568 18792
rect 4418 18685 4522 18731
rect 4418 18624 4568 18685
rect 4418 18578 4522 18624
rect 4418 18517 4568 18578
rect 4418 18471 4522 18517
rect 4418 18470 4568 18471
rect 4746 19807 4919 19820
rect 4792 19761 4919 19807
rect 4746 19699 4919 19761
rect 4792 19653 4919 19699
rect 4746 19591 4919 19653
rect 4792 19545 4919 19591
rect 4746 19483 4919 19545
rect 4792 19437 4919 19483
rect 4746 19375 4919 19437
rect 4792 19329 4919 19375
rect 4746 19267 4919 19329
rect 4792 19221 4919 19267
rect 4746 19159 4919 19221
rect 4792 19113 4919 19159
rect 4746 19052 4919 19113
rect 4792 19006 4919 19052
rect 4746 18945 4919 19006
rect 4792 18899 4919 18945
rect 4746 18838 4919 18899
rect 4792 18792 4919 18838
rect 4746 18731 4919 18792
rect 4792 18685 4919 18731
rect 4746 18624 4919 18685
rect 4792 18578 4919 18624
rect 4746 18517 4919 18578
rect 4792 18471 4919 18517
rect 4418 18406 4603 18470
rect 4746 18468 4919 18471
rect 5015 21818 5528 21844
rect 5015 21766 5459 21818
rect 5511 21766 5528 21818
rect 5015 21747 5528 21766
rect 5015 21675 5155 21747
rect 5015 21662 5188 21675
rect 5015 21616 5142 21662
rect 5015 21554 5188 21616
rect 5015 21508 5142 21554
rect 5015 21446 5188 21508
rect 5015 21400 5142 21446
rect 5015 21338 5188 21400
rect 5015 21292 5142 21338
rect 5015 21230 5188 21292
rect 5015 21184 5142 21230
rect 5015 21122 5188 21184
rect 5015 21076 5142 21122
rect 5015 21014 5188 21076
rect 5015 20968 5142 21014
rect 5015 20907 5188 20968
rect 5015 20861 5142 20907
rect 5015 20800 5188 20861
rect 5015 20754 5142 20800
rect 5015 20693 5188 20754
rect 5015 20647 5142 20693
rect 5015 20586 5188 20647
rect 5015 20540 5142 20586
rect 5015 20479 5188 20540
rect 5015 20433 5142 20479
rect 5015 20372 5188 20433
rect 5015 20326 5142 20372
rect 5015 20313 5188 20326
rect 5366 21667 5412 21675
rect 5366 21662 5517 21667
rect 5412 21616 5517 21662
rect 5366 21554 5517 21616
rect 5412 21508 5517 21554
rect 5366 21446 5517 21508
rect 5412 21400 5517 21446
rect 5366 21338 5517 21400
rect 5412 21292 5517 21338
rect 5366 21230 5517 21292
rect 5412 21184 5517 21230
rect 5366 21122 5517 21184
rect 5412 21076 5517 21122
rect 5366 21014 5517 21076
rect 5412 20968 5517 21014
rect 5366 20907 5517 20968
rect 5412 20861 5517 20907
rect 5366 20800 5517 20861
rect 5412 20754 5517 20800
rect 5366 20693 5517 20754
rect 5412 20647 5517 20693
rect 5366 20586 5517 20647
rect 5412 20540 5517 20586
rect 5366 20479 5517 20540
rect 5412 20433 5517 20479
rect 5366 20372 5517 20433
rect 5412 20326 5517 20372
rect 5366 20313 5517 20326
rect 5015 19820 5112 20313
rect 5186 20229 5368 20243
rect 5186 20219 5254 20229
rect 5300 20219 5368 20229
rect 5186 20167 5253 20219
rect 5305 20167 5368 20219
rect 5186 20108 5368 20167
rect 5186 19956 5368 20028
rect 5186 19904 5251 19956
rect 5303 19904 5368 19956
rect 5186 19892 5368 19904
rect 5431 19820 5517 20313
rect 5015 19807 5188 19820
rect 5015 19761 5142 19807
rect 5015 19699 5188 19761
rect 5015 19653 5142 19699
rect 5015 19591 5188 19653
rect 5015 19545 5142 19591
rect 5015 19483 5188 19545
rect 5015 19437 5142 19483
rect 5015 19375 5188 19437
rect 5015 19329 5142 19375
rect 5015 19267 5188 19329
rect 5015 19221 5142 19267
rect 5015 19159 5188 19221
rect 5015 19113 5142 19159
rect 5015 19052 5188 19113
rect 5015 19006 5142 19052
rect 5015 18945 5188 19006
rect 5015 18899 5142 18945
rect 5015 18838 5188 18899
rect 5015 18792 5142 18838
rect 5015 18731 5188 18792
rect 5015 18685 5142 18731
rect 5015 18624 5188 18685
rect 5015 18578 5142 18624
rect 5015 18517 5188 18578
rect 5015 18471 5142 18517
rect 5015 18468 5188 18471
rect 4746 18458 4792 18468
rect 5142 18458 5188 18468
rect 5366 19807 5517 19820
rect 5412 19761 5517 19807
rect 5366 19699 5517 19761
rect 5412 19653 5517 19699
rect 5366 19591 5517 19653
rect 5412 19545 5517 19591
rect 5366 19483 5517 19545
rect 5412 19437 5517 19483
rect 5366 19375 5517 19437
rect 5412 19329 5517 19375
rect 5366 19267 5517 19329
rect 5412 19221 5517 19267
rect 5366 19159 5517 19221
rect 5412 19113 5517 19159
rect 5366 19052 5517 19113
rect 5412 19006 5517 19052
rect 5366 18945 5517 19006
rect 5412 18899 5517 18945
rect 5366 18838 5517 18899
rect 5412 18792 5517 18838
rect 5366 18731 5517 18792
rect 5412 18685 5517 18731
rect 5366 18624 5517 18685
rect 5412 18578 5517 18624
rect 5366 18517 5517 18578
rect 5412 18471 5517 18517
rect 5366 18458 5517 18471
rect 4092 18386 4603 18406
rect 4092 18334 4224 18386
rect 4276 18334 4410 18386
rect 4462 18334 4603 18386
rect 4092 18314 4603 18334
rect 5388 18378 5517 18458
rect 5388 18326 5453 18378
rect 5505 18326 5517 18378
rect 5388 18314 5517 18326
rect 631 18178 5587 18212
rect 631 18175 1699 18178
rect 631 18129 754 18175
rect 800 18129 912 18175
rect 958 18129 1070 18175
rect 1116 18129 1228 18175
rect 1274 18129 1386 18175
rect 1432 18129 1544 18175
rect 1590 18129 1699 18175
rect 631 18126 1699 18129
rect 1751 18126 1990 18178
rect 2042 18175 2938 18178
rect 2042 18129 2151 18175
rect 2197 18129 2309 18175
rect 2355 18129 2467 18175
rect 2513 18129 2625 18175
rect 2671 18129 2783 18175
rect 2829 18129 2938 18175
rect 2042 18126 2938 18129
rect 2990 18126 3229 18178
rect 3281 18175 4176 18178
rect 3281 18129 3389 18175
rect 3435 18129 3547 18175
rect 3593 18129 3705 18175
rect 3751 18129 3863 18175
rect 3909 18129 4021 18175
rect 4067 18129 4176 18175
rect 3281 18126 4176 18129
rect 4228 18126 4467 18178
rect 4519 18175 5587 18178
rect 4519 18129 4628 18175
rect 4674 18129 4786 18175
rect 4832 18129 4944 18175
rect 4990 18129 5102 18175
rect 5148 18129 5260 18175
rect 5306 18129 5418 18175
rect 5464 18129 5587 18175
rect 4519 18126 5587 18129
rect 631 18092 5587 18126
rect 631 17836 702 18092
rect 847 17987 1115 18012
rect 847 17935 913 17987
rect 965 17985 1115 17987
rect 965 17939 975 17985
rect 1021 17939 1115 17985
rect 965 17935 1115 17939
rect 847 17915 1115 17935
rect 631 17720 805 17836
rect 631 17674 725 17720
rect 771 17674 805 17720
rect 631 17557 805 17674
rect 948 17824 1056 17836
rect 948 17668 973 17824
rect 1025 17668 1056 17824
rect 510 17260 578 17263
rect 510 17252 826 17260
rect 510 17112 521 17252
rect 567 17223 826 17252
rect 567 17177 780 17223
rect 567 17112 826 17177
rect 948 17223 1056 17668
rect 1194 17720 1308 18092
rect 1387 17987 1655 18012
rect 1387 17985 1537 17987
rect 1387 17939 1481 17985
rect 1527 17939 1537 17985
rect 1387 17935 1537 17939
rect 1589 17935 1655 17987
rect 1387 17915 1655 17935
rect 1800 17836 1941 18092
rect 2086 17987 2354 18012
rect 2086 17935 2152 17987
rect 2204 17985 2354 17987
rect 2204 17939 2214 17985
rect 2260 17939 2354 17985
rect 2204 17935 2354 17939
rect 2086 17915 2354 17935
rect 1194 17674 1228 17720
rect 1274 17674 1308 17720
rect 1194 17557 1308 17674
rect 1446 17824 1554 17836
rect 1446 17668 1477 17824
rect 1529 17668 1554 17824
rect 948 17177 1004 17223
rect 1050 17177 1056 17223
rect 948 17140 1056 17177
rect 1194 17223 1308 17260
rect 1194 17177 1228 17223
rect 1274 17177 1308 17223
rect 510 17031 826 17112
rect 1194 17031 1308 17177
rect 1446 17223 1554 17668
rect 1697 17720 2044 17836
rect 1697 17674 1731 17720
rect 1777 17674 1964 17720
rect 2010 17674 2044 17720
rect 1697 17557 2044 17674
rect 2187 17824 2295 17836
rect 2187 17668 2212 17824
rect 2264 17668 2295 17824
rect 1837 17260 1905 17263
rect 1446 17177 1452 17223
rect 1498 17177 1554 17223
rect 1446 17140 1554 17177
rect 1676 17252 2065 17260
rect 1676 17223 1848 17252
rect 1722 17177 1848 17223
rect 1676 17112 1848 17177
rect 1894 17223 2065 17252
rect 1894 17177 2019 17223
rect 1894 17112 2065 17177
rect 2187 17223 2295 17668
rect 2433 17720 2547 18092
rect 2626 17987 2894 18012
rect 2626 17985 2776 17987
rect 2626 17939 2720 17985
rect 2766 17939 2776 17985
rect 2626 17935 2776 17939
rect 2828 17935 2894 17987
rect 2626 17915 2894 17935
rect 3039 17836 3179 18092
rect 3324 17987 3592 18012
rect 3324 17935 3390 17987
rect 3442 17985 3592 17987
rect 3442 17939 3452 17985
rect 3498 17939 3592 17985
rect 3442 17935 3592 17939
rect 3324 17915 3592 17935
rect 2433 17674 2467 17720
rect 2513 17674 2547 17720
rect 2433 17557 2547 17674
rect 2685 17824 2793 17836
rect 2685 17668 2716 17824
rect 2768 17668 2793 17824
rect 2187 17177 2243 17223
rect 2289 17177 2295 17223
rect 2187 17140 2295 17177
rect 2433 17223 2547 17260
rect 2433 17177 2467 17223
rect 2513 17177 2547 17223
rect 1676 17031 2065 17112
rect 2433 17031 2547 17177
rect 2685 17223 2793 17668
rect 2936 17720 3282 17836
rect 2936 17674 2970 17720
rect 3016 17674 3202 17720
rect 3248 17674 3282 17720
rect 2936 17557 3282 17674
rect 3425 17824 3533 17836
rect 3425 17668 3450 17824
rect 3502 17668 3533 17824
rect 3076 17260 3144 17263
rect 2685 17177 2691 17223
rect 2737 17177 2793 17223
rect 2685 17140 2793 17177
rect 2915 17252 3303 17260
rect 2915 17223 3087 17252
rect 2961 17177 3087 17223
rect 2915 17112 3087 17177
rect 3133 17223 3303 17252
rect 3133 17177 3257 17223
rect 3133 17112 3303 17177
rect 3425 17223 3533 17668
rect 3671 17720 3785 18092
rect 3864 17987 4132 18012
rect 3864 17985 4014 17987
rect 3864 17939 3958 17985
rect 4004 17939 4014 17985
rect 3864 17935 4014 17939
rect 4066 17935 4132 17987
rect 3864 17915 4132 17935
rect 4277 17836 4418 18092
rect 4563 17987 4831 18012
rect 4563 17935 4629 17987
rect 4681 17985 4831 17987
rect 4681 17939 4691 17985
rect 4737 17939 4831 17985
rect 4681 17935 4831 17939
rect 4563 17915 4831 17935
rect 3671 17674 3705 17720
rect 3751 17674 3785 17720
rect 3671 17557 3785 17674
rect 3923 17824 4031 17836
rect 3923 17668 3954 17824
rect 4006 17668 4031 17824
rect 3425 17177 3481 17223
rect 3527 17177 3533 17223
rect 3425 17140 3533 17177
rect 3671 17223 3785 17260
rect 3671 17177 3705 17223
rect 3751 17177 3785 17223
rect 2915 17031 3303 17112
rect 3671 17031 3785 17177
rect 3923 17223 4031 17668
rect 4174 17720 4521 17836
rect 4174 17674 4208 17720
rect 4254 17674 4441 17720
rect 4487 17674 4521 17720
rect 4174 17557 4521 17674
rect 4664 17824 4772 17836
rect 4664 17668 4689 17824
rect 4741 17668 4772 17824
rect 4314 17260 4382 17263
rect 3923 17177 3929 17223
rect 3975 17177 4031 17223
rect 3923 17140 4031 17177
rect 4153 17252 4542 17260
rect 4153 17223 4325 17252
rect 4199 17177 4325 17223
rect 4153 17112 4325 17177
rect 4371 17223 4542 17252
rect 4371 17177 4496 17223
rect 4371 17112 4542 17177
rect 4664 17223 4772 17668
rect 4909 17720 5025 18092
rect 5103 17988 5372 18012
rect 5103 17985 5254 17988
rect 5103 17939 5197 17985
rect 5243 17939 5254 17985
rect 5103 17936 5254 17939
rect 5306 17936 5372 17988
rect 5103 17915 5372 17936
rect 5515 17836 5587 18092
rect 4909 17674 4944 17720
rect 4990 17674 5025 17720
rect 4909 17557 5025 17674
rect 5162 17824 5291 17836
rect 5162 17668 5174 17824
rect 5226 17720 5291 17824
rect 5243 17674 5291 17720
rect 5226 17668 5291 17674
rect 5162 17557 5291 17668
rect 5412 17720 5587 17836
rect 5412 17674 5447 17720
rect 5493 17674 5587 17720
rect 5412 17557 5587 17674
rect 5184 17260 5256 17557
rect 5553 17260 5621 17263
rect 4664 17177 4720 17223
rect 4766 17177 4772 17223
rect 4664 17140 4772 17177
rect 4909 17223 5025 17260
rect 4909 17177 4944 17223
rect 4990 17177 5025 17223
rect 4153 17031 4542 17112
rect 4909 17031 5025 17177
rect 5159 17223 5256 17260
rect 5159 17177 5168 17223
rect 5214 17177 5256 17223
rect 5159 17140 5256 17177
rect 5392 17252 5621 17260
rect 5392 17223 5564 17252
rect 5438 17177 5564 17223
rect 5392 17112 5564 17177
rect 5610 17112 5621 17252
rect 5392 17101 5621 17112
rect 5392 17031 5587 17101
rect 510 16940 5587 17031
rect 510 16888 915 16940
rect 967 16888 1535 16940
rect 1587 16888 2154 16940
rect 2206 16888 2774 16940
rect 2826 16888 3392 16940
rect 3444 16888 4012 16940
rect 4064 16888 4631 16940
rect 4683 16888 5251 16940
rect 5303 16888 5587 16940
rect 510 16856 5587 16888
rect 510 16810 754 16856
rect 800 16810 912 16856
rect 958 16810 1070 16856
rect 1116 16810 1228 16856
rect 1274 16810 1386 16856
rect 1432 16810 1544 16856
rect 1590 16810 1702 16856
rect 1748 16810 1993 16856
rect 2039 16810 2151 16856
rect 2197 16810 2309 16856
rect 2355 16810 2467 16856
rect 2513 16810 2625 16856
rect 2671 16810 2783 16856
rect 2829 16810 2941 16856
rect 2987 16810 3231 16856
rect 3277 16810 3389 16856
rect 3435 16810 3547 16856
rect 3593 16810 3705 16856
rect 3751 16810 3863 16856
rect 3909 16810 4021 16856
rect 4067 16810 4179 16856
rect 4225 16810 4470 16856
rect 4516 16810 4628 16856
rect 4674 16810 4786 16856
rect 4832 16810 4944 16856
rect 4990 16810 5102 16856
rect 5148 16810 5260 16856
rect 5306 16810 5418 16856
rect 5464 16810 5587 16856
rect 510 16759 5587 16810
rect 678 16623 2390 16648
rect 678 16571 728 16623
rect 780 16571 914 16623
rect 966 16571 1745 16623
rect 1797 16571 1931 16623
rect 1983 16571 2390 16623
rect 678 16551 2390 16571
rect 678 16435 2390 16439
rect 678 16415 2624 16435
rect 678 16363 1108 16415
rect 1160 16363 1294 16415
rect 1346 16363 2346 16415
rect 2398 16363 2532 16415
rect 2584 16363 2624 16415
rect 678 16343 2624 16363
rect 4824 16415 5132 16435
rect 4824 16363 4854 16415
rect 4906 16363 5040 16415
rect 5092 16363 5132 16415
rect 4824 16343 5132 16363
rect 678 16342 2390 16343
rect 929 16230 1058 16231
rect 368 16190 3328 16230
rect 368 16138 967 16190
rect 1019 16138 1761 16190
rect 1813 16138 1972 16190
rect 2024 16138 2182 16190
rect 2234 16138 2393 16190
rect 2445 16138 2605 16190
rect 2657 16138 2816 16190
rect 2868 16138 3026 16190
rect 3078 16138 3237 16190
rect 3289 16138 3328 16190
rect 368 16097 3328 16138
rect 3675 16190 4437 16230
rect 3675 16138 3713 16190
rect 3765 16138 3924 16190
rect 3976 16138 4136 16190
rect 4188 16138 4347 16190
rect 4399 16138 4437 16190
rect 3675 16097 4437 16138
rect 368 16093 2390 16097
rect 487 15953 1903 15976
rect 487 15901 499 15953
rect 551 15901 1903 15953
rect 487 15880 1903 15901
rect 2258 15936 2350 15977
rect 2258 15884 2278 15936
rect 2330 15884 2350 15936
rect 913 15781 1413 15782
rect 300 15765 346 15778
rect 277 15612 300 15642
rect 524 15765 570 15778
rect 346 15612 369 15642
rect 277 15560 297 15612
rect 349 15560 369 15612
rect 277 15426 300 15560
rect 346 15426 369 15560
rect 277 15374 297 15426
rect 349 15374 369 15426
rect 277 15334 300 15374
rect 277 15013 300 15043
rect 346 15334 369 15374
rect 346 15013 369 15043
rect 277 14961 297 15013
rect 349 14961 369 15013
rect 277 14827 300 14961
rect 346 14827 369 14961
rect 277 14775 297 14827
rect 349 14775 369 14827
rect 277 14735 300 14775
rect 277 13556 300 13586
rect 346 14735 369 14775
rect 346 13556 369 13586
rect 277 13504 297 13556
rect 349 13504 369 13556
rect 277 13370 300 13504
rect 346 13370 369 13504
rect 277 13318 297 13370
rect 349 13318 369 13370
rect 277 13278 300 13318
rect 346 13278 369 13318
rect 300 13056 346 13069
rect 489 13069 524 13331
rect 913 15741 1491 15781
rect 913 15707 1419 15741
rect 913 15591 1009 15707
rect 1399 15689 1419 15707
rect 1471 15689 1491 15741
rect 913 15545 948 15591
rect 994 15545 1009 15591
rect 913 15485 1009 15545
rect 1126 15591 1292 15627
rect 1126 15545 1211 15591
rect 1257 15545 1292 15591
rect 1126 15508 1292 15545
rect 1399 15555 1491 15689
rect 2258 15750 2350 15884
rect 2258 15698 2278 15750
rect 2330 15698 2350 15750
rect 2258 15658 2350 15698
rect 790 15368 1048 15405
rect 790 15365 990 15368
rect 790 15313 967 15365
rect 1036 15322 1048 15368
rect 1019 15313 1048 15322
rect 790 15272 1048 15313
rect 1126 15188 1198 15508
rect 1399 15503 1419 15555
rect 1471 15503 1491 15555
rect 1399 15462 1491 15503
rect 1627 15565 1935 15585
rect 1627 15513 1657 15565
rect 1709 15562 1843 15565
rect 1895 15562 1935 15565
rect 1899 15516 1935 15562
rect 1709 15513 1843 15516
rect 1895 15513 1935 15516
rect 1627 15493 1935 15513
rect 2318 15509 2478 15559
rect 1644 15311 1690 15324
rect 1644 15207 1690 15265
rect 818 15072 915 15176
rect 818 15026 853 15072
rect 899 15026 915 15072
rect 818 14909 915 15026
rect 1082 15072 1198 15188
rect 1082 15026 1117 15072
rect 1163 15026 1198 15072
rect 1082 14909 1198 15026
rect 842 14562 915 14909
rect 1126 14716 1198 14909
rect 1074 14702 1198 14716
rect 1074 14656 1108 14702
rect 1154 14656 1198 14702
rect 1074 14642 1198 14656
rect 1315 15177 1431 15188
rect 1315 15147 1449 15177
rect 1315 15095 1377 15147
rect 1429 15095 1449 15147
rect 1315 15072 1449 15095
rect 1315 15026 1350 15072
rect 1396 15026 1449 15072
rect 1315 14961 1449 15026
rect 1315 14909 1377 14961
rect 1429 14909 1449 14961
rect 1315 14869 1449 14909
rect 1644 15103 1690 15161
rect 1868 15311 1914 15493
rect 1868 15207 1914 15265
rect 1868 15103 1914 15161
rect 1644 14999 1690 15057
rect 1644 14895 1690 14953
rect 1315 14562 1387 14869
rect 842 14488 1387 14562
rect 1644 14791 1690 14849
rect 1847 15057 1868 15077
rect 2318 15463 2366 15509
rect 2412 15463 2478 15509
rect 2318 15345 2478 15463
rect 2318 15299 2366 15345
rect 2412 15299 2478 15345
rect 2318 15182 2478 15299
rect 2318 15136 2366 15182
rect 2412 15136 2478 15182
rect 1914 15057 1939 15077
rect 1847 15047 1939 15057
rect 1847 14995 1867 15047
rect 1919 14995 1939 15047
rect 1847 14953 1868 14995
rect 1914 14953 1939 14995
rect 1847 14895 1939 14953
rect 1847 14861 1868 14895
rect 1914 14861 1939 14895
rect 1847 14809 1867 14861
rect 1919 14809 1939 14861
rect 1847 14791 1939 14809
rect 1847 14769 1868 14791
rect 1644 14687 1690 14745
rect 1644 14583 1690 14641
rect 1644 14479 1690 14537
rect 748 14405 794 14418
rect 720 14359 748 14398
rect 972 14405 1018 14418
rect 794 14359 812 14398
rect 720 14358 812 14359
rect 720 14306 740 14358
rect 792 14306 812 14358
rect 720 14298 812 14306
rect 720 14252 748 14298
rect 794 14252 812 14298
rect 720 14191 812 14252
rect 720 14172 748 14191
rect 720 14120 740 14172
rect 794 14145 812 14191
rect 792 14120 812 14145
rect 720 14084 812 14120
rect 720 14079 748 14084
rect 794 14079 812 14084
rect 1196 14405 1242 14418
rect 972 14298 1018 14359
rect 972 14191 1018 14252
rect 972 14084 1018 14145
rect 748 13977 794 14038
rect 748 13870 794 13931
rect 748 13763 794 13824
rect 748 13655 794 13717
rect 748 13547 794 13609
rect 748 13439 794 13501
rect 748 13331 794 13393
rect 1173 14359 1196 14398
rect 1420 14405 1466 14418
rect 1242 14359 1265 14398
rect 1173 14358 1265 14359
rect 1173 14306 1193 14358
rect 1245 14306 1265 14358
rect 1173 14298 1265 14306
rect 1173 14252 1196 14298
rect 1242 14252 1265 14298
rect 1173 14191 1265 14252
rect 1173 14172 1196 14191
rect 1242 14172 1265 14191
rect 1173 14120 1193 14172
rect 1245 14120 1265 14172
rect 1173 14084 1265 14120
rect 1173 14079 1196 14084
rect 972 13977 1018 14038
rect 972 13870 1018 13931
rect 972 13763 1018 13824
rect 972 13655 1018 13717
rect 972 13547 1018 13609
rect 972 13439 1018 13501
rect 972 13331 1018 13393
rect 1242 14079 1265 14084
rect 1420 14298 1466 14359
rect 1420 14191 1466 14252
rect 1420 14084 1466 14145
rect 1196 13977 1242 14038
rect 1196 13870 1242 13931
rect 1196 13763 1242 13824
rect 1196 13655 1242 13717
rect 1196 13547 1242 13609
rect 1196 13439 1242 13501
rect 1196 13331 1242 13393
rect 570 13069 605 13331
rect 489 12896 605 13069
rect 748 13223 794 13285
rect 748 13115 794 13177
rect 748 13056 794 13069
rect 937 13285 972 13331
rect 1018 13285 1053 13331
rect 937 13223 1053 13285
rect 937 13177 972 13223
rect 1018 13177 1053 13223
rect 937 13115 1053 13177
rect 937 13069 972 13115
rect 1018 13069 1053 13115
rect 937 12896 1053 13069
rect 1196 13223 1242 13285
rect 1420 13977 1466 14038
rect 1420 13870 1466 13931
rect 1420 13763 1466 13824
rect 1420 13655 1466 13717
rect 1420 13547 1466 13609
rect 1420 13439 1466 13501
rect 1420 13331 1466 13393
rect 1420 13223 1466 13285
rect 1196 13115 1242 13177
rect 1196 13056 1242 13069
rect 1385 13177 1420 13184
rect 1644 14375 1690 14433
rect 1644 14270 1690 14329
rect 1644 14165 1690 14224
rect 1644 14060 1690 14119
rect 1644 13955 1690 14014
rect 1644 13850 1690 13909
rect 1644 13745 1690 13804
rect 1644 13640 1690 13699
rect 1644 13535 1690 13594
rect 1914 14769 1939 14791
rect 2318 15019 2478 15136
rect 2318 14973 2366 15019
rect 2412 14973 2478 15019
rect 2318 14856 2478 14973
rect 2318 14810 2366 14856
rect 2412 14810 2478 14856
rect 1868 14687 1914 14745
rect 1868 14583 1914 14641
rect 1868 14479 1914 14537
rect 1868 14375 1914 14433
rect 1868 14270 1914 14329
rect 1868 14165 1914 14224
rect 1868 14060 1914 14119
rect 1868 13955 1914 14014
rect 1868 13850 1914 13909
rect 1868 13745 1914 13804
rect 1868 13640 1914 13699
rect 1868 13586 1914 13594
rect 2318 14693 2478 14810
rect 2318 14647 2366 14693
rect 2412 14647 2478 14693
rect 2318 14529 2478 14647
rect 2318 14483 2366 14529
rect 2412 14483 2478 14529
rect 2318 14366 2478 14483
rect 2318 14320 2366 14366
rect 2412 14320 2478 14366
rect 2318 14203 2478 14320
rect 2318 14157 2366 14203
rect 2412 14157 2478 14203
rect 2318 14040 2478 14157
rect 2318 13994 2366 14040
rect 2412 13994 2478 14040
rect 2318 13876 2478 13994
rect 2318 13830 2366 13876
rect 2412 13830 2478 13876
rect 2318 13713 2478 13830
rect 2318 13667 2366 13713
rect 2412 13667 2478 13713
rect 1644 13430 1690 13489
rect 1644 13331 1690 13384
rect 1847 13556 1939 13586
rect 1847 13504 1867 13556
rect 1919 13504 1939 13556
rect 1847 13489 1868 13504
rect 1914 13489 1939 13504
rect 1847 13430 1939 13489
rect 1847 13384 1868 13430
rect 1914 13384 1939 13430
rect 1847 13370 1939 13384
rect 1644 13325 1725 13331
rect 1690 13279 1725 13325
rect 1644 13220 1725 13279
rect 1847 13318 1867 13370
rect 1919 13318 1939 13370
rect 1847 13279 1868 13318
rect 1914 13279 1939 13318
rect 1847 13278 1939 13279
rect 2318 13550 2478 13667
rect 2318 13504 2366 13550
rect 2412 13504 2478 13550
rect 2318 13387 2478 13504
rect 2318 13341 2366 13387
rect 2412 13341 2478 13387
rect 1466 13177 1644 13184
rect 1385 13174 1644 13177
rect 1690 13174 1725 13220
rect 1385 13115 1725 13174
rect 1385 13069 1420 13115
rect 1466 13069 1644 13115
rect 1690 13069 1725 13115
rect 1385 13064 1725 13069
rect 1420 13056 1466 13064
rect 1644 13056 1725 13064
rect 1868 13220 1914 13278
rect 1868 13115 1914 13174
rect 1868 13056 1914 13069
rect 2318 13223 2478 13341
rect 2318 13177 2366 13223
rect 2412 13177 2478 13223
rect 2318 13060 2478 13177
rect 489 12859 1576 12896
rect 489 12813 1516 12859
rect 1562 12813 1576 12859
rect 489 12776 1576 12813
rect 300 12607 346 12620
rect 277 12561 300 12591
rect 489 12607 605 12776
rect 748 12607 794 12619
rect 346 12561 369 12591
rect 277 12509 297 12561
rect 349 12509 369 12561
rect 489 12520 524 12607
rect 277 12375 300 12509
rect 346 12375 369 12509
rect 277 12323 297 12375
rect 349 12323 369 12375
rect 277 12283 300 12323
rect 277 11613 300 11643
rect 346 12283 369 12323
rect 346 11613 369 11643
rect 277 11561 297 11613
rect 349 11561 369 11613
rect 277 11427 300 11561
rect 346 11427 369 11561
rect 277 11375 297 11427
rect 349 11375 369 11427
rect 277 11335 300 11375
rect 277 10697 300 10727
rect 346 11335 369 11375
rect 346 10697 369 10727
rect 277 10645 297 10697
rect 349 10645 369 10697
rect 277 10511 300 10645
rect 346 10511 369 10645
rect 277 10459 297 10511
rect 349 10459 369 10511
rect 277 10419 300 10459
rect 346 10419 369 10459
rect 300 9898 346 9911
rect 570 12520 605 12607
rect 723 12606 815 12607
rect 723 12567 748 12606
rect 794 12567 815 12606
rect 723 12515 743 12567
rect 795 12515 815 12567
rect 937 12606 1053 12776
rect 1653 12619 1725 13056
rect 2318 13014 2366 13060
rect 2412 13014 2478 13060
rect 2318 12897 2478 13014
rect 2318 12851 2366 12897
rect 2412 12851 2478 12897
rect 2318 12733 2478 12851
rect 2318 12687 2366 12733
rect 2412 12687 2478 12733
rect 2073 12629 2165 12659
rect 2073 12621 2093 12629
rect 1196 12607 1242 12619
rect 1420 12610 1466 12619
rect 1644 12610 1725 12619
rect 937 12560 972 12606
rect 1018 12560 1053 12606
rect 937 12520 1053 12560
rect 1173 12606 1265 12607
rect 1173 12567 1196 12606
rect 1242 12567 1265 12606
rect 723 12502 815 12515
rect 723 12456 748 12502
rect 794 12456 815 12502
rect 723 12398 815 12456
rect 723 12381 748 12398
rect 794 12381 815 12398
rect 723 12329 743 12381
rect 795 12329 815 12381
rect 723 12294 815 12329
rect 723 12288 748 12294
rect 794 12288 815 12294
rect 972 12502 1018 12520
rect 972 12398 1018 12456
rect 972 12294 1018 12352
rect 748 12190 794 12248
rect 748 12086 794 12144
rect 748 11982 794 12040
rect 748 11878 794 11936
rect 748 11774 794 11832
rect 748 11670 794 11728
rect 748 11565 794 11624
rect 748 11460 794 11519
rect 748 11355 794 11414
rect 748 11250 794 11309
rect 748 11145 794 11204
rect 748 11040 794 11099
rect 748 10935 794 10994
rect 748 10830 794 10889
rect 748 10725 794 10784
rect 748 10620 794 10679
rect 748 10515 794 10574
rect 748 10410 794 10469
rect 748 10351 794 10364
rect 1173 12515 1193 12567
rect 1245 12515 1265 12567
rect 1173 12502 1265 12515
rect 1173 12456 1196 12502
rect 1242 12456 1265 12502
rect 1385 12606 1725 12610
rect 1385 12560 1420 12606
rect 1466 12560 1644 12606
rect 1690 12560 1725 12606
rect 1385 12502 1725 12560
rect 1385 12490 1420 12502
rect 1173 12398 1265 12456
rect 1173 12381 1196 12398
rect 1242 12381 1265 12398
rect 1173 12329 1193 12381
rect 1245 12329 1265 12381
rect 1173 12294 1265 12329
rect 1173 12288 1196 12294
rect 972 12190 1018 12248
rect 972 12086 1018 12144
rect 972 11982 1018 12040
rect 972 11878 1018 11936
rect 972 11774 1018 11832
rect 972 11670 1018 11728
rect 972 11565 1018 11624
rect 972 11460 1018 11519
rect 972 11355 1018 11414
rect 972 11250 1018 11309
rect 972 11145 1018 11204
rect 972 11040 1018 11099
rect 972 10935 1018 10994
rect 972 10830 1018 10889
rect 972 10725 1018 10784
rect 972 10620 1018 10679
rect 972 10515 1018 10574
rect 972 10410 1018 10469
rect 972 10351 1018 10364
rect 1242 12288 1265 12294
rect 1466 12490 1644 12502
rect 1420 12398 1466 12456
rect 1420 12294 1466 12352
rect 1196 12190 1242 12248
rect 1196 12086 1242 12144
rect 1196 11982 1242 12040
rect 1196 11878 1242 11936
rect 1196 11774 1242 11832
rect 1196 11670 1242 11728
rect 1196 11565 1242 11624
rect 1196 11460 1242 11519
rect 1196 11355 1242 11414
rect 1196 11250 1242 11309
rect 1196 11145 1242 11204
rect 1196 11040 1242 11099
rect 1196 10935 1242 10994
rect 1196 10830 1242 10889
rect 1196 10725 1242 10784
rect 1196 10620 1242 10679
rect 1196 10515 1242 10574
rect 1196 10410 1242 10469
rect 1196 10351 1242 10364
rect 1420 12190 1466 12248
rect 1420 12086 1466 12144
rect 1420 11982 1466 12040
rect 1420 11878 1466 11936
rect 1420 11774 1466 11832
rect 1420 11670 1466 11728
rect 1420 11565 1466 11624
rect 1420 11460 1466 11519
rect 1420 11355 1466 11414
rect 1420 11250 1466 11309
rect 1420 11145 1466 11204
rect 1420 11040 1466 11099
rect 1420 10935 1466 10994
rect 1420 10830 1466 10889
rect 1420 10725 1466 10784
rect 1420 10620 1466 10679
rect 1420 10515 1466 10574
rect 1420 10410 1466 10469
rect 1420 10351 1466 10364
rect 1690 12490 1725 12502
rect 1833 12606 2093 12621
rect 1833 12561 1868 12606
rect 1914 12577 2093 12606
rect 2145 12621 2165 12629
rect 2318 12621 2478 12687
rect 2145 12577 2478 12621
rect 1914 12571 2478 12577
rect 1833 12509 1854 12561
rect 1914 12560 2208 12571
rect 1906 12525 2208 12560
rect 2254 12570 2478 12571
rect 2254 12525 2366 12570
rect 1906 12524 2366 12525
rect 2412 12524 2478 12570
rect 1906 12509 2478 12524
rect 1833 12502 2478 12509
rect 1644 12398 1690 12456
rect 1644 12294 1690 12352
rect 1644 12190 1690 12248
rect 1644 12086 1690 12144
rect 1644 11982 1690 12040
rect 1644 11878 1690 11936
rect 1644 11774 1690 11832
rect 1644 11670 1690 11728
rect 1644 11565 1690 11624
rect 1644 11460 1690 11519
rect 1644 11355 1690 11414
rect 1644 11250 1690 11309
rect 1644 11145 1690 11204
rect 1644 11040 1690 11099
rect 1644 10935 1690 10994
rect 1644 10830 1690 10889
rect 1644 10725 1690 10784
rect 1644 10620 1690 10679
rect 1644 10515 1690 10574
rect 1644 10410 1690 10469
rect 1833 12456 1868 12502
rect 1914 12456 2478 12502
rect 1833 12443 2478 12456
rect 1833 12398 2093 12443
rect 1833 12375 1868 12398
rect 1914 12391 2093 12398
rect 2145 12407 2478 12443
rect 2145 12391 2208 12407
rect 1833 12323 1854 12375
rect 1914 12361 2208 12391
rect 2254 12361 2366 12407
rect 2412 12361 2478 12407
rect 1914 12352 2478 12361
rect 1906 12323 2478 12352
rect 1833 12294 2478 12323
rect 1833 12248 1868 12294
rect 1914 12248 2478 12294
rect 1833 12244 2478 12248
rect 1833 12198 2208 12244
rect 2254 12198 2366 12244
rect 2412 12198 2478 12244
rect 1833 12190 2478 12198
rect 1833 12144 1868 12190
rect 1914 12144 2478 12190
rect 1833 12086 2478 12144
rect 1833 12040 1868 12086
rect 1914 12081 2478 12086
rect 1914 12040 2208 12081
rect 1833 12035 2208 12040
rect 2254 12080 2478 12081
rect 2254 12035 2366 12080
rect 1833 12034 2366 12035
rect 2412 12034 2478 12080
rect 1833 11982 2478 12034
rect 1833 11936 1868 11982
rect 1914 11936 2478 11982
rect 1833 11918 2478 11936
rect 1833 11878 2208 11918
rect 1833 11832 1868 11878
rect 1914 11872 2208 11878
rect 2254 11917 2478 11918
rect 2254 11872 2366 11917
rect 1914 11871 2366 11872
rect 2412 11871 2478 11917
rect 1914 11853 2478 11871
rect 1914 11832 2093 11853
rect 1833 11801 2093 11832
rect 2145 11801 2478 11853
rect 1833 11774 2478 11801
rect 1833 11728 1868 11774
rect 1914 11754 2478 11774
rect 1914 11728 2208 11754
rect 1833 11708 2208 11728
rect 2254 11708 2366 11754
rect 2412 11708 2478 11754
rect 1833 11670 2478 11708
rect 1833 11624 1868 11670
rect 1914 11667 2478 11670
rect 1914 11624 2093 11667
rect 1833 11615 2093 11624
rect 2145 11615 2478 11667
rect 1833 11613 2478 11615
rect 1833 11561 1854 11613
rect 1906 11591 2478 11613
rect 1906 11565 2208 11591
rect 1833 11519 1868 11561
rect 1914 11545 2208 11565
rect 2254 11545 2366 11591
rect 2412 11545 2478 11591
rect 1914 11519 2478 11545
rect 1833 11460 2478 11519
rect 1833 11427 1868 11460
rect 1914 11428 2478 11460
rect 1833 11375 1854 11427
rect 1914 11414 2208 11428
rect 1906 11382 2208 11414
rect 2254 11427 2478 11428
rect 2254 11382 2366 11427
rect 1906 11381 2366 11382
rect 2412 11381 2478 11427
rect 1906 11375 2478 11381
rect 1833 11355 2478 11375
rect 1833 11309 1868 11355
rect 1914 11309 2478 11355
rect 1833 11264 2478 11309
rect 1833 11250 2208 11264
rect 1833 11204 1868 11250
rect 1914 11218 2208 11250
rect 2254 11218 2366 11264
rect 2412 11218 2478 11264
rect 1914 11204 2478 11218
rect 1833 11145 2478 11204
rect 1833 11099 1868 11145
rect 1914 11101 2478 11145
rect 1914 11099 2208 11101
rect 1833 11055 2208 11099
rect 2254 11055 2366 11101
rect 2412 11055 2478 11101
rect 1833 11040 2478 11055
rect 1833 10994 1868 11040
rect 1914 10994 2478 11040
rect 1833 10938 2478 10994
rect 1833 10937 2208 10938
rect 1833 10935 2093 10937
rect 1833 10889 1868 10935
rect 1914 10889 2093 10935
rect 1833 10885 2093 10889
rect 2145 10892 2208 10937
rect 2254 10892 2366 10938
rect 2412 10892 2478 10938
rect 2145 10885 2478 10892
rect 1833 10830 2478 10885
rect 1833 10784 1868 10830
rect 1914 10784 2478 10830
rect 1833 10775 2478 10784
rect 1833 10751 2208 10775
rect 1833 10725 2093 10751
rect 1833 10697 1868 10725
rect 1914 10699 2093 10725
rect 2145 10729 2208 10751
rect 2254 10729 2366 10775
rect 2412 10729 2478 10775
rect 2145 10699 2478 10729
rect 1833 10645 1854 10697
rect 1914 10679 2478 10699
rect 1906 10645 2478 10679
rect 1833 10620 2478 10645
rect 1833 10574 1868 10620
rect 1914 10611 2478 10620
rect 1914 10574 2208 10611
rect 1833 10565 2208 10574
rect 2254 10565 2366 10611
rect 2412 10565 2478 10611
rect 1833 10515 2478 10565
rect 1833 10511 1868 10515
rect 1833 10459 1854 10511
rect 1914 10469 2478 10515
rect 1906 10459 2478 10469
rect 1833 10410 2478 10459
rect 1833 10409 1868 10410
rect 1644 10351 1690 10364
rect 1914 10409 2478 10410
rect 1868 10351 1914 10364
rect 941 10265 1229 10279
rect 941 10219 976 10265
rect 1022 10255 1229 10265
rect 941 10203 978 10219
rect 1030 10203 1229 10255
rect 941 10183 1229 10203
rect 5344 10246 5438 11053
rect 5344 10194 5365 10246
rect 5417 10194 5438 10246
rect 524 9898 570 9911
rect 682 10052 2527 10103
rect 5344 10076 5438 10194
rect 682 10006 1741 10052
rect 1787 10006 2527 10052
rect 682 9984 2527 10006
rect 5345 10060 5437 10076
rect 5345 10008 5365 10060
rect 5417 10008 5437 10060
rect 682 9983 2481 9984
rect 682 9797 798 9983
rect 1629 9898 1675 9911
rect 377 9780 798 9797
rect 377 9734 412 9780
rect 458 9734 798 9780
rect 377 9677 798 9734
rect 898 9845 990 9875
rect 898 9798 918 9845
rect 898 9752 911 9798
rect 970 9793 990 9845
rect 1616 9852 1629 9875
rect 1853 9898 1899 9911
rect 1675 9852 1708 9875
rect 1616 9845 1708 9852
rect 957 9752 990 9793
rect 898 9678 990 9752
rect 898 9632 911 9678
rect 957 9659 990 9678
rect 898 9607 918 9632
rect 970 9607 990 9659
rect 1135 9803 1181 9811
rect 1135 9798 1220 9803
rect 1181 9752 1220 9798
rect 1135 9678 1220 9752
rect 1181 9632 1220 9678
rect 1135 9619 1220 9632
rect 252 9566 394 9577
rect 898 9567 990 9607
rect 252 9526 598 9566
rect 252 9525 300 9526
rect 346 9525 598 9526
rect 252 9473 296 9525
rect 348 9473 508 9525
rect 560 9473 598 9525
rect 252 9432 598 9473
rect 252 9429 394 9432
rect 1148 9420 1220 9619
rect 1616 9793 1636 9845
rect 1688 9793 1708 9845
rect 1616 9778 1708 9793
rect 1616 9732 1629 9778
rect 1675 9732 1708 9778
rect 1853 9778 1899 9852
rect 1616 9659 1708 9732
rect 1616 9607 1636 9659
rect 1688 9607 1708 9659
rect 1616 9567 1708 9607
rect 1817 9732 1853 9756
rect 2481 9856 2527 9938
rect 1899 9732 1933 9756
rect 1629 9427 1675 9440
rect 1018 9346 1503 9420
rect 801 9234 847 9247
rect 801 9124 847 9188
rect 1018 9234 1090 9346
rect 1018 9188 1025 9234
rect 1071 9188 1090 9234
rect 573 9104 881 9124
rect 573 9052 603 9104
rect 655 9052 789 9104
rect 841 9078 881 9104
rect 573 9032 801 9052
rect 847 9032 881 9078
rect 1018 9078 1090 9188
rect 1249 9234 1295 9247
rect 1249 9127 1295 9188
rect 1018 9032 1025 9078
rect 1071 9032 1090 9078
rect 801 9019 847 9032
rect 1018 9029 1090 9032
rect 1221 9087 1313 9127
rect 1221 9035 1241 9087
rect 1293 9078 1313 9087
rect 1221 9032 1249 9035
rect 1295 9032 1313 9078
rect 1025 9019 1071 9029
rect 277 9015 369 9018
rect 265 8988 381 9015
rect 265 8936 297 8988
rect 349 8936 381 8988
rect 265 8932 300 8936
rect 346 8932 381 8936
rect 265 8814 381 8932
rect 265 8802 300 8814
rect 346 8802 381 8814
rect 265 8750 297 8802
rect 349 8750 381 8802
rect 550 8887 956 8906
rect 550 8870 875 8887
rect 550 8818 647 8870
rect 699 8818 833 8870
rect 921 8841 956 8887
rect 885 8818 956 8841
rect 1221 8901 1313 9032
rect 1221 8849 1241 8901
rect 1293 8849 1313 8901
rect 1221 8819 1313 8849
rect 1431 9027 1503 9346
rect 1629 9271 1675 9381
rect 1431 8981 1444 9027
rect 1490 8981 1503 9027
rect 1593 9225 1629 9239
rect 1817 9427 1933 9732
rect 2481 9729 2527 9810
rect 2481 9602 2527 9683
rect 1817 9381 1853 9427
rect 1899 9381 1933 9427
rect 1817 9271 1933 9381
rect 2077 9427 2123 9440
rect 2077 9314 2123 9381
rect 1675 9225 1709 9239
rect 1593 9087 1709 9225
rect 1593 9035 1630 9087
rect 1682 9035 1709 9087
rect 1593 8995 1709 9035
rect 1817 9225 1853 9271
rect 1899 9225 1933 9271
rect 2043 9273 2135 9314
rect 2043 9239 2063 9273
rect 2115 9271 2135 9273
rect 1609 8994 1703 8995
rect 550 8797 956 8818
rect 265 8732 381 8750
rect 1039 8738 1131 8778
rect 276 8731 370 8732
rect 277 8710 369 8731
rect 1039 8686 1059 8738
rect 1111 8686 1131 8738
rect 1039 8643 1131 8686
rect 801 8630 847 8643
rect 461 8530 553 8570
rect 461 8478 481 8530
rect 533 8478 553 8530
rect 461 8371 553 8478
rect 801 8527 847 8584
rect 1025 8630 1131 8643
rect 1071 8584 1131 8630
rect 1025 8552 1131 8584
rect 801 8510 882 8527
rect 847 8464 882 8510
rect 801 8451 882 8464
rect 1025 8510 1059 8552
rect 1111 8500 1131 8552
rect 1071 8470 1131 8500
rect 1249 8630 1347 8643
rect 1295 8584 1347 8630
rect 1249 8510 1347 8584
rect 1025 8451 1071 8464
rect 1295 8464 1347 8510
rect 1249 8451 1347 8464
rect 461 8344 732 8371
rect 461 8292 481 8344
rect 533 8334 732 8344
rect 533 8292 673 8334
rect 461 8288 673 8292
rect 719 8288 732 8334
rect 461 8251 732 8288
rect 810 8348 882 8451
rect 810 8334 1197 8348
rect 810 8288 1117 8334
rect 1163 8288 1197 8334
rect 810 8274 1197 8288
rect 810 8170 882 8274
rect 1275 8170 1347 8451
rect 1431 8259 1503 8981
rect 1610 8901 1702 8994
rect 1610 8849 1630 8901
rect 1682 8849 1702 8901
rect 1610 8819 1702 8849
rect 1817 8915 1933 9225
rect 2041 9221 2063 9239
rect 2123 9239 2135 9271
rect 2481 9252 2527 9556
rect 2705 9984 2751 9997
rect 2751 9940 2864 9970
rect 5345 9967 5437 10008
rect 2751 9938 2792 9940
rect 2705 9888 2792 9938
rect 2844 9888 2864 9940
rect 2705 9856 2864 9888
rect 2751 9810 2864 9856
rect 2705 9754 2864 9810
rect 2705 9729 2792 9754
rect 2751 9702 2792 9729
rect 2844 9702 2864 9754
rect 2751 9683 2864 9702
rect 2705 9662 2864 9683
rect 2705 9661 2788 9662
rect 2705 9602 2751 9661
rect 2705 9543 2751 9556
rect 2123 9225 2157 9239
rect 2115 9221 2157 9225
rect 2041 9087 2157 9221
rect 2041 9035 2063 9087
rect 2115 9035 2157 9087
rect 2041 8995 2157 9035
rect 2481 9145 2527 9206
rect 2481 9038 2527 9099
rect 2481 8931 2527 8992
rect 1817 8795 2157 8915
rect 1431 8213 1444 8259
rect 1490 8213 1503 8259
rect 1431 8202 1503 8213
rect 1629 8712 1675 8725
rect 1629 8592 1675 8666
rect 801 8157 882 8170
rect 322 8131 390 8142
rect 322 7991 333 8131
rect 379 7991 390 8131
rect 322 7901 390 7991
rect 847 8111 882 8157
rect 1025 8157 1071 8170
rect 801 8058 882 8111
rect 1017 8111 1025 8143
rect 1249 8157 1347 8170
rect 1071 8111 1110 8143
rect 1017 8103 1110 8111
rect 801 8037 847 8058
rect 1017 8051 1037 8103
rect 1089 8051 1110 8103
rect 1017 8037 1110 8051
rect 1017 8010 1025 8037
rect 801 7978 847 7991
rect 1023 7991 1025 8010
rect 1071 8011 1110 8037
rect 1295 8111 1347 8157
rect 1249 8037 1347 8111
rect 1071 8010 1106 8011
rect 1071 7991 1095 8010
rect 1023 7901 1095 7991
rect 1295 7991 1347 8037
rect 1249 7978 1347 7991
rect 322 7827 1095 7901
rect 1275 7901 1347 7978
rect 1629 8136 1675 8546
rect 1629 8016 1675 8090
rect 1629 7901 1675 7970
rect 1275 7827 1675 7901
rect 1853 8712 1899 8725
rect 1853 8592 1899 8666
rect 1853 8136 1899 8546
rect 1853 8016 1899 8090
rect 1853 7831 1899 7970
rect 2041 8712 2157 8795
rect 2041 8666 2077 8712
rect 2123 8666 2157 8712
rect 2041 8592 2157 8666
rect 2041 8546 2077 8592
rect 2123 8546 2157 8592
rect 2041 8136 2157 8546
rect 2041 8090 2077 8136
rect 2123 8090 2157 8136
rect 2041 8016 2157 8090
rect 2041 7970 2077 8016
rect 2123 7970 2157 8016
rect 2041 7957 2157 7970
rect 2481 8824 2527 8885
rect 2481 8717 2527 8778
rect 2481 8610 2527 8671
rect 2481 8502 2527 8564
rect 2481 8394 2527 8456
rect 2481 8286 2527 8348
rect 2481 8178 2527 8240
rect 2481 8070 2527 8132
rect 2481 7962 2527 8024
rect 2481 7903 2527 7916
rect 2705 9252 2751 9265
rect 2705 9145 2751 9206
rect 2705 9047 2751 9099
rect 2705 9038 2864 9047
rect 2751 9017 2864 9038
rect 2751 8992 2792 9017
rect 2705 8965 2792 8992
rect 2844 8965 2864 9017
rect 2705 8931 2864 8965
rect 2751 8885 2864 8931
rect 2705 8831 2864 8885
rect 2705 8824 2792 8831
rect 2751 8779 2792 8824
rect 2844 8779 2864 8831
rect 2751 8778 2864 8779
rect 2705 8739 2864 8778
rect 2705 8717 2751 8739
rect 2705 8610 2751 8671
rect 2705 8502 2751 8564
rect 2705 8394 2751 8456
rect 2705 8286 2751 8348
rect 2705 8178 2751 8240
rect 2705 8070 2751 8132
rect 2705 7962 2751 8024
rect 2705 7903 2751 7916
rect 1853 7820 2650 7831
rect 1853 7774 2593 7820
rect 2639 7774 2650 7820
rect 1853 7757 2650 7774
rect 3416 7668 3620 7806
rect 1511 6327 1603 6368
rect 1511 6275 1531 6327
rect 1583 6275 1603 6327
rect 1511 6141 1603 6275
rect 1511 6089 1531 6141
rect 1583 6089 1603 6141
rect 1511 6049 1603 6089
rect 4639 5597 4715 5609
rect 4639 5441 4651 5597
rect 4703 5441 4715 5597
rect 4639 5429 4715 5441
rect 5125 5597 5201 5609
rect 5125 5441 5137 5597
rect 5189 5441 5201 5597
rect 5125 5429 5201 5441
rect 2257 3610 2349 3650
rect 2257 3558 2277 3610
rect 2329 3558 2349 3610
rect 2257 3424 2349 3558
rect 2257 3372 2277 3424
rect 2329 3372 2349 3424
rect 2257 3331 2349 3372
rect 2397 913 2470 1034
rect 2621 913 2741 1033
rect 3346 913 3466 1033
rect 2621 376 2741 566
rect 3346 376 3466 566
rect 5547 556 5623 568
rect 5547 192 5559 556
rect 5611 192 5623 556
rect 5547 180 5623 192
rect 828 -94 1008 -82
rect 828 -146 840 -94
rect 996 -146 1008 -94
rect 828 -158 1008 -146
rect 3000 -2259 3076 -2247
rect 3000 -2415 3012 -2259
rect 3064 -2415 3076 -2259
rect 3000 -2427 3076 -2415
<< via1 >>
rect 918 28925 970 28963
rect 1532 28925 1584 28963
rect 2157 28925 2209 28963
rect 2771 28925 2823 28963
rect 3395 28925 3447 28963
rect 4009 28925 4061 28963
rect 4634 28925 4686 28963
rect 5248 28925 5300 28963
rect 918 28911 964 28925
rect 964 28911 970 28925
rect 1532 28911 1538 28925
rect 1538 28911 1584 28925
rect 2157 28911 2203 28925
rect 2203 28911 2209 28925
rect 2771 28911 2777 28925
rect 2777 28911 2823 28925
rect 3395 28911 3441 28925
rect 3441 28911 3447 28925
rect 4009 28911 4015 28925
rect 4015 28911 4061 28925
rect 4634 28911 4680 28925
rect 4680 28911 4686 28925
rect 5248 28911 5254 28925
rect 5254 28911 5300 28925
rect 918 28725 970 28777
rect 1532 28725 1584 28777
rect 2157 28725 2209 28777
rect 2771 28725 2823 28777
rect 3395 28725 3447 28777
rect 4009 28725 4061 28777
rect 4634 28725 4686 28777
rect 5248 28725 5300 28777
rect 914 28360 918 28393
rect 918 28360 964 28393
rect 964 28360 966 28393
rect 914 28237 966 28360
rect 914 27585 918 27618
rect 918 27585 964 27618
rect 964 27585 966 27618
rect 914 27462 966 27585
rect 1536 28360 1538 28393
rect 1538 28360 1584 28393
rect 1584 28360 1588 28393
rect 1536 28237 1588 28360
rect 1536 27585 1538 27618
rect 1538 27585 1584 27618
rect 1584 27585 1588 27618
rect 1536 27462 1588 27585
rect 2153 28360 2157 28393
rect 2157 28360 2203 28393
rect 2203 28360 2205 28393
rect 2153 28237 2205 28360
rect 2153 27585 2157 27618
rect 2157 27585 2203 27618
rect 2203 27585 2205 27618
rect 2153 27462 2205 27585
rect 2775 28360 2777 28393
rect 2777 28360 2823 28393
rect 2823 28360 2827 28393
rect 2775 28237 2827 28360
rect 2775 27585 2777 27618
rect 2777 27585 2823 27618
rect 2823 27585 2827 27618
rect 2775 27462 2827 27585
rect 3391 28360 3395 28393
rect 3395 28360 3441 28393
rect 3441 28360 3443 28393
rect 3391 28237 3443 28360
rect 3391 27585 3395 27618
rect 3395 27585 3441 27618
rect 3441 27585 3443 27618
rect 3391 27462 3443 27585
rect 4013 28360 4015 28393
rect 4015 28360 4061 28393
rect 4061 28360 4065 28393
rect 4013 28237 4065 28360
rect 4013 27585 4015 27618
rect 4015 27585 4061 27618
rect 4061 27585 4065 27618
rect 4013 27462 4065 27585
rect 4630 28360 4634 28393
rect 4634 28360 4680 28393
rect 4680 28360 4682 28393
rect 4630 28237 4682 28360
rect 4630 27585 4634 27618
rect 4634 27585 4680 27618
rect 4680 27585 4682 27618
rect 4630 27462 4682 27585
rect 5226 28360 5265 28393
rect 5265 28360 5278 28393
rect 5226 28341 5278 28360
rect 5226 28179 5265 28207
rect 5265 28179 5278 28207
rect 5226 28155 5278 28179
rect 5216 27585 5219 27618
rect 5219 27585 5265 27618
rect 5265 27585 5268 27618
rect 5216 27462 5268 27585
rect 499 27041 551 27093
rect 699 26242 751 26398
rect 1129 26242 1181 26398
rect 1321 26242 1373 26398
rect 1751 26242 1803 26398
rect 1938 26242 1990 26398
rect 2368 26242 2420 26398
rect 2560 26242 2612 26398
rect 2990 26242 3042 26398
rect 3176 26242 3228 26398
rect 3606 26242 3658 26398
rect 3798 26242 3850 26398
rect 4228 26242 4280 26398
rect 4415 26242 4467 26398
rect 4845 26242 4897 26398
rect 5041 26242 5093 26398
rect 5459 26242 5511 26398
rect 1117 25202 1169 25358
rect 1333 25202 1385 25358
rect 1225 24657 1277 24684
rect 1225 24424 1228 24657
rect 1228 24424 1274 24657
rect 1274 24424 1277 24657
rect 909 23924 961 23926
rect 909 23878 912 23924
rect 912 23878 958 23924
rect 958 23878 961 23924
rect 909 23770 961 23878
rect 1541 23924 1593 23926
rect 1541 23878 1544 23924
rect 1544 23878 1590 23924
rect 1590 23878 1593 23924
rect 1541 23770 1593 23878
rect 2356 25202 2408 25358
rect 2572 25202 2624 25358
rect 2464 24657 2516 24684
rect 2464 24424 2467 24657
rect 2467 24424 2513 24657
rect 2513 24424 2516 24657
rect 2148 23924 2200 23926
rect 2148 23878 2151 23924
rect 2151 23878 2197 23924
rect 2197 23878 2200 23924
rect 2148 23770 2200 23878
rect 1124 22173 1176 22225
rect 1326 22173 1378 22225
rect 2780 23924 2832 23926
rect 2780 23878 2783 23924
rect 2783 23878 2829 23924
rect 2829 23878 2832 23924
rect 2780 23770 2832 23878
rect 3594 25202 3646 25358
rect 3810 25202 3862 25358
rect 3702 24657 3754 24684
rect 3702 24424 3705 24657
rect 3705 24424 3751 24657
rect 3751 24424 3754 24657
rect 3386 23924 3438 23926
rect 3386 23878 3389 23924
rect 3389 23878 3435 23924
rect 3435 23878 3438 23924
rect 3386 23770 3438 23878
rect 2363 22173 2415 22225
rect 2565 22173 2617 22225
rect 4018 23924 4070 23926
rect 4018 23878 4021 23924
rect 4021 23878 4067 23924
rect 4067 23878 4070 23924
rect 4018 23770 4070 23878
rect 4833 25202 4885 25358
rect 5053 25202 5105 25358
rect 4941 24657 4993 24684
rect 4941 24424 4944 24657
rect 4944 24424 4990 24657
rect 4990 24424 4993 24657
rect 4625 23924 4677 23926
rect 4625 23878 4628 23924
rect 4628 23878 4674 23924
rect 4674 23878 4677 23924
rect 4625 23770 4677 23878
rect 3601 22173 3653 22225
rect 3803 22173 3855 22225
rect 5257 23924 5309 23926
rect 5257 23878 5260 23924
rect 5260 23878 5306 23924
rect 5306 23878 5309 23924
rect 5257 23770 5309 23878
rect 4840 22173 4892 22225
rect 5042 22173 5094 22225
rect 831 21975 883 22027
rect 1619 21975 1671 22027
rect 2070 21975 2122 22027
rect 2858 21975 2910 22027
rect 3308 21975 3360 22027
rect 4096 21975 4148 22027
rect 4547 21975 4599 22027
rect 5314 21975 5366 22027
rect 699 21767 751 21819
rect 913 20183 918 20219
rect 918 20183 964 20219
rect 964 20183 965 20219
rect 913 20167 965 20183
rect 915 19952 967 19955
rect 915 19906 918 19952
rect 918 19906 964 19952
rect 964 19906 967 19952
rect 915 19903 967 19906
rect 1751 21767 1803 21819
rect 1938 21767 1990 21819
rect 1537 20183 1538 20219
rect 1538 20183 1584 20219
rect 1584 20183 1589 20219
rect 1537 20167 1589 20183
rect 1535 19952 1587 19955
rect 1535 19906 1538 19952
rect 1538 19906 1584 19952
rect 1584 19906 1587 19952
rect 1535 19903 1587 19906
rect 714 18326 766 18378
rect 2152 20183 2157 20219
rect 2157 20183 2203 20219
rect 2203 20183 2204 20219
rect 2152 20167 2204 20183
rect 2154 19952 2206 19955
rect 2154 19906 2157 19952
rect 2157 19906 2203 19952
rect 2203 19906 2206 19952
rect 2154 19903 2206 19906
rect 2990 21767 3042 21819
rect 3176 21767 3228 21819
rect 2776 20183 2777 20219
rect 2777 20183 2823 20219
rect 2823 20183 2828 20219
rect 2776 20167 2828 20183
rect 2774 19952 2826 19955
rect 2774 19906 2777 19952
rect 2777 19906 2823 19952
rect 2823 19906 2826 19952
rect 2774 19903 2826 19906
rect 1747 18334 1799 18386
rect 1933 18334 1985 18386
rect 3390 20183 3395 20219
rect 3395 20183 3441 20219
rect 3441 20183 3442 20219
rect 3390 20167 3442 20183
rect 3392 19952 3444 19955
rect 3392 19906 3395 19952
rect 3395 19906 3441 19952
rect 3441 19906 3444 19952
rect 3392 19903 3444 19906
rect 4228 21767 4280 21819
rect 4415 21767 4467 21819
rect 4014 20183 4015 20219
rect 4015 20183 4061 20219
rect 4061 20183 4066 20219
rect 4014 20167 4066 20183
rect 4012 19952 4064 19955
rect 4012 19906 4015 19952
rect 4015 19906 4061 19952
rect 4061 19906 4064 19952
rect 4012 19903 4064 19906
rect 2985 18334 3037 18386
rect 3171 18334 3223 18386
rect 4629 20183 4634 20219
rect 4634 20183 4680 20219
rect 4680 20183 4681 20219
rect 4629 20167 4681 20183
rect 4631 19952 4683 19955
rect 4631 19906 4634 19952
rect 4634 19906 4680 19952
rect 4680 19906 4683 19952
rect 4631 19903 4683 19906
rect 5459 21766 5511 21818
rect 5253 20183 5254 20219
rect 5254 20183 5300 20219
rect 5300 20183 5305 20219
rect 5253 20167 5305 20183
rect 5251 19952 5303 19956
rect 5251 19906 5254 19952
rect 5254 19906 5300 19952
rect 5300 19906 5303 19952
rect 5251 19904 5303 19906
rect 4224 18334 4276 18386
rect 4410 18334 4462 18386
rect 5453 18326 5505 18378
rect 1699 18175 1751 18178
rect 1699 18129 1702 18175
rect 1702 18129 1748 18175
rect 1748 18129 1751 18175
rect 1699 18126 1751 18129
rect 1990 18175 2042 18178
rect 2938 18175 2990 18178
rect 1990 18129 1993 18175
rect 1993 18129 2039 18175
rect 2039 18129 2042 18175
rect 2938 18129 2941 18175
rect 2941 18129 2987 18175
rect 2987 18129 2990 18175
rect 1990 18126 2042 18129
rect 2938 18126 2990 18129
rect 3229 18175 3281 18178
rect 4176 18175 4228 18178
rect 3229 18129 3231 18175
rect 3231 18129 3277 18175
rect 3277 18129 3281 18175
rect 4176 18129 4179 18175
rect 4179 18129 4225 18175
rect 4225 18129 4228 18175
rect 3229 18126 3281 18129
rect 4176 18126 4228 18129
rect 4467 18175 4519 18178
rect 4467 18129 4470 18175
rect 4470 18129 4516 18175
rect 4516 18129 4519 18175
rect 4467 18126 4519 18129
rect 913 17935 965 17987
rect 973 17720 1025 17824
rect 973 17674 975 17720
rect 975 17674 1021 17720
rect 1021 17674 1025 17720
rect 973 17668 1025 17674
rect 1537 17935 1589 17987
rect 2152 17935 2204 17987
rect 1477 17720 1529 17824
rect 1477 17674 1481 17720
rect 1481 17674 1527 17720
rect 1527 17674 1529 17720
rect 1477 17668 1529 17674
rect 2212 17720 2264 17824
rect 2212 17674 2214 17720
rect 2214 17674 2260 17720
rect 2260 17674 2264 17720
rect 2212 17668 2264 17674
rect 2776 17935 2828 17987
rect 3390 17935 3442 17987
rect 2716 17720 2768 17824
rect 2716 17674 2720 17720
rect 2720 17674 2766 17720
rect 2766 17674 2768 17720
rect 2716 17668 2768 17674
rect 3450 17720 3502 17824
rect 3450 17674 3452 17720
rect 3452 17674 3498 17720
rect 3498 17674 3502 17720
rect 3450 17668 3502 17674
rect 4014 17935 4066 17987
rect 4629 17935 4681 17987
rect 3954 17720 4006 17824
rect 3954 17674 3958 17720
rect 3958 17674 4004 17720
rect 4004 17674 4006 17720
rect 3954 17668 4006 17674
rect 4689 17720 4741 17824
rect 4689 17674 4691 17720
rect 4691 17674 4737 17720
rect 4737 17674 4741 17720
rect 4689 17668 4741 17674
rect 5254 17936 5306 17988
rect 5174 17720 5226 17824
rect 5174 17674 5197 17720
rect 5197 17674 5226 17720
rect 5174 17668 5226 17674
rect 915 16888 967 16940
rect 1535 16888 1587 16940
rect 2154 16888 2206 16940
rect 2774 16888 2826 16940
rect 3392 16888 3444 16940
rect 4012 16888 4064 16940
rect 4631 16888 4683 16940
rect 5251 16888 5303 16940
rect 728 16571 780 16623
rect 914 16571 966 16623
rect 1745 16571 1797 16623
rect 1931 16571 1983 16623
rect 1108 16363 1160 16415
rect 1294 16363 1346 16415
rect 2346 16363 2398 16415
rect 2532 16363 2584 16415
rect 4854 16363 4906 16415
rect 5040 16363 5092 16415
rect 967 16138 1019 16190
rect 1761 16138 1813 16190
rect 1972 16138 2024 16190
rect 2182 16138 2234 16190
rect 2393 16138 2445 16190
rect 2605 16138 2657 16190
rect 2816 16138 2868 16190
rect 3026 16138 3078 16190
rect 3237 16138 3289 16190
rect 3713 16138 3765 16190
rect 3924 16138 3976 16190
rect 4136 16138 4188 16190
rect 4347 16138 4399 16190
rect 499 15901 551 15953
rect 2278 15884 2330 15936
rect 297 15560 300 15612
rect 300 15560 346 15612
rect 346 15560 349 15612
rect 297 15374 300 15426
rect 300 15374 346 15426
rect 346 15374 349 15426
rect 297 14961 300 15013
rect 300 14961 346 15013
rect 346 14961 349 15013
rect 297 14775 300 14827
rect 300 14775 346 14827
rect 346 14775 349 14827
rect 297 13504 300 13556
rect 300 13504 346 13556
rect 346 13504 349 13556
rect 297 13318 300 13370
rect 300 13318 346 13370
rect 346 13318 349 13370
rect 1419 15689 1471 15741
rect 2278 15698 2330 15750
rect 967 15322 990 15365
rect 990 15322 1019 15365
rect 967 15313 1019 15322
rect 1419 15503 1471 15555
rect 1657 15562 1709 15565
rect 1843 15562 1895 15565
rect 1657 15516 1665 15562
rect 1665 15516 1709 15562
rect 1843 15516 1895 15562
rect 1657 15513 1709 15516
rect 1843 15513 1895 15516
rect 1377 15095 1429 15147
rect 1377 14909 1429 14961
rect 1867 14999 1919 15047
rect 1867 14995 1868 14999
rect 1868 14995 1914 14999
rect 1914 14995 1919 14999
rect 1867 14849 1868 14861
rect 1868 14849 1914 14861
rect 1914 14849 1919 14861
rect 1867 14809 1919 14849
rect 740 14306 792 14358
rect 740 14145 748 14172
rect 748 14145 792 14172
rect 740 14120 792 14145
rect 1193 14306 1245 14358
rect 1193 14145 1196 14172
rect 1196 14145 1242 14172
rect 1242 14145 1245 14172
rect 1193 14120 1245 14145
rect 1867 13535 1919 13556
rect 1867 13504 1868 13535
rect 1868 13504 1914 13535
rect 1914 13504 1919 13535
rect 1867 13325 1919 13370
rect 1867 13318 1868 13325
rect 1868 13318 1914 13325
rect 1914 13318 1919 13325
rect 297 12509 300 12561
rect 300 12509 346 12561
rect 346 12509 349 12561
rect 297 12323 300 12375
rect 300 12323 346 12375
rect 346 12323 349 12375
rect 297 11561 300 11613
rect 300 11561 346 11613
rect 346 11561 349 11613
rect 297 11375 300 11427
rect 300 11375 346 11427
rect 346 11375 349 11427
rect 297 10645 300 10697
rect 300 10645 346 10697
rect 346 10645 349 10697
rect 297 10459 300 10511
rect 300 10459 346 10511
rect 346 10459 349 10511
rect 743 12560 748 12567
rect 748 12560 794 12567
rect 794 12560 795 12567
rect 743 12515 795 12560
rect 743 12352 748 12381
rect 748 12352 794 12381
rect 794 12352 795 12381
rect 743 12329 795 12352
rect 1193 12560 1196 12567
rect 1196 12560 1242 12567
rect 1242 12560 1245 12567
rect 1193 12515 1245 12560
rect 1193 12352 1196 12381
rect 1196 12352 1242 12381
rect 1242 12352 1245 12381
rect 1193 12329 1245 12352
rect 2093 12577 2145 12629
rect 1854 12560 1868 12561
rect 1868 12560 1906 12561
rect 1854 12509 1906 12560
rect 2093 12391 2145 12443
rect 1854 12352 1868 12375
rect 1868 12352 1906 12375
rect 1854 12323 1906 12352
rect 2093 11801 2145 11853
rect 2093 11615 2145 11667
rect 1854 11565 1906 11613
rect 1854 11561 1868 11565
rect 1868 11561 1906 11565
rect 1854 11414 1868 11427
rect 1868 11414 1906 11427
rect 1854 11375 1906 11414
rect 2093 10885 2145 10937
rect 2093 10699 2145 10751
rect 1854 10679 1868 10697
rect 1868 10679 1906 10697
rect 1854 10645 1906 10679
rect 1854 10469 1868 10511
rect 1868 10469 1906 10511
rect 1854 10459 1906 10469
rect 978 10219 1022 10255
rect 1022 10219 1030 10255
rect 978 10203 1030 10219
rect 5365 10194 5417 10246
rect 5365 10008 5417 10060
rect 918 9798 970 9845
rect 918 9793 957 9798
rect 957 9793 970 9798
rect 918 9632 957 9659
rect 957 9632 970 9659
rect 918 9607 970 9632
rect 296 9480 300 9525
rect 300 9480 346 9525
rect 346 9480 348 9525
rect 296 9473 348 9480
rect 508 9473 560 9525
rect 1636 9793 1688 9845
rect 1636 9607 1688 9659
rect 603 9052 655 9104
rect 789 9078 841 9104
rect 789 9052 801 9078
rect 801 9052 841 9078
rect 1241 9078 1293 9087
rect 1241 9035 1249 9078
rect 1249 9035 1293 9078
rect 297 8978 349 8988
rect 297 8936 300 8978
rect 300 8936 346 8978
rect 346 8936 349 8978
rect 297 8768 300 8802
rect 300 8768 346 8802
rect 346 8768 349 8802
rect 297 8750 349 8768
rect 647 8818 699 8870
rect 833 8841 875 8870
rect 875 8841 885 8870
rect 833 8818 885 8841
rect 1241 8849 1293 8901
rect 1630 9035 1682 9087
rect 2063 9271 2115 9273
rect 1059 8686 1111 8738
rect 481 8478 533 8530
rect 1059 8510 1111 8552
rect 1059 8500 1071 8510
rect 1071 8500 1111 8510
rect 481 8292 533 8344
rect 1630 8849 1682 8901
rect 2063 9225 2077 9271
rect 2077 9225 2115 9271
rect 2792 9888 2844 9940
rect 2792 9702 2844 9754
rect 2063 9221 2115 9225
rect 2063 9035 2115 9087
rect 1037 8051 1089 8103
rect 2792 8965 2844 9017
rect 2792 8779 2844 8831
rect 1531 6275 1583 6327
rect 1531 6089 1583 6141
rect 4651 5441 4703 5597
rect 5137 5441 5189 5597
rect 2277 3558 2329 3610
rect 2277 3372 2329 3424
rect 5559 536 5611 556
rect 5559 208 5562 536
rect 5562 208 5608 536
rect 5608 208 5611 536
rect 5559 192 5611 208
rect 840 -146 996 -94
rect 3012 -2415 3064 -2259
<< metal2 >>
rect 697 27568 753 28985
rect 877 28965 1005 28987
rect 877 28909 916 28965
rect 972 28909 1005 28965
rect 877 28779 1005 28909
rect 877 28723 916 28779
rect 972 28723 1005 28779
rect 877 28704 1005 28723
rect 902 28393 978 28405
rect 902 28237 914 28393
rect 966 28344 978 28393
rect 1127 28344 1183 28985
rect 966 28288 1183 28344
rect 966 28237 978 28288
rect 902 28225 978 28237
rect 902 27618 978 27630
rect 902 27568 914 27618
rect 697 27512 914 27568
rect 487 27093 563 27105
rect 487 27041 499 27093
rect 551 27041 563 27093
rect 487 27029 563 27041
rect 497 15965 553 27029
rect 697 26410 753 27512
rect 902 27462 914 27512
rect 966 27462 978 27618
rect 902 27450 978 27462
rect 1127 26410 1183 28288
rect 1319 28344 1375 28985
rect 1497 28965 1625 28987
rect 1497 28909 1530 28965
rect 1586 28909 1625 28965
rect 1497 28779 1625 28909
rect 1497 28723 1530 28779
rect 1586 28723 1625 28779
rect 1497 28704 1625 28723
rect 1524 28393 1600 28405
rect 1524 28344 1536 28393
rect 1319 28288 1536 28344
rect 1319 26410 1375 28288
rect 1524 28237 1536 28288
rect 1588 28237 1600 28393
rect 1524 28225 1600 28237
rect 1524 27618 1600 27630
rect 1524 27462 1536 27618
rect 1588 27568 1600 27618
rect 1749 27568 1805 28985
rect 1588 27512 1805 27568
rect 1588 27462 1600 27512
rect 1524 27450 1600 27462
rect 1749 26410 1805 27512
rect 1936 27568 1992 28985
rect 2116 28965 2244 28987
rect 2116 28909 2155 28965
rect 2211 28909 2244 28965
rect 2116 28779 2244 28909
rect 2116 28723 2155 28779
rect 2211 28723 2244 28779
rect 2116 28704 2244 28723
rect 2141 28393 2217 28405
rect 2141 28237 2153 28393
rect 2205 28344 2217 28393
rect 2366 28344 2422 28985
rect 2205 28288 2422 28344
rect 2205 28237 2217 28288
rect 2141 28225 2217 28237
rect 2141 27618 2217 27630
rect 2141 27568 2153 27618
rect 1936 27512 2153 27568
rect 1936 26410 1992 27512
rect 2141 27462 2153 27512
rect 2205 27462 2217 27618
rect 2141 27450 2217 27462
rect 2366 26410 2422 28288
rect 2558 28344 2614 28985
rect 2736 28965 2864 28987
rect 2736 28909 2769 28965
rect 2825 28909 2864 28965
rect 2736 28779 2864 28909
rect 2736 28723 2769 28779
rect 2825 28723 2864 28779
rect 2736 28704 2864 28723
rect 2763 28393 2839 28405
rect 2763 28344 2775 28393
rect 2558 28288 2775 28344
rect 2558 26410 2614 28288
rect 2763 28237 2775 28288
rect 2827 28237 2839 28393
rect 2763 28225 2839 28237
rect 2763 27618 2839 27630
rect 2763 27462 2775 27618
rect 2827 27568 2839 27618
rect 2988 27568 3044 28985
rect 2827 27512 3044 27568
rect 2827 27462 2839 27512
rect 2763 27450 2839 27462
rect 2988 26410 3044 27512
rect 3174 27568 3230 28985
rect 3354 28965 3482 28987
rect 3354 28909 3393 28965
rect 3449 28909 3482 28965
rect 3354 28779 3482 28909
rect 3354 28723 3393 28779
rect 3449 28723 3482 28779
rect 3354 28704 3482 28723
rect 3379 28393 3455 28405
rect 3379 28237 3391 28393
rect 3443 28344 3455 28393
rect 3604 28344 3660 28985
rect 3443 28288 3660 28344
rect 3443 28237 3455 28288
rect 3379 28225 3455 28237
rect 3379 27618 3455 27630
rect 3379 27568 3391 27618
rect 3174 27512 3391 27568
rect 3174 26410 3230 27512
rect 3379 27462 3391 27512
rect 3443 27462 3455 27618
rect 3379 27450 3455 27462
rect 3604 26410 3660 28288
rect 3796 28344 3852 28985
rect 3974 28965 4102 28987
rect 3974 28909 4007 28965
rect 4063 28909 4102 28965
rect 3974 28779 4102 28909
rect 3974 28723 4007 28779
rect 4063 28723 4102 28779
rect 3974 28704 4102 28723
rect 4001 28393 4077 28405
rect 4001 28344 4013 28393
rect 3796 28288 4013 28344
rect 3796 26410 3852 28288
rect 4001 28237 4013 28288
rect 4065 28237 4077 28393
rect 4001 28225 4077 28237
rect 4001 27618 4077 27630
rect 4001 27462 4013 27618
rect 4065 27568 4077 27618
rect 4226 27568 4282 28985
rect 4065 27512 4282 27568
rect 4065 27462 4077 27512
rect 4001 27450 4077 27462
rect 4226 26410 4282 27512
rect 4413 27568 4469 28985
rect 4593 28965 4721 28987
rect 4593 28909 4632 28965
rect 4688 28909 4721 28965
rect 4593 28779 4721 28909
rect 4593 28723 4632 28779
rect 4688 28723 4721 28779
rect 4593 28704 4721 28723
rect 4618 28393 4694 28405
rect 4618 28237 4630 28393
rect 4682 28344 4694 28393
rect 4843 28344 4899 28985
rect 4682 28288 4899 28344
rect 4682 28237 4694 28288
rect 4618 28225 4694 28237
rect 4618 27618 4694 27630
rect 4618 27568 4630 27618
rect 4413 27512 4630 27568
rect 4413 26410 4469 27512
rect 4618 27462 4630 27512
rect 4682 27462 4694 27618
rect 4618 27450 4694 27462
rect 4843 26410 4899 28288
rect 5039 28344 5095 29035
rect 5212 28965 5341 28987
rect 5212 28909 5246 28965
rect 5302 28909 5341 28965
rect 5212 28779 5341 28909
rect 5212 28723 5246 28779
rect 5302 28723 5341 28779
rect 5212 28704 5341 28723
rect 5206 28393 5298 28433
rect 5206 28344 5226 28393
rect 5039 28341 5226 28344
rect 5278 28341 5298 28393
rect 5039 28288 5298 28341
rect 5039 26410 5095 28288
rect 5206 28207 5298 28288
rect 5206 28155 5226 28207
rect 5278 28155 5298 28207
rect 5206 28115 5298 28155
rect 5204 27618 5280 27630
rect 5204 27462 5216 27618
rect 5268 27568 5280 27618
rect 5457 27568 5513 29035
rect 5268 27512 5513 27568
rect 5268 27462 5280 27512
rect 5204 27450 5280 27462
rect 5457 26410 5513 27512
rect 687 26398 763 26410
rect 687 26242 699 26398
rect 751 26242 763 26398
rect 687 26230 763 26242
rect 1117 26398 1193 26410
rect 1117 26242 1129 26398
rect 1181 26242 1193 26398
rect 1117 26230 1193 26242
rect 1309 26398 1385 26410
rect 1309 26242 1321 26398
rect 1373 26242 1385 26398
rect 1309 26230 1385 26242
rect 1739 26398 1815 26410
rect 1739 26242 1751 26398
rect 1803 26242 1815 26398
rect 1739 26230 1815 26242
rect 1926 26398 2002 26410
rect 1926 26242 1938 26398
rect 1990 26242 2002 26398
rect 1926 26230 2002 26242
rect 2356 26398 2432 26410
rect 2356 26242 2368 26398
rect 2420 26242 2432 26398
rect 2356 26230 2432 26242
rect 2548 26398 2624 26410
rect 2548 26242 2560 26398
rect 2612 26242 2624 26398
rect 2548 26230 2624 26242
rect 2978 26398 3054 26410
rect 2978 26242 2990 26398
rect 3042 26242 3054 26398
rect 2978 26230 3054 26242
rect 3164 26398 3240 26410
rect 3164 26242 3176 26398
rect 3228 26242 3240 26398
rect 3164 26230 3240 26242
rect 3594 26398 3670 26410
rect 3594 26242 3606 26398
rect 3658 26242 3670 26398
rect 3594 26230 3670 26242
rect 3786 26398 3862 26410
rect 3786 26242 3798 26398
rect 3850 26242 3862 26398
rect 3786 26230 3862 26242
rect 4216 26398 4292 26410
rect 4216 26242 4228 26398
rect 4280 26242 4292 26398
rect 4216 26230 4292 26242
rect 4403 26398 4479 26410
rect 4403 26242 4415 26398
rect 4467 26242 4479 26398
rect 4403 26230 4479 26242
rect 4833 26398 4909 26410
rect 4833 26242 4845 26398
rect 4897 26242 4909 26398
rect 4833 26230 4909 26242
rect 5029 26398 5105 26410
rect 5029 26242 5041 26398
rect 5093 26242 5105 26398
rect 5029 26230 5105 26242
rect 5447 26398 5523 26410
rect 5447 26242 5459 26398
rect 5511 26242 5523 26398
rect 5447 26230 5523 26242
rect 697 21831 753 26230
rect 1127 25370 1183 26230
rect 1105 25358 1183 25370
rect 1105 25202 1117 25358
rect 1169 25202 1183 25358
rect 1105 25190 1183 25202
rect 1319 25370 1375 26230
rect 1319 25358 1397 25370
rect 1319 25202 1333 25358
rect 1385 25202 1397 25358
rect 1319 25190 1397 25202
rect 1213 24686 1289 24696
rect 1213 24422 1223 24686
rect 1279 24422 1289 24686
rect 1213 24412 1289 24422
rect 897 23926 973 23938
rect 897 23770 909 23926
rect 961 23770 973 23926
rect 897 23758 973 23770
rect 1529 23926 1605 23938
rect 1529 23770 1541 23926
rect 1593 23770 1605 23926
rect 1529 23758 1605 23770
rect 907 22157 963 23758
rect 1112 22225 1390 22237
rect 1112 22173 1124 22225
rect 1176 22173 1326 22225
rect 1378 22173 1390 22225
rect 1112 22161 1390 22173
rect 907 22101 1030 22157
rect 819 22027 895 22039
rect 819 22016 831 22027
rect 883 22016 895 22027
rect 819 21856 829 22016
rect 885 21856 895 22016
rect 819 21846 895 21856
rect 687 21819 763 21831
rect 687 21767 699 21819
rect 751 21767 763 21819
rect 687 21755 763 21767
rect 678 21224 770 21277
rect 678 21186 772 21224
rect 678 21130 697 21186
rect 753 21130 772 21186
rect 678 21091 772 21130
rect 678 20243 770 21091
rect 974 20415 1030 22101
rect 974 20359 1138 20415
rect 678 20219 1001 20243
rect 678 20167 913 20219
rect 965 20167 1001 20219
rect 678 20146 1001 20167
rect 678 18613 770 20146
rect 903 19957 979 19967
rect 1082 19957 1138 20359
rect 903 19955 1138 19957
rect 903 19903 915 19955
rect 967 19903 1138 19955
rect 903 19901 1138 19903
rect 903 19891 979 19901
rect 678 18516 977 18613
rect 702 18378 778 18390
rect 702 18326 714 18378
rect 766 18326 778 18378
rect 702 16648 778 18326
rect 901 17987 977 18516
rect 901 17935 913 17987
rect 965 17935 977 17987
rect 901 17915 977 17935
rect 1082 17836 1138 19901
rect 961 17824 1138 17836
rect 961 17668 973 17824
rect 1025 17668 1138 17824
rect 961 17656 1138 17668
rect 877 16942 1005 17038
rect 877 16886 913 16942
rect 969 16886 1005 16942
rect 877 16809 1005 16886
rect 1223 16761 1279 22161
rect 1539 22157 1595 23758
rect 1472 22101 1595 22157
rect 1472 20415 1528 22101
rect 1607 22027 1683 22039
rect 1607 22016 1619 22027
rect 1671 22016 1683 22027
rect 1607 21856 1617 22016
rect 1673 21856 1683 22016
rect 1607 21846 1683 21856
rect 1749 21831 1805 26230
rect 1936 21831 1992 26230
rect 2366 25370 2422 26230
rect 2344 25358 2422 25370
rect 2344 25202 2356 25358
rect 2408 25202 2422 25358
rect 2344 25190 2422 25202
rect 2558 25370 2614 26230
rect 2558 25358 2636 25370
rect 2558 25202 2572 25358
rect 2624 25202 2636 25358
rect 2558 25190 2636 25202
rect 2452 24686 2528 24696
rect 2452 24422 2462 24686
rect 2518 24422 2528 24686
rect 2452 24412 2528 24422
rect 2136 23926 2212 23938
rect 2136 23770 2148 23926
rect 2200 23770 2212 23926
rect 2136 23758 2212 23770
rect 2768 23926 2844 23938
rect 2768 23770 2780 23926
rect 2832 23770 2844 23926
rect 2768 23758 2844 23770
rect 2146 22157 2202 23758
rect 2351 22225 2629 22237
rect 2351 22173 2363 22225
rect 2415 22173 2565 22225
rect 2617 22173 2629 22225
rect 2351 22161 2629 22173
rect 2146 22101 2269 22157
rect 2058 22027 2134 22039
rect 2058 22016 2070 22027
rect 2122 22016 2134 22027
rect 2058 21856 2068 22016
rect 2124 21856 2134 22016
rect 2058 21846 2134 21856
rect 1739 21819 1815 21831
rect 1739 21767 1751 21819
rect 1803 21767 1815 21819
rect 1739 21755 1815 21767
rect 1926 21819 2002 21831
rect 1926 21767 1938 21819
rect 1990 21767 2002 21819
rect 1926 21755 2002 21767
rect 1364 20359 1528 20415
rect 1732 20905 1824 21277
rect 1732 20867 1826 20905
rect 1732 20811 1751 20867
rect 1807 20811 1826 20867
rect 1732 20772 1826 20811
rect 1364 19957 1420 20359
rect 1732 20243 1824 20772
rect 1917 20576 2009 21277
rect 1916 20538 2010 20576
rect 1916 20482 1935 20538
rect 1991 20482 2010 20538
rect 1916 20443 2010 20482
rect 1501 20219 1824 20243
rect 1501 20167 1537 20219
rect 1589 20167 1824 20219
rect 1501 20146 1824 20167
rect 1523 19957 1599 19967
rect 1364 19955 1599 19957
rect 1364 19903 1535 19955
rect 1587 19903 1599 19955
rect 1364 19901 1599 19903
rect 1364 17836 1420 19901
rect 1523 19891 1599 19901
rect 1732 18613 1824 20146
rect 1525 18516 1824 18613
rect 1917 20243 2009 20443
rect 2213 20415 2269 22101
rect 2213 20359 2377 20415
rect 1917 20219 2240 20243
rect 1917 20167 2152 20219
rect 2204 20167 2240 20219
rect 1917 20146 2240 20167
rect 1917 18613 2009 20146
rect 2142 19957 2218 19967
rect 2321 19957 2377 20359
rect 2142 19955 2377 19957
rect 2142 19903 2154 19955
rect 2206 19903 2377 19955
rect 2142 19901 2377 19903
rect 2142 19891 2218 19901
rect 1917 18516 2216 18613
rect 1525 17987 1601 18516
rect 1717 18386 2025 18406
rect 1717 18334 1747 18386
rect 1799 18334 1933 18386
rect 1985 18334 2025 18386
rect 1717 18314 2025 18334
rect 1525 17935 1537 17987
rect 1589 17935 1601 17987
rect 1525 17915 1601 17935
rect 1687 18180 1763 18202
rect 1687 18020 1697 18180
rect 1753 18020 1763 18180
rect 1687 17920 1763 18020
rect 1364 17824 1541 17836
rect 1364 17668 1477 17824
rect 1529 17668 1541 17824
rect 1364 17656 1541 17668
rect 1497 16942 1625 17038
rect 1497 16886 1533 16942
rect 1589 16886 1625 16942
rect 1497 16809 1625 16886
rect 702 16643 814 16648
rect 698 16623 1006 16643
rect 698 16571 728 16623
rect 780 16571 914 16623
rect 966 16571 1006 16623
rect 698 16551 1006 16571
rect 487 15953 563 15965
rect 487 15901 499 15953
rect 551 15901 563 15953
rect 487 15889 563 15901
rect 277 15614 369 15642
rect 277 15558 295 15614
rect 351 15558 369 15614
rect 277 15428 369 15558
rect 277 15372 295 15428
rect 351 15372 369 15428
rect 277 15334 369 15372
rect 277 15015 369 15043
rect 277 14959 295 15015
rect 351 14959 369 15015
rect 277 14829 369 14959
rect 277 14773 295 14829
rect 351 14773 369 14829
rect 277 14735 369 14773
rect 719 14358 814 16551
rect 1207 16439 1297 16761
rect 1172 16435 1297 16439
rect 1078 16415 1386 16435
rect 1078 16363 1108 16415
rect 1160 16363 1294 16415
rect 1346 16363 1386 16415
rect 1078 16343 1386 16363
rect 1172 16342 1297 16343
rect 928 16192 1058 16231
rect 928 16136 965 16192
rect 1021 16136 1058 16192
rect 928 16097 1058 16136
rect 719 14306 740 14358
rect 792 14306 814 14358
rect 719 14172 814 14306
rect 719 14120 740 14172
rect 792 14120 814 14172
rect 277 13558 369 13586
rect 277 13502 295 13558
rect 351 13502 369 13558
rect 277 13372 369 13502
rect 277 13316 295 13372
rect 351 13316 369 13372
rect 277 13278 369 13316
rect 719 12607 814 14120
rect 946 15365 1040 16097
rect 946 15313 967 15365
rect 1019 15313 1040 15365
rect 277 12563 369 12591
rect 277 12507 295 12563
rect 351 12507 369 12563
rect 277 12377 369 12507
rect 277 12321 295 12377
rect 351 12321 369 12377
rect 277 12283 369 12321
rect 719 12567 815 12607
rect 719 12515 743 12567
rect 795 12515 815 12567
rect 719 12381 815 12515
rect 719 12329 743 12381
rect 795 12329 815 12381
rect 719 12289 815 12329
rect 277 11615 369 11643
rect 277 11559 295 11615
rect 351 11559 369 11615
rect 277 11429 369 11559
rect 277 11373 295 11429
rect 351 11373 369 11429
rect 277 11335 369 11373
rect 277 10699 369 10727
rect 277 10643 295 10699
rect 351 10643 369 10699
rect 277 10513 369 10643
rect 277 10457 295 10513
rect 351 10457 369 10513
rect 277 10419 369 10457
rect 946 10276 1040 15313
rect 1172 14358 1266 16342
rect 1514 15782 1608 16809
rect 1826 16643 1916 18314
rect 1978 18180 2054 18202
rect 1978 18020 1988 18180
rect 2044 18020 2054 18180
rect 1978 17920 2054 18020
rect 2140 17987 2216 18516
rect 2140 17935 2152 17987
rect 2204 17935 2216 17987
rect 2140 17915 2216 17935
rect 2321 17836 2377 19901
rect 2200 17824 2377 17836
rect 2200 17668 2212 17824
rect 2264 17668 2377 17824
rect 2200 17656 2377 17668
rect 2116 16942 2244 17038
rect 2116 16886 2152 16942
rect 2208 16886 2244 16942
rect 2116 16809 2244 16886
rect 2462 16761 2518 22161
rect 2778 22157 2834 23758
rect 2711 22101 2834 22157
rect 2711 20415 2767 22101
rect 2846 22027 2922 22039
rect 2846 22016 2858 22027
rect 2910 22016 2922 22027
rect 2846 21856 2856 22016
rect 2912 21856 2922 22016
rect 2846 21846 2922 21856
rect 2988 21831 3044 26230
rect 3174 21831 3230 26230
rect 3604 25370 3660 26230
rect 3582 25358 3660 25370
rect 3582 25202 3594 25358
rect 3646 25202 3660 25358
rect 3582 25190 3660 25202
rect 3796 25370 3852 26230
rect 3796 25358 3874 25370
rect 3796 25202 3810 25358
rect 3862 25202 3874 25358
rect 3796 25190 3874 25202
rect 3690 24686 3766 24696
rect 3690 24422 3700 24686
rect 3756 24422 3766 24686
rect 3690 24412 3766 24422
rect 3374 23926 3450 23938
rect 3374 23770 3386 23926
rect 3438 23770 3450 23926
rect 3374 23758 3450 23770
rect 4006 23926 4082 23938
rect 4006 23770 4018 23926
rect 4070 23770 4082 23926
rect 4006 23758 4082 23770
rect 3384 22157 3440 23758
rect 3589 22225 3867 22237
rect 3589 22173 3601 22225
rect 3653 22173 3803 22225
rect 3855 22173 3867 22225
rect 3589 22161 3867 22173
rect 3384 22101 3507 22157
rect 3296 22027 3372 22039
rect 3296 22016 3308 22027
rect 3360 22016 3372 22027
rect 3296 21856 3306 22016
rect 3362 21856 3372 22016
rect 3296 21846 3372 21856
rect 2978 21819 3054 21831
rect 2978 21767 2990 21819
rect 3042 21767 3054 21819
rect 2978 21755 3054 21767
rect 3164 21819 3240 21831
rect 3164 21767 3176 21819
rect 3228 21767 3240 21819
rect 3164 21755 3240 21767
rect 2603 20359 2767 20415
rect 2603 19957 2659 20359
rect 2971 20254 3063 21277
rect 2970 20243 3064 20254
rect 2740 20219 3064 20243
rect 2740 20167 2776 20219
rect 2828 20216 3064 20219
rect 2828 20167 2989 20216
rect 2740 20160 2989 20167
rect 3045 20160 3064 20216
rect 2740 20146 3064 20160
rect 2970 20121 3064 20146
rect 3155 20243 3247 21277
rect 3451 20415 3507 22101
rect 3451 20359 3615 20415
rect 3155 20219 3478 20243
rect 3155 20167 3390 20219
rect 3442 20167 3478 20219
rect 3155 20146 3478 20167
rect 2762 19957 2838 19967
rect 2603 19955 2838 19957
rect 2603 19903 2774 19955
rect 2826 19903 2838 19955
rect 2603 19901 2838 19903
rect 2603 17836 2659 19901
rect 2762 19891 2838 19901
rect 2971 18613 3063 20121
rect 2764 18516 3063 18613
rect 3155 19603 3247 20146
rect 3380 19957 3456 19967
rect 3559 19957 3615 20359
rect 3380 19955 3615 19957
rect 3380 19903 3392 19955
rect 3444 19903 3615 19955
rect 3380 19901 3615 19903
rect 3380 19891 3456 19901
rect 3155 19565 3249 19603
rect 3155 19509 3174 19565
rect 3230 19509 3249 19565
rect 3155 19470 3249 19509
rect 3155 18613 3247 19470
rect 3155 18516 3454 18613
rect 2764 17987 2840 18516
rect 2955 18386 3263 18406
rect 2955 18334 2985 18386
rect 3037 18334 3171 18386
rect 3223 18334 3263 18386
rect 2955 18314 3263 18334
rect 2764 17935 2776 17987
rect 2828 17935 2840 17987
rect 2764 17915 2840 17935
rect 2926 18180 3002 18202
rect 2926 18020 2936 18180
rect 2992 18020 3002 18180
rect 2926 17920 3002 18020
rect 2603 17824 2780 17836
rect 2603 17668 2716 17824
rect 2768 17668 2780 17824
rect 2603 17656 2780 17668
rect 2736 16942 2864 17038
rect 2736 16886 2772 16942
rect 2828 16886 2864 16942
rect 2736 16809 2864 16886
rect 1715 16623 2023 16643
rect 1715 16571 1745 16623
rect 1797 16571 1931 16623
rect 1983 16571 2023 16623
rect 1715 16551 2023 16571
rect 2446 16435 2535 16761
rect 3065 16645 3154 18314
rect 3217 18180 3293 18202
rect 3217 18020 3227 18180
rect 3283 18020 3293 18180
rect 3217 17920 3293 18020
rect 3378 17987 3454 18516
rect 3378 17935 3390 17987
rect 3442 17935 3454 17987
rect 3378 17915 3454 17935
rect 3559 17836 3615 19901
rect 3438 17824 3615 17836
rect 3438 17668 3450 17824
rect 3502 17668 3615 17824
rect 3438 17656 3615 17668
rect 3354 16942 3482 17038
rect 3354 16886 3390 16942
rect 3446 16886 3482 16942
rect 3354 16809 3482 16886
rect 3700 16759 3756 22161
rect 4016 22157 4072 23758
rect 3949 22101 4072 22157
rect 3949 20415 4005 22101
rect 4084 22027 4160 22039
rect 4084 22016 4096 22027
rect 4148 22016 4160 22027
rect 4084 21856 4094 22016
rect 4150 21856 4160 22016
rect 4084 21846 4160 21856
rect 4226 21831 4282 26230
rect 4413 21831 4469 26230
rect 4843 25370 4899 26230
rect 4821 25358 4899 25370
rect 4821 25202 4833 25358
rect 4885 25202 4899 25358
rect 4821 25190 4899 25202
rect 5039 25370 5095 26230
rect 5039 25358 5117 25370
rect 5039 25202 5053 25358
rect 5105 25202 5117 25358
rect 5039 25190 5117 25202
rect 4929 24686 5005 24696
rect 4929 24422 4939 24686
rect 4995 24422 5005 24686
rect 4929 24412 5005 24422
rect 4613 23926 4689 23938
rect 4613 23770 4625 23926
rect 4677 23770 4689 23926
rect 4613 23758 4689 23770
rect 5245 23926 5321 23938
rect 5245 23770 5257 23926
rect 5309 23770 5321 23926
rect 5245 23758 5321 23770
rect 4623 22157 4679 23758
rect 4828 22225 5106 22237
rect 4828 22173 4840 22225
rect 4892 22173 5042 22225
rect 5094 22173 5106 22225
rect 4828 22161 5106 22173
rect 4623 22101 4746 22157
rect 4535 22027 4611 22039
rect 4535 22016 4547 22027
rect 4599 22016 4611 22027
rect 4535 21856 4545 22016
rect 4601 21856 4611 22016
rect 4535 21846 4611 21856
rect 4216 21819 4292 21831
rect 4216 21767 4228 21819
rect 4280 21767 4292 21819
rect 4216 21755 4292 21767
rect 4403 21819 4479 21831
rect 4403 21767 4415 21819
rect 4467 21767 4479 21819
rect 4403 21755 4479 21767
rect 3841 20359 4005 20415
rect 3841 19957 3897 20359
rect 4209 20243 4301 21277
rect 3978 20219 4301 20243
rect 3978 20167 4014 20219
rect 4066 20167 4301 20219
rect 3978 20146 4301 20167
rect 4000 19957 4076 19967
rect 3841 19955 4076 19957
rect 3841 19903 4012 19955
rect 4064 19903 4076 19955
rect 3841 19901 4076 19903
rect 3841 17836 3897 19901
rect 4000 19891 4076 19901
rect 4209 19290 4301 20146
rect 4394 20243 4486 21277
rect 4690 20415 4746 22101
rect 4690 20359 4854 20415
rect 4394 20219 4717 20243
rect 4394 20167 4629 20219
rect 4681 20167 4717 20219
rect 4394 20146 4717 20167
rect 4209 19252 4303 19290
rect 4209 19196 4228 19252
rect 4284 19196 4303 19252
rect 4209 19157 4303 19196
rect 4209 18613 4301 19157
rect 4394 18964 4486 20146
rect 4619 19957 4695 19967
rect 4798 19957 4854 20359
rect 4619 19955 4854 19957
rect 4619 19903 4631 19955
rect 4683 19903 4854 19955
rect 4619 19901 4854 19903
rect 4619 19891 4695 19901
rect 4393 18926 4487 18964
rect 4393 18870 4412 18926
rect 4468 18870 4487 18926
rect 4393 18831 4487 18870
rect 4002 18516 4301 18613
rect 4394 18613 4486 18831
rect 4394 18516 4693 18613
rect 4002 17987 4078 18516
rect 4194 18386 4502 18406
rect 4194 18334 4224 18386
rect 4276 18334 4410 18386
rect 4462 18334 4502 18386
rect 4194 18314 4502 18334
rect 4002 17935 4014 17987
rect 4066 17935 4078 17987
rect 4002 17915 4078 17935
rect 4164 18180 4240 18202
rect 4164 18020 4174 18180
rect 4230 18020 4240 18180
rect 4164 17920 4240 18020
rect 3841 17824 4018 17836
rect 3841 17668 3954 17824
rect 4006 17668 4018 17824
rect 3841 17656 4018 17668
rect 3974 16942 4102 17038
rect 3974 16886 4010 16942
rect 4066 16886 4102 16942
rect 3974 16809 4102 16886
rect 4303 16646 4393 18314
rect 4455 18180 4531 18202
rect 4455 18020 4465 18180
rect 4521 18020 4531 18180
rect 4455 17920 4531 18020
rect 4617 17987 4693 18516
rect 4617 17935 4629 17987
rect 4681 17935 4693 17987
rect 4617 17915 4693 17935
rect 4798 17836 4854 19901
rect 4677 17824 4854 17836
rect 4677 17668 4689 17824
rect 4741 17668 4854 17824
rect 4677 17656 4854 17668
rect 4593 16942 4721 17038
rect 4593 16886 4629 16942
rect 4685 16886 4721 16942
rect 4593 16809 4721 16886
rect 4939 16759 4995 22161
rect 5255 22157 5311 23758
rect 5166 22101 5311 22157
rect 5166 20415 5222 22101
rect 5302 22027 5378 22039
rect 5302 22016 5314 22027
rect 5366 22016 5378 22027
rect 5302 21856 5312 22016
rect 5368 21856 5378 22016
rect 5302 21846 5378 21856
rect 5457 21830 5513 26230
rect 5447 21818 5523 21830
rect 5447 21766 5459 21818
rect 5511 21766 5523 21818
rect 5447 21754 5523 21766
rect 5080 20359 5222 20415
rect 5080 19957 5136 20359
rect 5447 20243 5541 21277
rect 5217 20219 5541 20243
rect 5217 20167 5253 20219
rect 5305 20167 5541 20219
rect 5217 20146 5541 20167
rect 5239 19957 5315 19968
rect 5080 19956 5315 19957
rect 5080 19904 5251 19956
rect 5303 19904 5315 19956
rect 5080 19901 5315 19904
rect 5080 17836 5136 19901
rect 5239 19892 5315 19901
rect 5447 18613 5541 20146
rect 5242 18611 5541 18613
rect 5242 18555 5466 18611
rect 5522 18555 5541 18611
rect 5242 18516 5541 18555
rect 5242 17988 5318 18516
rect 5242 17936 5254 17988
rect 5306 17936 5318 17988
rect 5242 17915 5318 17936
rect 5441 18378 5517 18390
rect 5441 18326 5453 18378
rect 5505 18326 5517 18378
rect 5080 17824 5238 17836
rect 5080 17668 5174 17824
rect 5226 17668 5238 17824
rect 5080 17656 5238 17668
rect 5212 16942 5341 17038
rect 5212 16886 5249 16942
rect 5305 16886 5341 16942
rect 5212 16809 5341 16886
rect 5441 16435 5517 18326
rect 2316 16415 2624 16435
rect 2316 16363 2346 16415
rect 2398 16363 2532 16415
rect 2584 16363 2624 16415
rect 2316 16343 2624 16363
rect 4824 16415 5517 16435
rect 4824 16363 4854 16415
rect 4906 16363 5040 16415
rect 5092 16363 5517 16415
rect 4824 16343 5517 16363
rect 2446 16342 2535 16343
rect 1723 16192 3328 16230
rect 1723 16136 1759 16192
rect 1815 16136 1970 16192
rect 2026 16136 2180 16192
rect 2236 16136 2391 16192
rect 2447 16136 2603 16192
rect 2659 16136 2814 16192
rect 2870 16136 3024 16192
rect 3080 16136 3235 16192
rect 3291 16136 3328 16192
rect 1723 16097 3328 16136
rect 3675 16192 4437 16230
rect 3675 16136 3711 16192
rect 3767 16136 3922 16192
rect 3978 16136 4134 16192
rect 4190 16136 4345 16192
rect 4401 16136 4437 16192
rect 3675 16097 4437 16136
rect 1398 15741 1608 15782
rect 1398 15689 1419 15741
rect 1471 15689 1608 15741
rect 1398 15685 1608 15689
rect 1398 15555 1492 15685
rect 1398 15503 1419 15555
rect 1471 15503 1492 15555
rect 1398 15462 1492 15503
rect 1627 15567 1935 15585
rect 1627 15511 1655 15567
rect 1711 15511 1841 15567
rect 1897 15511 1935 15567
rect 1627 15493 1935 15511
rect 1357 15149 1449 15177
rect 1357 15093 1375 15149
rect 1431 15093 1449 15149
rect 1357 14963 1449 15093
rect 1357 14907 1375 14963
rect 1431 14907 1449 14963
rect 1357 14869 1449 14907
rect 1847 15049 1939 15077
rect 1847 14993 1865 15049
rect 1921 14993 1939 15049
rect 1847 14863 1939 14993
rect 1847 14807 1865 14863
rect 1921 14807 1939 14863
rect 1847 14769 1939 14807
rect 1172 14306 1193 14358
rect 1245 14306 1266 14358
rect 1172 14172 1266 14306
rect 1172 14120 1193 14172
rect 1245 14120 1266 14172
rect 1172 12567 1266 14120
rect 1847 13558 1939 13586
rect 1847 13502 1865 13558
rect 1921 13502 1939 13558
rect 1847 13372 1939 13502
rect 1847 13316 1865 13372
rect 1921 13316 1939 13372
rect 1847 13278 1939 13316
rect 2072 12631 2166 15979
rect 2258 15945 2350 15976
rect 1172 12515 1193 12567
rect 1245 12515 1266 12567
rect 1172 12381 1266 12515
rect 1172 12329 1193 12381
rect 1245 12329 1266 12381
rect 1172 12289 1266 12329
rect 1834 12563 1926 12591
rect 1834 12507 1852 12563
rect 1908 12507 1926 12563
rect 1834 12377 1926 12507
rect 1834 12321 1852 12377
rect 1908 12321 1926 12377
rect 1834 12283 1926 12321
rect 2072 12575 2091 12631
rect 2147 12575 2166 12631
rect 2072 12445 2166 12575
rect 2072 12389 2091 12445
rect 2147 12389 2166 12445
rect 2072 11855 2166 12389
rect 2072 11799 2091 11855
rect 2147 11799 2166 11855
rect 2072 11669 2166 11799
rect 1834 11615 1926 11643
rect 1834 11559 1852 11615
rect 1908 11559 1926 11615
rect 1834 11429 1926 11559
rect 1834 11373 1852 11429
rect 1908 11373 1926 11429
rect 1834 11335 1926 11373
rect 2072 11613 2091 11669
rect 2147 11613 2166 11669
rect 2072 10939 2166 11613
rect 2072 10883 2091 10939
rect 2147 10883 2166 10939
rect 2072 10753 2166 10883
rect 1834 10699 1926 10727
rect 1834 10643 1852 10699
rect 1908 10643 1926 10699
rect 1834 10513 1926 10643
rect 1834 10457 1852 10513
rect 1908 10457 1926 10513
rect 1834 10419 1926 10457
rect 2072 10697 2091 10753
rect 2147 10697 2166 10753
rect 943 10255 1070 10276
rect 2072 10264 2166 10697
rect 2256 15936 2351 15945
rect 2256 15884 2278 15936
rect 2330 15884 2351 15936
rect 2256 15750 2351 15884
rect 2256 15698 2278 15750
rect 2330 15698 2351 15750
rect 943 10203 978 10255
rect 1030 10203 1913 10255
rect 943 10199 1913 10203
rect 943 10183 1070 10199
rect 898 9847 990 9875
rect 898 9791 916 9847
rect 972 9791 990 9847
rect 898 9661 990 9791
rect 1616 9847 1708 9875
rect 1616 9791 1634 9847
rect 1690 9791 1708 9847
rect 898 9605 916 9661
rect 972 9605 990 9661
rect 898 9567 990 9605
rect 1420 9702 1514 9740
rect 1420 9646 1439 9702
rect 1495 9646 1514 9702
rect 258 9527 598 9566
rect 258 9471 294 9527
rect 350 9471 506 9527
rect 562 9471 598 9527
rect 258 9432 598 9471
rect 1420 9516 1514 9646
rect 1616 9661 1708 9791
rect 1616 9605 1634 9661
rect 1690 9605 1708 9661
rect 1616 9567 1708 9605
rect 1420 9460 1439 9516
rect 1495 9460 1514 9516
rect 573 9106 881 9124
rect 573 9050 601 9106
rect 657 9050 787 9106
rect 843 9050 881 9106
rect 573 9032 881 9050
rect 1221 9089 1313 9127
rect 1221 9033 1239 9089
rect 1295 9033 1313 9089
rect 277 8990 369 9018
rect 277 8934 295 8990
rect 351 8934 369 8990
rect 277 8804 369 8934
rect 1221 8903 1313 9033
rect 831 8890 926 8894
rect 277 8748 295 8804
rect 351 8748 369 8804
rect 617 8870 926 8890
rect 617 8818 647 8870
rect 699 8818 833 8870
rect 885 8818 926 8870
rect 1221 8847 1239 8903
rect 1295 8847 1313 8903
rect 1221 8819 1313 8847
rect 617 8798 926 8818
rect 277 8710 369 8748
rect 461 8530 553 8570
rect 461 8478 481 8530
rect 533 8478 553 8530
rect 461 8434 553 8478
rect 460 8344 554 8434
rect 460 8292 481 8344
rect 533 8292 554 8344
rect 460 8 554 8292
rect 831 7826 926 8798
rect 1039 8740 1131 8778
rect 1039 8684 1057 8740
rect 1113 8684 1131 8740
rect 1039 8554 1131 8684
rect 1039 8498 1057 8554
rect 1113 8498 1131 8554
rect 1039 8470 1131 8498
rect 1017 8128 1110 8143
rect 1420 8128 1514 9460
rect 1610 9089 1702 9127
rect 1610 9033 1628 9089
rect 1684 9033 1702 9089
rect 1610 8903 1702 9033
rect 1610 8847 1628 8903
rect 1684 8847 1702 8903
rect 1610 8819 1702 8847
rect 1016 8103 1514 8128
rect 1016 8051 1037 8103
rect 1089 8051 1514 8103
rect 1016 8031 1514 8051
rect 1017 8011 1110 8031
rect 831 7735 1156 7826
rect 1061 5893 1156 7735
rect 1857 7696 1913 10199
rect 2043 9273 2135 9313
rect 2043 9221 2063 9273
rect 2115 9221 2135 9273
rect 2043 9128 2135 9221
rect 2042 9089 2135 9128
rect 2042 9033 2061 9089
rect 2117 9033 2135 9089
rect 2042 8903 2135 9033
rect 2042 8847 2061 8903
rect 2117 8847 2135 8903
rect 2042 8809 2135 8847
rect 1857 7640 2004 7696
rect 845 5795 1156 5893
rect 1508 6367 1602 6374
rect 1508 6327 1603 6367
rect 1508 6275 1531 6327
rect 1583 6275 1603 6327
rect 1508 6141 1603 6275
rect 1508 6089 1531 6141
rect 1583 6089 1603 6141
rect 1508 6049 1603 6089
rect 1948 6083 2004 7640
rect 2256 7648 2351 15698
rect 2441 12631 2535 15979
rect 2441 12575 2460 12631
rect 2516 12575 2535 12631
rect 2441 12445 2535 12575
rect 2441 12389 2460 12445
rect 2516 12389 2535 12445
rect 2441 11855 2535 12389
rect 2441 11799 2460 11855
rect 2516 11799 2535 11855
rect 2441 11669 2535 11799
rect 2441 11613 2460 11669
rect 2516 11613 2535 11669
rect 2441 10939 2535 11613
rect 2441 10883 2460 10939
rect 2516 10883 2535 10939
rect 2441 10753 2535 10883
rect 2441 10697 2460 10753
rect 2516 10697 2535 10753
rect 2441 10264 2535 10697
rect 5345 10246 5437 10286
rect 5345 10198 5365 10246
rect 5344 10194 5365 10198
rect 5417 10198 5437 10246
rect 5417 10194 5438 10198
rect 5344 10060 5438 10194
rect 5344 10008 5365 10060
rect 5417 10008 5438 10060
rect 2772 9942 2864 9970
rect 2772 9886 2790 9942
rect 2846 9886 2864 9942
rect 2772 9756 2864 9886
rect 2772 9700 2790 9756
rect 2846 9700 2864 9756
rect 2772 9662 2864 9700
rect 2772 9019 2864 9047
rect 2772 8963 2790 9019
rect 2846 8963 2864 9019
rect 2772 8833 2864 8963
rect 2772 8777 2790 8833
rect 2846 8777 2864 8833
rect 2772 8739 2864 8777
rect 4233 8346 4327 8525
rect 4692 8467 4786 8646
rect 4692 8370 5050 8467
rect 4233 8249 4435 8346
rect 4956 8229 5050 8370
rect 2256 7566 2859 7648
rect 845 1465 940 5795
rect 1508 5771 1602 6049
rect 1308 5647 1602 5771
rect 1877 6027 2004 6083
rect 845 1287 958 1465
rect 878 -82 958 1287
rect 1308 -1 1402 5647
rect 1877 1860 1933 6027
rect 2298 5006 2354 5866
rect 2764 5052 2859 7566
rect 4395 5916 4715 6050
rect 5344 6002 5438 10008
rect 4639 5597 4715 5916
rect 4639 5441 4651 5597
rect 4703 5441 4715 5597
rect 4639 5429 4715 5441
rect 5125 5905 5438 6002
rect 5125 5597 5201 5905
rect 5125 5441 5137 5597
rect 5189 5441 5201 5597
rect 5125 5429 5201 5441
rect 2131 4996 2354 5006
rect 2131 4940 2141 4996
rect 2301 4940 2354 4996
rect 2480 4974 2859 5052
rect 2131 4930 2311 4940
rect 2480 4655 2575 4974
rect 2256 4533 2575 4655
rect 2256 3610 2351 4533
rect 2256 3558 2277 3610
rect 2329 3558 2351 3610
rect 2256 3424 2351 3558
rect 2256 3372 2277 3424
rect 2329 3372 2351 3424
rect 2256 3331 2351 3372
rect 1877 1804 1984 1860
rect 1928 993 1984 1804
rect 1928 917 2054 993
rect 828 -94 1008 -82
rect 828 -146 840 -94
rect 996 -146 1008 -94
rect 828 -158 1008 -146
rect 1998 -1900 2054 917
rect 5547 558 5623 568
rect 5547 190 5557 558
rect 5613 190 5623 558
rect 5547 180 5623 190
rect 1998 -1956 3066 -1900
rect 3010 -2247 3066 -1956
rect 3000 -2259 3076 -2247
rect 3000 -2415 3012 -2259
rect 3064 -2415 3076 -2259
rect 3000 -2427 3076 -2415
<< via2 >>
rect 916 28963 972 28965
rect 916 28911 918 28963
rect 918 28911 970 28963
rect 970 28911 972 28963
rect 916 28909 972 28911
rect 916 28777 972 28779
rect 916 28725 918 28777
rect 918 28725 970 28777
rect 970 28725 972 28777
rect 916 28723 972 28725
rect 1530 28963 1586 28965
rect 1530 28911 1532 28963
rect 1532 28911 1584 28963
rect 1584 28911 1586 28963
rect 1530 28909 1586 28911
rect 1530 28777 1586 28779
rect 1530 28725 1532 28777
rect 1532 28725 1584 28777
rect 1584 28725 1586 28777
rect 1530 28723 1586 28725
rect 2155 28963 2211 28965
rect 2155 28911 2157 28963
rect 2157 28911 2209 28963
rect 2209 28911 2211 28963
rect 2155 28909 2211 28911
rect 2155 28777 2211 28779
rect 2155 28725 2157 28777
rect 2157 28725 2209 28777
rect 2209 28725 2211 28777
rect 2155 28723 2211 28725
rect 2769 28963 2825 28965
rect 2769 28911 2771 28963
rect 2771 28911 2823 28963
rect 2823 28911 2825 28963
rect 2769 28909 2825 28911
rect 2769 28777 2825 28779
rect 2769 28725 2771 28777
rect 2771 28725 2823 28777
rect 2823 28725 2825 28777
rect 2769 28723 2825 28725
rect 3393 28963 3449 28965
rect 3393 28911 3395 28963
rect 3395 28911 3447 28963
rect 3447 28911 3449 28963
rect 3393 28909 3449 28911
rect 3393 28777 3449 28779
rect 3393 28725 3395 28777
rect 3395 28725 3447 28777
rect 3447 28725 3449 28777
rect 3393 28723 3449 28725
rect 4007 28963 4063 28965
rect 4007 28911 4009 28963
rect 4009 28911 4061 28963
rect 4061 28911 4063 28963
rect 4007 28909 4063 28911
rect 4007 28777 4063 28779
rect 4007 28725 4009 28777
rect 4009 28725 4061 28777
rect 4061 28725 4063 28777
rect 4007 28723 4063 28725
rect 4632 28963 4688 28965
rect 4632 28911 4634 28963
rect 4634 28911 4686 28963
rect 4686 28911 4688 28963
rect 4632 28909 4688 28911
rect 4632 28777 4688 28779
rect 4632 28725 4634 28777
rect 4634 28725 4686 28777
rect 4686 28725 4688 28777
rect 4632 28723 4688 28725
rect 5246 28963 5302 28965
rect 5246 28911 5248 28963
rect 5248 28911 5300 28963
rect 5300 28911 5302 28963
rect 5246 28909 5302 28911
rect 5246 28777 5302 28779
rect 5246 28725 5248 28777
rect 5248 28725 5300 28777
rect 5300 28725 5302 28777
rect 5246 28723 5302 28725
rect 1223 24684 1279 24686
rect 1223 24424 1225 24684
rect 1225 24424 1277 24684
rect 1277 24424 1279 24684
rect 1223 24422 1279 24424
rect 829 21975 831 22016
rect 831 21975 883 22016
rect 883 21975 885 22016
rect 829 21856 885 21975
rect 697 21130 753 21186
rect 913 16940 969 16942
rect 913 16888 915 16940
rect 915 16888 967 16940
rect 967 16888 969 16940
rect 913 16886 969 16888
rect 1617 21975 1619 22016
rect 1619 21975 1671 22016
rect 1671 21975 1673 22016
rect 1617 21856 1673 21975
rect 2462 24684 2518 24686
rect 2462 24424 2464 24684
rect 2464 24424 2516 24684
rect 2516 24424 2518 24684
rect 2462 24422 2518 24424
rect 2068 21975 2070 22016
rect 2070 21975 2122 22016
rect 2122 21975 2124 22016
rect 2068 21856 2124 21975
rect 1751 20811 1807 20867
rect 1935 20482 1991 20538
rect 1697 18178 1753 18180
rect 1697 18126 1699 18178
rect 1699 18126 1751 18178
rect 1751 18126 1753 18178
rect 1697 18020 1753 18126
rect 1533 16940 1589 16942
rect 1533 16888 1535 16940
rect 1535 16888 1587 16940
rect 1587 16888 1589 16940
rect 1533 16886 1589 16888
rect 295 15612 351 15614
rect 295 15560 297 15612
rect 297 15560 349 15612
rect 349 15560 351 15612
rect 295 15558 351 15560
rect 295 15426 351 15428
rect 295 15374 297 15426
rect 297 15374 349 15426
rect 349 15374 351 15426
rect 295 15372 351 15374
rect 295 15013 351 15015
rect 295 14961 297 15013
rect 297 14961 349 15013
rect 349 14961 351 15013
rect 295 14959 351 14961
rect 295 14827 351 14829
rect 295 14775 297 14827
rect 297 14775 349 14827
rect 349 14775 351 14827
rect 295 14773 351 14775
rect 965 16190 1021 16192
rect 965 16138 967 16190
rect 967 16138 1019 16190
rect 1019 16138 1021 16190
rect 965 16136 1021 16138
rect 295 13556 351 13558
rect 295 13504 297 13556
rect 297 13504 349 13556
rect 349 13504 351 13556
rect 295 13502 351 13504
rect 295 13370 351 13372
rect 295 13318 297 13370
rect 297 13318 349 13370
rect 349 13318 351 13370
rect 295 13316 351 13318
rect 295 12561 351 12563
rect 295 12509 297 12561
rect 297 12509 349 12561
rect 349 12509 351 12561
rect 295 12507 351 12509
rect 295 12375 351 12377
rect 295 12323 297 12375
rect 297 12323 349 12375
rect 349 12323 351 12375
rect 295 12321 351 12323
rect 295 11613 351 11615
rect 295 11561 297 11613
rect 297 11561 349 11613
rect 349 11561 351 11613
rect 295 11559 351 11561
rect 295 11427 351 11429
rect 295 11375 297 11427
rect 297 11375 349 11427
rect 349 11375 351 11427
rect 295 11373 351 11375
rect 295 10697 351 10699
rect 295 10645 297 10697
rect 297 10645 349 10697
rect 349 10645 351 10697
rect 295 10643 351 10645
rect 295 10511 351 10513
rect 295 10459 297 10511
rect 297 10459 349 10511
rect 349 10459 351 10511
rect 295 10457 351 10459
rect 1988 18178 2044 18180
rect 1988 18126 1990 18178
rect 1990 18126 2042 18178
rect 2042 18126 2044 18178
rect 1988 18020 2044 18126
rect 2152 16940 2208 16942
rect 2152 16888 2154 16940
rect 2154 16888 2206 16940
rect 2206 16888 2208 16940
rect 2152 16886 2208 16888
rect 2856 21975 2858 22016
rect 2858 21975 2910 22016
rect 2910 21975 2912 22016
rect 2856 21856 2912 21975
rect 3700 24684 3756 24686
rect 3700 24424 3702 24684
rect 3702 24424 3754 24684
rect 3754 24424 3756 24684
rect 3700 24422 3756 24424
rect 3306 21975 3308 22016
rect 3308 21975 3360 22016
rect 3360 21975 3362 22016
rect 3306 21856 3362 21975
rect 2989 20160 3045 20216
rect 3174 19509 3230 19565
rect 2936 18178 2992 18180
rect 2936 18126 2938 18178
rect 2938 18126 2990 18178
rect 2990 18126 2992 18178
rect 2936 18020 2992 18126
rect 2772 16940 2828 16942
rect 2772 16888 2774 16940
rect 2774 16888 2826 16940
rect 2826 16888 2828 16940
rect 2772 16886 2828 16888
rect 3227 18178 3283 18180
rect 3227 18126 3229 18178
rect 3229 18126 3281 18178
rect 3281 18126 3283 18178
rect 3227 18020 3283 18126
rect 3390 16940 3446 16942
rect 3390 16888 3392 16940
rect 3392 16888 3444 16940
rect 3444 16888 3446 16940
rect 3390 16886 3446 16888
rect 4094 21975 4096 22016
rect 4096 21975 4148 22016
rect 4148 21975 4150 22016
rect 4094 21856 4150 21975
rect 4939 24684 4995 24686
rect 4939 24424 4941 24684
rect 4941 24424 4993 24684
rect 4993 24424 4995 24684
rect 4939 24422 4995 24424
rect 4545 21975 4547 22016
rect 4547 21975 4599 22016
rect 4599 21975 4601 22016
rect 4545 21856 4601 21975
rect 4228 19196 4284 19252
rect 4412 18870 4468 18926
rect 4174 18178 4230 18180
rect 4174 18126 4176 18178
rect 4176 18126 4228 18178
rect 4228 18126 4230 18178
rect 4174 18020 4230 18126
rect 4010 16940 4066 16942
rect 4010 16888 4012 16940
rect 4012 16888 4064 16940
rect 4064 16888 4066 16940
rect 4010 16886 4066 16888
rect 4465 18178 4521 18180
rect 4465 18126 4467 18178
rect 4467 18126 4519 18178
rect 4519 18126 4521 18178
rect 4465 18020 4521 18126
rect 4629 16940 4685 16942
rect 4629 16888 4631 16940
rect 4631 16888 4683 16940
rect 4683 16888 4685 16940
rect 4629 16886 4685 16888
rect 5312 21975 5314 22016
rect 5314 21975 5366 22016
rect 5366 21975 5368 22016
rect 5312 21856 5368 21975
rect 5466 18555 5522 18611
rect 5249 16940 5305 16942
rect 5249 16888 5251 16940
rect 5251 16888 5303 16940
rect 5303 16888 5305 16940
rect 5249 16886 5305 16888
rect 1759 16190 1815 16192
rect 1759 16138 1761 16190
rect 1761 16138 1813 16190
rect 1813 16138 1815 16190
rect 1759 16136 1815 16138
rect 1970 16190 2026 16192
rect 1970 16138 1972 16190
rect 1972 16138 2024 16190
rect 2024 16138 2026 16190
rect 1970 16136 2026 16138
rect 2180 16190 2236 16192
rect 2180 16138 2182 16190
rect 2182 16138 2234 16190
rect 2234 16138 2236 16190
rect 2180 16136 2236 16138
rect 2391 16190 2447 16192
rect 2391 16138 2393 16190
rect 2393 16138 2445 16190
rect 2445 16138 2447 16190
rect 2391 16136 2447 16138
rect 2603 16190 2659 16192
rect 2603 16138 2605 16190
rect 2605 16138 2657 16190
rect 2657 16138 2659 16190
rect 2603 16136 2659 16138
rect 2814 16190 2870 16192
rect 2814 16138 2816 16190
rect 2816 16138 2868 16190
rect 2868 16138 2870 16190
rect 2814 16136 2870 16138
rect 3024 16190 3080 16192
rect 3024 16138 3026 16190
rect 3026 16138 3078 16190
rect 3078 16138 3080 16190
rect 3024 16136 3080 16138
rect 3235 16190 3291 16192
rect 3235 16138 3237 16190
rect 3237 16138 3289 16190
rect 3289 16138 3291 16190
rect 3235 16136 3291 16138
rect 3711 16190 3767 16192
rect 3711 16138 3713 16190
rect 3713 16138 3765 16190
rect 3765 16138 3767 16190
rect 3711 16136 3767 16138
rect 3922 16190 3978 16192
rect 3922 16138 3924 16190
rect 3924 16138 3976 16190
rect 3976 16138 3978 16190
rect 3922 16136 3978 16138
rect 4134 16190 4190 16192
rect 4134 16138 4136 16190
rect 4136 16138 4188 16190
rect 4188 16138 4190 16190
rect 4134 16136 4190 16138
rect 4345 16190 4401 16192
rect 4345 16138 4347 16190
rect 4347 16138 4399 16190
rect 4399 16138 4401 16190
rect 4345 16136 4401 16138
rect 1655 15565 1711 15567
rect 1655 15513 1657 15565
rect 1657 15513 1709 15565
rect 1709 15513 1711 15565
rect 1655 15511 1711 15513
rect 1841 15565 1897 15567
rect 1841 15513 1843 15565
rect 1843 15513 1895 15565
rect 1895 15513 1897 15565
rect 1841 15511 1897 15513
rect 1375 15147 1431 15149
rect 1375 15095 1377 15147
rect 1377 15095 1429 15147
rect 1429 15095 1431 15147
rect 1375 15093 1431 15095
rect 1375 14961 1431 14963
rect 1375 14909 1377 14961
rect 1377 14909 1429 14961
rect 1429 14909 1431 14961
rect 1375 14907 1431 14909
rect 1865 15047 1921 15049
rect 1865 14995 1867 15047
rect 1867 14995 1919 15047
rect 1919 14995 1921 15047
rect 1865 14993 1921 14995
rect 1865 14861 1921 14863
rect 1865 14809 1867 14861
rect 1867 14809 1919 14861
rect 1919 14809 1921 14861
rect 1865 14807 1921 14809
rect 1865 13556 1921 13558
rect 1865 13504 1867 13556
rect 1867 13504 1919 13556
rect 1919 13504 1921 13556
rect 1865 13502 1921 13504
rect 1865 13370 1921 13372
rect 1865 13318 1867 13370
rect 1867 13318 1919 13370
rect 1919 13318 1921 13370
rect 1865 13316 1921 13318
rect 1852 12561 1908 12563
rect 1852 12509 1854 12561
rect 1854 12509 1906 12561
rect 1906 12509 1908 12561
rect 1852 12507 1908 12509
rect 1852 12375 1908 12377
rect 1852 12323 1854 12375
rect 1854 12323 1906 12375
rect 1906 12323 1908 12375
rect 1852 12321 1908 12323
rect 2091 12629 2147 12631
rect 2091 12577 2093 12629
rect 2093 12577 2145 12629
rect 2145 12577 2147 12629
rect 2091 12575 2147 12577
rect 2091 12443 2147 12445
rect 2091 12391 2093 12443
rect 2093 12391 2145 12443
rect 2145 12391 2147 12443
rect 2091 12389 2147 12391
rect 2091 11853 2147 11855
rect 2091 11801 2093 11853
rect 2093 11801 2145 11853
rect 2145 11801 2147 11853
rect 2091 11799 2147 11801
rect 1852 11613 1908 11615
rect 1852 11561 1854 11613
rect 1854 11561 1906 11613
rect 1906 11561 1908 11613
rect 1852 11559 1908 11561
rect 1852 11427 1908 11429
rect 1852 11375 1854 11427
rect 1854 11375 1906 11427
rect 1906 11375 1908 11427
rect 1852 11373 1908 11375
rect 2091 11667 2147 11669
rect 2091 11615 2093 11667
rect 2093 11615 2145 11667
rect 2145 11615 2147 11667
rect 2091 11613 2147 11615
rect 2091 10937 2147 10939
rect 2091 10885 2093 10937
rect 2093 10885 2145 10937
rect 2145 10885 2147 10937
rect 2091 10883 2147 10885
rect 1852 10697 1908 10699
rect 1852 10645 1854 10697
rect 1854 10645 1906 10697
rect 1906 10645 1908 10697
rect 1852 10643 1908 10645
rect 1852 10511 1908 10513
rect 1852 10459 1854 10511
rect 1854 10459 1906 10511
rect 1906 10459 1908 10511
rect 1852 10457 1908 10459
rect 2091 10751 2147 10753
rect 2091 10699 2093 10751
rect 2093 10699 2145 10751
rect 2145 10699 2147 10751
rect 2091 10697 2147 10699
rect 916 9845 972 9847
rect 916 9793 918 9845
rect 918 9793 970 9845
rect 970 9793 972 9845
rect 916 9791 972 9793
rect 1634 9845 1690 9847
rect 1634 9793 1636 9845
rect 1636 9793 1688 9845
rect 1688 9793 1690 9845
rect 1634 9791 1690 9793
rect 916 9659 972 9661
rect 916 9607 918 9659
rect 918 9607 970 9659
rect 970 9607 972 9659
rect 916 9605 972 9607
rect 1439 9646 1495 9702
rect 294 9525 350 9527
rect 294 9473 296 9525
rect 296 9473 348 9525
rect 348 9473 350 9525
rect 294 9471 350 9473
rect 506 9525 562 9527
rect 506 9473 508 9525
rect 508 9473 560 9525
rect 560 9473 562 9525
rect 506 9471 562 9473
rect 1634 9659 1690 9661
rect 1634 9607 1636 9659
rect 1636 9607 1688 9659
rect 1688 9607 1690 9659
rect 1634 9605 1690 9607
rect 1439 9460 1495 9516
rect 601 9104 657 9106
rect 601 9052 603 9104
rect 603 9052 655 9104
rect 655 9052 657 9104
rect 601 9050 657 9052
rect 787 9104 843 9106
rect 787 9052 789 9104
rect 789 9052 841 9104
rect 841 9052 843 9104
rect 787 9050 843 9052
rect 1239 9087 1295 9089
rect 1239 9035 1241 9087
rect 1241 9035 1293 9087
rect 1293 9035 1295 9087
rect 1239 9033 1295 9035
rect 295 8988 351 8990
rect 295 8936 297 8988
rect 297 8936 349 8988
rect 349 8936 351 8988
rect 295 8934 351 8936
rect 295 8802 351 8804
rect 295 8750 297 8802
rect 297 8750 349 8802
rect 349 8750 351 8802
rect 295 8748 351 8750
rect 1239 8901 1295 8903
rect 1239 8849 1241 8901
rect 1241 8849 1293 8901
rect 1293 8849 1295 8901
rect 1239 8847 1295 8849
rect 1057 8738 1113 8740
rect 1057 8686 1059 8738
rect 1059 8686 1111 8738
rect 1111 8686 1113 8738
rect 1057 8684 1113 8686
rect 1057 8552 1113 8554
rect 1057 8500 1059 8552
rect 1059 8500 1111 8552
rect 1111 8500 1113 8552
rect 1057 8498 1113 8500
rect 1628 9087 1684 9089
rect 1628 9035 1630 9087
rect 1630 9035 1682 9087
rect 1682 9035 1684 9087
rect 1628 9033 1684 9035
rect 1628 8901 1684 8903
rect 1628 8849 1630 8901
rect 1630 8849 1682 8901
rect 1682 8849 1684 8901
rect 1628 8847 1684 8849
rect 2061 9087 2117 9089
rect 2061 9035 2063 9087
rect 2063 9035 2115 9087
rect 2115 9035 2117 9087
rect 2061 9033 2117 9035
rect 2061 8847 2117 8903
rect 2460 12575 2516 12631
rect 2460 12389 2516 12445
rect 2460 11799 2516 11855
rect 2460 11613 2516 11669
rect 2460 10883 2516 10939
rect 2460 10697 2516 10753
rect 2790 9940 2846 9942
rect 2790 9888 2792 9940
rect 2792 9888 2844 9940
rect 2844 9888 2846 9940
rect 2790 9886 2846 9888
rect 2790 9754 2846 9756
rect 2790 9702 2792 9754
rect 2792 9702 2844 9754
rect 2844 9702 2846 9754
rect 2790 9700 2846 9702
rect 2790 9017 2846 9019
rect 2790 8965 2792 9017
rect 2792 8965 2844 9017
rect 2844 8965 2846 9017
rect 2790 8963 2846 8965
rect 2790 8831 2846 8833
rect 2790 8779 2792 8831
rect 2792 8779 2844 8831
rect 2844 8779 2846 8831
rect 2790 8777 2846 8779
rect 2141 4940 2301 4996
rect 5557 556 5613 558
rect 5557 192 5559 556
rect 5559 192 5611 556
rect 5611 192 5613 556
rect 5557 190 5613 192
<< metal3 >>
rect 322 28965 5618 29107
rect 322 28909 916 28965
rect 972 28909 1530 28965
rect 1586 28909 2155 28965
rect 2211 28909 2769 28965
rect 2825 28909 3393 28965
rect 3449 28909 4007 28965
rect 4063 28909 4632 28965
rect 4688 28909 5246 28965
rect 5302 28909 5618 28965
rect 322 28779 5618 28909
rect 322 28723 916 28779
rect 972 28723 1530 28779
rect 1586 28723 2155 28779
rect 2211 28723 2769 28779
rect 2825 28723 3393 28779
rect 3449 28723 4007 28779
rect 4063 28723 4632 28779
rect 4688 28723 5246 28779
rect 5302 28723 5618 28779
rect 322 27298 5618 28723
rect -269 24686 7633 24696
rect -269 24422 1223 24686
rect 1279 24422 2462 24686
rect 2518 24422 3700 24686
rect 3756 24422 4939 24686
rect 4995 24422 7633 24686
rect -269 24412 7633 24422
rect -1 22016 5603 23398
rect -1 21856 829 22016
rect 885 21856 1617 22016
rect 1673 21856 2068 22016
rect 2124 21856 2856 22016
rect 2912 21856 3306 22016
rect 3362 21856 4094 22016
rect 4150 21856 4545 22016
rect 4601 21856 5312 22016
rect 5368 21856 5603 22016
rect -1 21417 5603 21856
rect 4966 21416 5603 21417
rect 322 21186 5603 21306
rect 322 21130 697 21186
rect 753 21130 5603 21186
rect 322 21091 5603 21130
rect 322 20867 5603 20984
rect 322 20811 1751 20867
rect 1807 20811 5603 20867
rect 322 20769 5603 20811
rect 322 20538 5603 20663
rect 322 20482 1935 20538
rect 1991 20482 5603 20538
rect 322 20448 5603 20482
rect 1916 20443 2010 20448
rect 322 20216 5603 20341
rect 322 20160 2989 20216
rect 3045 20160 5603 20216
rect 322 20126 5603 20160
rect 2970 20121 3064 20126
rect 322 19565 5603 19649
rect 322 19509 3174 19565
rect 3230 19509 5603 19565
rect 322 19434 5603 19509
rect 322 19252 5603 19327
rect 322 19196 4228 19252
rect 4284 19196 5603 19252
rect 322 19112 5603 19196
rect 322 18926 5603 19005
rect 322 18870 4412 18926
rect 4468 18870 5603 18926
rect 322 18790 5603 18870
rect 322 18611 5603 18683
rect 322 18555 5466 18611
rect 5522 18555 5603 18611
rect 322 18468 5603 18555
rect 322 18180 5603 18362
rect 322 18020 1697 18180
rect 1753 18020 1988 18180
rect 2044 18020 2936 18180
rect 2992 18020 3227 18180
rect 3283 18020 4174 18180
rect 4230 18020 4465 18180
rect 4521 18020 5603 18180
rect 322 17920 5603 18020
rect 322 16942 5603 17264
rect 322 16886 913 16942
rect 969 16886 1533 16942
rect 1589 16886 2152 16942
rect 2208 16886 2772 16942
rect 2828 16886 3390 16942
rect 3446 16886 4010 16942
rect 4066 16886 4629 16942
rect 4685 16886 5249 16942
rect 5305 16886 5603 16942
rect 322 16809 5603 16886
rect 377 16192 5517 16235
rect 377 16136 965 16192
rect 1021 16136 1759 16192
rect 1815 16136 1970 16192
rect 2026 16136 2180 16192
rect 2236 16136 2391 16192
rect 2447 16136 2603 16192
rect 2659 16136 2814 16192
rect 2870 16136 3024 16192
rect 3080 16136 3235 16192
rect 3291 16136 3711 16192
rect 3767 16136 3922 16192
rect 3978 16136 4134 16192
rect 4190 16136 4345 16192
rect 4401 16136 5517 16192
rect 377 16006 5517 16136
rect 276 15614 2779 15720
rect 276 15558 295 15614
rect 351 15567 2779 15614
rect 351 15558 1655 15567
rect 276 15511 1655 15558
rect 1711 15511 1841 15567
rect 1897 15511 2779 15567
rect 276 15428 2779 15511
rect 276 15372 295 15428
rect 351 15372 2779 15428
rect 276 15149 2779 15372
rect 276 15093 1375 15149
rect 1431 15093 2779 15149
rect 276 15049 2779 15093
rect 276 15015 1865 15049
rect 276 14959 295 15015
rect 351 14993 1865 15015
rect 1921 14993 2779 15049
rect 351 14963 2779 14993
rect 351 14959 1375 14963
rect 276 14907 1375 14959
rect 1431 14907 2779 14963
rect 276 14863 2779 14907
rect 276 14829 1865 14863
rect 276 14773 295 14829
rect 351 14807 1865 14829
rect 1921 14807 2779 14863
rect 351 14773 2779 14807
rect 276 13558 2779 14773
rect 276 13502 295 13558
rect 351 13502 1865 13558
rect 1921 13502 2779 13558
rect 276 13372 2779 13502
rect 276 13316 295 13372
rect 351 13316 1865 13372
rect 1921 13316 2779 13372
rect 276 12998 2779 13316
rect 5493 12998 5794 15720
rect 276 12631 2779 12712
rect 276 12575 2091 12631
rect 2147 12575 2460 12631
rect 2516 12575 2779 12631
rect 276 12563 2779 12575
rect 276 12507 295 12563
rect 351 12507 1852 12563
rect 1908 12507 2779 12563
rect 276 12445 2779 12507
rect 276 12389 2091 12445
rect 2147 12389 2460 12445
rect 2516 12389 2779 12445
rect 276 12377 2779 12389
rect 276 12321 295 12377
rect 351 12321 1852 12377
rect 1908 12321 2779 12377
rect 276 11855 2779 12321
rect 276 11799 2091 11855
rect 2147 11799 2460 11855
rect 2516 11799 2779 11855
rect 276 11669 2779 11799
rect 276 11615 2091 11669
rect 276 11559 295 11615
rect 351 11559 1852 11615
rect 1908 11613 2091 11615
rect 2147 11613 2460 11669
rect 2516 11613 2779 11669
rect 1908 11559 2779 11613
rect 276 11429 2779 11559
rect 276 11373 295 11429
rect 351 11373 1852 11429
rect 1908 11373 2779 11429
rect 276 10939 2779 11373
rect 276 10883 2091 10939
rect 2147 10883 2460 10939
rect 2516 10883 2779 10939
rect 276 10753 2779 10883
rect 276 10699 2091 10753
rect 276 10643 295 10699
rect 351 10643 1852 10699
rect 1908 10697 2091 10699
rect 2147 10697 2460 10753
rect 2516 10697 2779 10753
rect 1908 10643 2779 10697
rect 276 10513 2779 10643
rect 276 10457 295 10513
rect 351 10457 1852 10513
rect 1908 10457 2779 10513
rect 276 9970 2779 10457
rect 276 9942 2865 9970
rect 276 9886 2790 9942
rect 2846 9886 2865 9942
rect 276 9847 2865 9886
rect 276 9791 916 9847
rect 972 9791 1634 9847
rect 1690 9791 2865 9847
rect 276 9756 2865 9791
rect 276 9702 2790 9756
rect 276 9661 1439 9702
rect 276 9605 916 9661
rect 972 9646 1439 9661
rect 1495 9700 2790 9702
rect 2846 9700 2865 9756
rect 1495 9661 2865 9700
rect 1495 9646 1634 9661
rect 972 9605 1634 9646
rect 1690 9605 2779 9661
rect 276 9566 2779 9605
rect 258 9527 2779 9566
rect 258 9471 294 9527
rect 350 9471 506 9527
rect 562 9516 2779 9527
rect 562 9471 1439 9516
rect 258 9460 1439 9471
rect 1495 9460 2779 9516
rect 258 9432 2779 9460
rect 276 9310 2779 9432
rect 276 9106 2779 9160
rect 276 9050 601 9106
rect 657 9050 787 9106
rect 843 9089 2779 9106
rect 843 9050 1239 9089
rect 276 9033 1239 9050
rect 1295 9033 1628 9089
rect 1684 9033 2061 9089
rect 2117 9047 2779 9089
rect 2117 9033 2865 9047
rect 276 9019 2865 9033
rect 276 8990 2790 9019
rect 276 8934 295 8990
rect 351 8963 2790 8990
rect 2846 8963 2865 9019
rect 351 8934 2865 8963
rect 276 8903 2865 8934
rect 276 8847 1239 8903
rect 1295 8847 1628 8903
rect 1684 8847 2061 8903
rect 2117 8847 2865 8903
rect 276 8833 2865 8847
rect 276 8804 2790 8833
rect 276 8748 295 8804
rect 351 8777 2790 8804
rect 2846 8777 2865 8833
rect 351 8748 2865 8777
rect 276 8740 2865 8748
rect 276 8684 1057 8740
rect 1113 8738 2865 8740
rect 1113 8684 2779 8738
rect 276 8554 2779 8684
rect 276 8498 1057 8554
rect 1113 8498 2779 8554
rect 276 8443 2779 8498
rect 318 4996 2311 5012
rect 318 4940 2141 4996
rect 2301 4940 2311 4996
rect 318 4924 2311 4940
rect 5627 3135 5794 4496
rect 5547 558 5623 568
rect 5547 190 5557 558
rect 5613 190 5623 558
rect 5547 180 5623 190
rect 5636 156 5794 611
use din_128x8m81  din_128x8m81_0
timestamp 1755005639
transform 1 0 323 0 1 7812
box -46 -15 2450 8740
use M1_NACTIVE4310590548725_128x8m81  M1_NACTIVE4310590548725_128x8m81_0
timestamp 1755005639
transform 1 0 5585 0 1 372
box 0 0 1 1
use M2_M1$$45012012_128x8m81  M2_M1$$45012012_128x8m81_0
timestamp 1755005639
transform 1 0 2525 0 1 16164
box 0 0 1 1
use M2_M1$$45013036_128x8m81  M2_M1$$45013036_128x8m81_0
timestamp 1755005639
transform 1 0 4056 0 1 16164
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_0
timestamp 1755005639
transform 0 -1 5163 1 0 5519
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_1
timestamp 1755005639
transform 0 -1 4677 1 0 5519
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_0
timestamp 1755005639
transform 0 -1 918 1 0 -120
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_1
timestamp 1755005639
transform 1 0 3038 0 1 -2337
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_0
timestamp 1755005639
transform 1 0 525 0 1 27067
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_1
timestamp 1755005639
transform 1 0 740 0 1 18352
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_2
timestamp 1755005639
transform 1 0 5479 0 1 18352
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_3
timestamp 1755005639
transform 1 0 525 0 1 15927
box 0 0 1 1
use M2_M14310590548726_128x8m81  M2_M14310590548726_128x8m81_0
timestamp 1755005639
transform 1 0 5585 0 1 374
box 0 0 1 1
use m2_saout01_128x8m81  m2_saout01_128x8m81_0
timestamp 1755005639
transform 1 0 686 0 1 28987
box -89 -63 4849 2153
use M3_M2$$43370540_128x8m81  M3_M2$$43370540_128x8m81_0
timestamp 1755005639
transform 1 0 4056 0 1 16164
box 0 0 1 1
use M3_M2$$44741676_128x8m81  M3_M2$$44741676_128x8m81_0
timestamp 1755005639
transform 1 0 2525 0 1 16164
box 0 0 1 1
use M3_M2431059054874_128x8m81  M3_M2431059054874_128x8m81_0
timestamp 1755005639
transform 1 0 2221 0 1 4968
box 0 0 1 1
use M3_M24310590548727_128x8m81  M3_M24310590548727_128x8m81_0
timestamp 1755005639
transform 1 0 5585 0 1 374
box 0 0 1 1
use mux821_128x8m81  mux821_128x8m81_0
timestamp 1755005639
transform 1 0 553 0 1 16669
box -9 164 5035 12234
use outbuf_oe_128x8m81  outbuf_oe_128x8m81_0
timestamp 1755005639
transform 1 0 632 0 1 5516
box -532 -359 5177 3324
use sa_128x8m81  sa_128x8m81_0
timestamp 1755005639
transform 1 0 632 0 1 8615
box -357 -196 5034 8146
use sacntl_2_128x8m81  sacntl_2_128x8m81_0
timestamp 1755005639
transform 1 0 632 0 1 30
box -530 -24 5176 5655
use via1_2_x2_128x8m81  via1_2_x2_128x8m81_0
timestamp 1755005639
transform 1 0 2073 0 1 12351
box 0 0 1 1
use via1_2_x2_128x8m81  via1_2_x2_128x8m81_1
timestamp 1755005639
transform 1 0 2073 0 1 11575
box 0 0 1 1
use via1_2_x2_128x8m81  via1_2_x2_128x8m81_2
timestamp 1755005639
transform 1 0 2073 0 1 10659
box 0 0 1 1
use via1_x2_128x8m81  via1_x2_128x8m81_0
timestamp 1755005639
transform -1 0 2350 0 -1 15976
box 0 0 1 1
use via1_x2_128x8m81  via1_x2_128x8m81_1
timestamp 1755005639
transform -1 0 1603 0 -1 6367
box 0 0 1 1
use via1_x2_128x8m81  via1_x2_128x8m81_2
timestamp 1755005639
transform 1 0 2257 0 1 3332
box 0 0 1 1
use via1_x2_128x8m81  via1_x2_128x8m81_3
timestamp 1755005639
transform 1 0 5345 0 1 9968
box 0 0 1 1
use via1_x2_128x8m81  via1_x2_128x8m81_4
timestamp 1755005639
transform 1 0 461 0 1 8252
box 0 0 1 1
use via1_x2_R90_128x8m81  via1_x2_R90_128x8m81_0
timestamp 1755005639
transform 0 -1 5132 1 0 16343
box 0 0 1 1
use via1_x2_R90_128x8m81  via1_x2_R90_128x8m81_1
timestamp 1755005639
transform 0 -1 2025 1 0 18314
box 0 0 1 1
use via1_x2_R90_128x8m81  via1_x2_R90_128x8m81_2
timestamp 1755005639
transform 0 -1 3263 1 0 18314
box 0 0 1 1
use via1_x2_R90_128x8m81  via1_x2_R90_128x8m81_3
timestamp 1755005639
transform 0 -1 4502 1 0 18314
box 0 0 1 1
use via1_x2_R90_128x8m81  via1_x2_R90_128x8m81_4
timestamp 1755005639
transform 0 -1 925 1 0 8798
box 0 0 1 1
use via2_128x8m81  via2_128x8m81_0
timestamp 1755005639
transform 1 0 5448 0 1 18517
box 0 0 1 1
use via2_128x8m81  via2_128x8m81_1
timestamp 1755005639
transform 1 0 4394 0 1 18832
box 0 0 1 1
use via2_128x8m81  via2_128x8m81_2
timestamp 1755005639
transform 1 0 4210 0 1 19158
box 0 0 1 1
use via2_128x8m81  via2_128x8m81_3
timestamp 1755005639
transform 1 0 2971 0 1 20122
box 0 0 1 1
use via2_128x8m81  via2_128x8m81_4
timestamp 1755005639
transform 1 0 3156 0 1 19471
box 0 0 1 1
use via2_128x8m81  via2_128x8m81_5
timestamp 1755005639
transform 1 0 1917 0 1 20444
box 0 0 1 1
use via2_128x8m81  via2_128x8m81_6
timestamp 1755005639
transform 1 0 1733 0 1 20773
box 0 0 1 1
use via2_128x8m81  via2_128x8m81_7
timestamp 1755005639
transform 1 0 679 0 1 21092
box 0 0 1 1
use via2_x2_128x8m81  via2_x2_128x8m81_0
timestamp 1755005639
transform 1 0 2442 0 1 12351
box 0 0 1 1
use via2_x2_128x8m81  via2_x2_128x8m81_1
timestamp 1755005639
transform 1 0 2442 0 1 11575
box 0 0 1 1
use via2_x2_128x8m81  via2_x2_128x8m81_2
timestamp 1755005639
transform 1 0 2442 0 1 10659
box 0 0 1 1
use wen_wm1_128x8m81  wen_wm1_128x8m81_0
timestamp 1755005639
transform 1 0 322 0 1 -3369
box -156 -24 4946 3287
<< labels >>
rlabel metal3 s 810 18914 810 18914 4 ypass[1]
port 1 nsew
rlabel metal3 s 810 19231 810 19231 4 ypass[2]
port 2 nsew
rlabel metal3 s 810 19548 810 19548 4 ypass[3]
port 3 nsew
rlabel metal3 s 810 20204 810 20204 4 ypass[4]
port 4 nsew
rlabel metal3 s 810 20528 810 20528 4 ypass[5]
port 5 nsew
rlabel metal3 s 810 20845 810 20845 4 ypass[6]
port 6 nsew
rlabel metal3 s 810 21162 810 21162 4 ypass[7]
port 7 nsew
rlabel metal3 s 881 1467 881 1467 4 men
port 8 nsew
rlabel metal3 s 2918 1090 2918 1090 4 vss
port 9 nsew
rlabel metal3 s 2918 2179 2918 2179 4 vss
port 9 nsew
rlabel metal3 s 810 20204 810 20204 4 ypass[4]
port 4 nsew
rlabel metal3 s 3030 3831 3030 3831 4 vdd
port 10 nsew
rlabel metal3 s 2121 406 2121 406 4 vdd
port 10 nsew
rlabel metal3 s 2796 5470 2796 5470 4 vss
port 9 nsew
rlabel metal3 s 1878 11036 1878 11036 4 vss
port 9 nsew
rlabel metal3 s 810 21162 810 21162 4 ypass[7]
port 7 nsew
rlabel metal3 s 810 20845 810 20845 4 ypass[6]
port 6 nsew
rlabel metal3 s 810 20528 810 20528 4 ypass[5]
port 5 nsew
rlabel metal3 s 810 19548 810 19548 4 ypass[3]
port 3 nsew
rlabel metal3 s 810 19231 810 19231 4 ypass[2]
port 2 nsew
rlabel metal3 s 810 18914 810 18914 4 ypass[1]
port 1 nsew
rlabel metal3 s 810 18592 810 18592 4 ypass[0]
port 11 nsew
rlabel metal3 s 933 28902 933 28902 4 vdd
port 10 nsew
rlabel metal3 s 949 22015 949 22015 4 vss
port 9 nsew
rlabel metal3 s 933 18163 933 18163 4 vdd
port 10 nsew
rlabel metal3 s 973 16898 973 16898 4 vss
port 9 nsew
rlabel metal3 s 1807 13768 1807 13768 4 vdd
port 10 nsew
rlabel metal3 s 3303 7647 3303 7647 4 vdd
port 10 nsew
rlabel metal3 s 810 18592 810 18592 4 ypass[0]
port 11 nsew
flabel metal3 s 460 -586 460 -586 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 7098 460 7098 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 3309 460 3309 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 451 460 451 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 -2915 460 -2915 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 616 -1999 616 -1999 0 FreeSans 600 0 0 0 GWEN
port 13 nsew
flabel metal3 s 460 2469 460 2469 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 23368 460 23368 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 -2245 460 -2245 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 6326 460 6326 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 12529 460 12529 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 -1323 460 -1323 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 1081 460 1081 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 17115 460 17115 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 -1766 460 -1766 0 FreeSans 600 0 0 0 VSS
port 14 nsew
flabel metal3 s 460 8536 460 8536 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 13222 460 13222 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 460 18052 460 18052 0 FreeSans 600 0 0 0 VDD
port 12 nsew
flabel metal3 s 644 4966 644 4966 0 FreeSans 600 0 0 0 GWE
port 15 nsew
rlabel metal2 s 4862 28732 4862 28732 4 bb[1]
port 16 nsew
rlabel metal2 s 5073 28732 5073 28732 4 bb[0]
port 17 nsew
rlabel metal2 s 3832 28737 3832 28737 4 bb[2]
port 18 nsew
rlabel metal2 s 3632 28741 3632 28741 4 bb[3]
port 19 nsew
rlabel metal2 s 2593 28734 2593 28734 4 bb[4]
port 20 nsew
rlabel metal2 s 2387 28734 2387 28734 4 bb[5]
port 21 nsew
rlabel metal2 s 1155 28741 1155 28741 4 bb[7]
port 22 nsew
rlabel metal2 s 1355 28734 1355 28734 4 bb[6]
port 23 nsew
rlabel metal2 s 5499 28732 5499 28732 4 b[0]
port 24 nsew
rlabel metal2 s 4449 28732 4449 28732 4 b[1]
port 25 nsew
rlabel metal2 s 3006 28732 3006 28732 4 b[4]
port 26 nsew
rlabel metal2 s 1972 28732 1972 28732 4 b[5]
port 27 nsew
rlabel metal2 s 1770 28732 1770 28732 4 b[6]
port 28 nsew
rlabel metal2 s 736 28732 736 28732 4 b[7]
port 29 nsew
rlabel metal2 s 4251 28732 4251 28732 4 b[2]
port 30 nsew
rlabel metal2 s 3211 28732 3211 28732 4 b[3]
port 31 nsew
rlabel metal2 s 731 28732 731 28732 4 b[7]
port 29 nsew
rlabel metal2 s 488 1730 488 1730 4 datain
port 32 nsew
rlabel metal2 s 1768 28732 1768 28732 4 b[6]
port 28 nsew
rlabel metal2 s 1976 28732 1976 28732 4 b[5]
port 27 nsew
rlabel metal2 s 3004 28732 3004 28732 4 b[4]
port 26 nsew
rlabel metal2 s 3208 28732 3208 28732 4 b[3]
port 31 nsew
rlabel metal2 s 4249 28732 4249 28732 4 b[2]
port 30 nsew
rlabel metal2 s 4451 28732 4451 28732 4 b[1]
port 25 nsew
rlabel metal2 s 5497 28732 5497 28732 4 b[0]
port 24 nsew
rlabel metal2 s 1353 28734 1353 28734 4 bb[6]
port 23 nsew
rlabel metal2 s 1151 28741 1151 28741 4 bb[7]
port 22 nsew
rlabel metal2 s 2391 28734 2391 28734 4 bb[5]
port 21 nsew
rlabel metal2 s 1351 1131 1351 1131 4 q
port 33 nsew
rlabel metal2 s 2591 28734 2591 28734 4 bb[4]
port 20 nsew
rlabel metal2 s 3628 28741 3628 28741 4 bb[3]
port 19 nsew
rlabel metal2 s 3828 28737 3828 28737 4 bb[2]
port 18 nsew
rlabel metal2 s 5071 28732 5071 28732 4 bb[0]
port 17 nsew
rlabel metal2 s 4864 28732 4864 28732 4 bb[1]
port 16 nsew
rlabel metal2 s 1351 1131 1351 1131 4 q
port 33 nsew
rlabel metal1 s 993 27082 993 27082 4 pcb
port 34 nsew
rlabel metal1 s 698 8320 698 8320 4 datain
port 32 nsew
rlabel metal1 s 993 27079 993 27079 4 pcb
port 34 nsew
rlabel metal1 s 1801 15942 1801 15942 4 pcb
port 34 nsew
flabel metal1 s 722 -3358 722 -3358 0 FreeSans 600 0 0 0 WEN
port 35 nsew
<< properties >>
string FIXED_BBOX 2864 27052 2910 29928
string GDS_END 999192
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 989456
string path 14.435 135.260 14.435 149.640 
<< end >>
