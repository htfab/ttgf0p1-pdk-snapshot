magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 770 1486
<< nmos >>
rect 120 209 176 385
rect 280 209 336 385
rect 440 209 496 385
<< pmos >>
rect 120 1015 176 1191
rect 280 1015 336 1191
rect 440 1015 496 1191
<< ndiff >>
rect 32 268 120 385
rect 32 222 45 268
rect 91 222 120 268
rect 32 209 120 222
rect 176 209 280 385
rect 336 371 440 385
rect 336 325 365 371
rect 411 325 440 371
rect 336 209 440 325
rect 496 268 620 385
rect 496 222 561 268
rect 607 222 620 268
rect 496 209 620 222
<< pdiff >>
rect 32 1075 120 1191
rect 32 1029 45 1075
rect 91 1029 120 1075
rect 32 1015 120 1029
rect 176 1178 280 1191
rect 176 1132 205 1178
rect 251 1132 280 1178
rect 176 1015 280 1132
rect 336 1075 440 1191
rect 336 1029 365 1075
rect 411 1029 440 1075
rect 336 1015 440 1029
rect 496 1075 620 1191
rect 496 1029 561 1075
rect 607 1029 620 1075
rect 496 1015 620 1029
<< ndiffc >>
rect 45 222 91 268
rect 365 325 411 371
rect 561 222 607 268
<< pdiffc >>
rect 45 1029 91 1075
rect 205 1132 251 1178
rect 365 1029 411 1075
rect 561 1029 607 1075
<< psubdiff >>
rect 28 87 656 100
rect 28 41 69 87
rect 615 41 656 87
rect 28 28 656 41
<< nsubdiff >>
rect 28 1359 656 1372
rect 28 1313 69 1359
rect 615 1313 656 1359
rect 28 1300 656 1313
<< psubdiffcont >>
rect 69 41 615 87
<< nsubdiffcont >>
rect 69 1313 615 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 120 716 176 1015
rect 280 716 336 1015
rect 32 703 176 716
rect 32 657 45 703
rect 91 657 176 703
rect 32 644 176 657
rect 224 703 336 716
rect 224 657 237 703
rect 283 657 336 703
rect 224 644 336 657
rect 120 385 176 644
rect 280 385 336 644
rect 440 716 496 1015
rect 440 703 522 716
rect 440 657 463 703
rect 509 657 522 703
rect 440 644 522 657
rect 440 385 496 644
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
<< polycontact >>
rect 45 657 91 703
rect 237 657 283 703
rect 463 657 509 703
<< metal1 >>
rect 0 1359 684 1400
rect 0 1313 69 1359
rect 615 1313 684 1359
rect 0 1178 684 1313
rect 0 1132 205 1178
rect 251 1132 684 1178
rect 45 1075 411 1086
rect 91 1029 365 1075
rect 45 1018 411 1029
rect 42 703 94 972
rect 42 657 45 703
rect 91 657 94 703
rect 42 314 94 657
rect 234 703 286 972
rect 234 657 237 703
rect 283 657 286 703
rect 234 314 286 657
rect 460 703 512 1086
rect 460 657 463 703
rect 509 657 512 703
rect 460 428 512 657
rect 558 1075 610 1086
rect 558 1029 561 1075
rect 607 1029 610 1075
rect 558 382 610 1029
rect 365 371 610 382
rect 411 325 610 371
rect 365 314 610 325
rect 0 222 45 268
rect 91 222 561 268
rect 607 222 684 268
rect 0 87 684 222
rect 0 41 69 87
rect 615 41 684 87
rect 0 0 684 41
<< labels >>
rlabel metal1 s 0 0 684 268 4 vss
port 3 nsew
rlabel metal1 s 0 1132 684 1400 4 vdd
port 5 nsew
rlabel metal1 s 42 314 94 972 4 i0
port 7 nsew
rlabel metal1 s 558 314 610 1086 4 nq
port 9 nsew
rlabel metal1 s 234 314 286 972 4 i1
port 11 nsew
rlabel metal1 s 460 428 512 1086 4 i2
port 13 nsew
<< end >>
