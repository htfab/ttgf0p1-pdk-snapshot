magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
use pnp_10p00x00p42_0  pnp_10p00x00p42_0_0
timestamp 1755005639
transform 1 0 400 0 1 1360
box -338 -1296 338 1296
<< labels >>
flabel metal1 s 363 365 363 365 0 FreeSans 200 0 0 0 I1_default_E
port 1 nsew
flabel metal1 s 67 69 67 69 0 FreeSans 200 0 0 0 I1_default_C
port 2 nsew
flabel metal1 s 67 2577 67 2577 0 FreeSans 200 0 0 0 I1_default_C
port 2 nsew
flabel metal1 s 659 69 659 69 0 FreeSans 200 0 0 0 I1_default_C
port 2 nsew
flabel metal1 s 67 69 67 69 0 FreeSans 200 0 0 0 I1_default_C
port 2 nsew
flabel metal1 s 215 217 215 217 0 FreeSans 200 0 0 0 I1_default_B
port 3 nsew
flabel metal1 s 215 217 215 217 0 FreeSans 200 0 0 0 I1_default_B
port 3 nsew
flabel metal1 s 511 217 511 217 0 FreeSans 200 0 0 0 I1_default_B
port 3 nsew
flabel metal1 s 215 2429 215 2429 0 FreeSans 200 0 0 0 I1_default_B
port 3 nsew
<< properties >>
string GDS_END 11560
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_pr/gds/pnp_10p00x00p42.gds
string GDS_START 10866
<< end >>
