magic
tech gf180mcuD
magscale 1 10
timestamp 1751830969
<< nwell >>
rect -83 354 1545 870
<< pwell >>
rect -86 -86 1542 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 756 68 812 268
rect 916 68 972 268
rect 1076 68 1132 268
rect 1236 68 1292 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
rect 1076 440 1132 716
rect 1236 440 1292 716
<< ndiff >>
rect 28 249 116 268
rect 28 203 41 249
rect 87 203 116 249
rect 28 68 116 203
rect 172 127 276 268
rect 172 81 201 127
rect 247 81 276 127
rect 172 68 276 81
rect 332 249 436 268
rect 332 203 361 249
rect 407 203 436 249
rect 332 68 436 203
rect 492 127 596 268
rect 492 81 521 127
rect 567 81 596 127
rect 492 68 596 81
rect 652 249 756 268
rect 652 203 681 249
rect 727 203 756 249
rect 652 68 756 203
rect 812 249 916 268
rect 812 203 841 249
rect 887 203 916 249
rect 812 68 916 203
rect 972 152 1076 268
rect 972 106 1001 152
rect 1047 106 1076 152
rect 972 68 1076 106
rect 1132 249 1236 268
rect 1132 203 1161 249
rect 1207 203 1236 249
rect 1132 68 1236 203
rect 1292 152 1428 268
rect 1292 106 1321 152
rect 1367 106 1428 152
rect 1292 68 1428 106
<< pdiff >>
rect 28 703 116 716
rect 28 458 41 703
rect 87 458 116 703
rect 28 440 116 458
rect 172 542 276 716
rect 172 496 201 542
rect 247 496 276 542
rect 172 440 276 496
rect 332 703 436 716
rect 332 657 361 703
rect 407 657 436 703
rect 332 440 436 657
rect 492 542 596 716
rect 492 496 521 542
rect 567 496 596 542
rect 492 440 596 496
rect 652 703 756 716
rect 652 657 681 703
rect 727 657 756 703
rect 652 440 756 657
rect 812 542 916 716
rect 812 496 841 542
rect 887 496 916 542
rect 812 440 916 496
rect 972 703 1076 716
rect 972 657 1001 703
rect 1047 657 1076 703
rect 972 440 1076 657
rect 1132 667 1236 716
rect 1132 453 1161 667
rect 1207 453 1236 667
rect 1132 440 1236 453
rect 1292 703 1428 716
rect 1292 453 1321 703
rect 1367 453 1428 703
rect 1292 440 1428 453
<< ndiffc >>
rect 41 203 87 249
rect 201 81 247 127
rect 361 203 407 249
rect 521 81 567 127
rect 681 203 727 249
rect 841 203 887 249
rect 1001 106 1047 152
rect 1161 203 1207 249
rect 1321 106 1367 152
<< pdiffc >>
rect 41 458 87 703
rect 201 496 247 542
rect 361 657 407 703
rect 521 496 567 542
rect 681 657 727 703
rect 841 496 887 542
rect 1001 657 1047 703
rect 1161 453 1207 667
rect 1321 453 1367 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 1076 716 1132 760
rect 1236 716 1292 760
rect 116 411 172 440
rect 276 411 332 440
rect 436 411 492 440
rect 596 411 652 440
rect 116 386 652 411
rect 116 340 129 386
rect 629 340 652 386
rect 116 320 652 340
rect 116 268 172 320
rect 276 268 332 320
rect 436 268 492 320
rect 596 268 652 320
rect 756 410 812 440
rect 916 410 972 440
rect 1076 410 1132 440
rect 1236 410 1292 440
rect 756 391 1292 410
rect 756 345 779 391
rect 1108 345 1292 391
rect 756 319 1292 345
rect 756 268 812 319
rect 916 268 972 319
rect 1076 268 1132 319
rect 1236 268 1292 319
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
rect 1076 24 1132 68
rect 1236 24 1292 68
<< polycontact >>
rect 129 340 629 386
rect 779 345 1108 391
<< metal1 >>
rect 0 724 1456 844
rect 41 703 87 724
rect 361 703 407 724
rect 361 646 407 657
rect 681 703 727 724
rect 681 646 727 657
rect 1001 703 1047 724
rect 1321 703 1367 724
rect 1001 646 1047 657
rect 1161 667 1207 678
rect 164 496 201 542
rect 247 496 521 542
rect 567 496 841 542
rect 887 496 1161 542
rect 41 447 87 458
rect 116 386 629 411
rect 116 340 129 386
rect 116 320 629 340
rect 779 391 1108 410
rect 779 319 1108 345
rect 41 249 87 263
rect 361 249 407 263
rect 681 249 727 263
rect 1161 249 1233 453
rect 1321 427 1367 453
rect 87 203 361 249
rect 407 203 681 249
rect 817 203 841 249
rect 887 203 1161 249
rect 1207 203 1233 249
rect 41 190 87 203
rect 361 190 407 203
rect 681 152 727 203
rect 201 127 247 138
rect 201 60 247 81
rect 521 127 567 138
rect 681 106 1001 152
rect 1047 106 1321 152
rect 1367 106 1378 152
rect 521 60 567 81
rect 0 -60 1456 60
<< labels >>
flabel metal1 s 0 724 1456 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1456 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel nwell s 13 734 113 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel metal1 1161 203 1233 453 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 116 320 629 411 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 779 319 1108 410 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1456 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
