magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< obsm1 >>
rect -32 13108 52 69957
<< obsm2 >>
rect 0 49200 20 65000
<< metal3 >>
rect 0 68400 20 69678
rect 0 66800 20 68200
rect 0 65200 20 66600
rect 0 63600 20 65000
rect 0 62000 20 63400
rect 0 60400 20 61800
rect 0 58800 20 60200
rect 0 57200 20 58600
rect 0 55600 20 57000
rect 0 54000 20 55400
rect 0 52400 20 53800
rect 0 50800 20 52200
rect 0 49200 20 50600
rect 0 46000 20 49000
rect 0 42800 20 45800
rect 0 41200 20 42600
rect 0 39600 20 41000
rect 0 36400 20 39400
rect 0 33200 20 36200
rect 0 30000 20 33000
rect 0 26800 20 29800
rect 0 25200 20 26600
rect 0 23600 20 25000
rect 0 20400 20 23400
rect 0 17200 20 20200
rect 0 14000 20 17000
<< metal4 >>
rect 0 68400 20 69678
rect 0 66800 20 68200
rect 0 65200 20 66600
rect 0 63600 20 65000
rect 0 62000 20 63400
rect 0 60400 20 61800
rect 0 58800 20 60200
rect 0 57200 20 58600
rect 0 55600 20 57000
rect 0 54000 20 55400
rect 0 52400 20 53800
rect 0 50800 20 52200
rect 0 49200 20 50600
rect 0 46000 20 49000
rect 0 42800 20 45800
rect 0 41200 20 42600
rect 0 39600 20 41000
rect 0 36400 20 39400
rect 0 33200 20 36200
rect 0 30000 20 33000
rect 0 26800 20 29800
rect 0 25200 20 26600
rect 0 23600 20 25000
rect 0 20400 20 23400
rect 0 17200 20 20200
rect 0 14000 20 17000
<< metal5 >>
rect 0 68400 20 69678
rect 0 66800 20 68200
rect 0 65200 20 66600
rect 0 63600 20 65000
rect 0 62000 20 63400
rect 0 60400 20 61800
rect 0 58800 20 60200
rect 0 57200 20 58600
rect 0 55600 20 57000
rect 0 54000 20 55400
rect 0 52400 20 53800
rect 0 50800 20 52200
rect 0 49200 20 50600
rect 0 46000 20 49000
rect 0 42800 20 45800
rect 0 41200 20 42600
rect 0 39600 20 41000
rect 0 36400 20 39400
rect 0 33200 20 36200
rect 0 30000 20 33000
rect 0 26800 20 29800
rect 0 25200 20 26600
rect 0 23600 20 25000
rect 0 20400 20 23400
rect 0 17200 20 20200
rect 0 14000 20 17000
<< labels >>
rlabel metal3 s 0 66800 20 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 58800 20 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 55600 20 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 54000 20 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 52400 20 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 42800 20 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 41200 20 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 36400 20 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 33200 20 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 30000 20 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 26800 20 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 66800 20 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 58800 20 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 55600 20 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 54000 20 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 52400 20 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 42800 20 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 41200 20 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 36400 20 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 33200 20 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 30000 20 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 26800 20 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 66800 20 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 58800 20 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 55600 20 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 54000 20 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 52400 20 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 42800 20 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 41200 20 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 36400 20 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 33200 20 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 30000 20 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 26800 20 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 23600 20 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 23600 20 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 23600 20 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 68400 20 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 65200 20 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 60400 20 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 57200 20 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 46000 20 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 39600 20 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 25200 20 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 20400 20 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 17200 20 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 68400 20 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 65200 20 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 60400 20 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 57200 20 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 46000 20 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 39600 20 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 25200 20 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 20400 20 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 17200 20 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 68400 20 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 65200 20 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 60400 20 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 57200 20 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 46000 20 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 39600 20 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 25200 20 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 20400 20 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 17200 20 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 14000 20 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 14000 20 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 14000 20 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 62000 20 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 62000 20 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 0 62000 20 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 0 50800 20 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 50800 20 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 50800 20 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 63600 20 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 0 63600 20 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 63600 20 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 49200 20 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 0 49200 20 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 49200 20 50600 6 VSS
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20 70000
string LEFclass PAD SPACER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 17631666
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17626542
<< end >>
