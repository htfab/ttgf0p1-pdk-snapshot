magic
tech gf180mcuD
magscale 1 10
timestamp 1753952639
<< nwell >>
rect -86 354 2998 870
<< pwell >>
rect -86 -86 2998 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 756 68 812 268
rect 916 68 972 268
rect 1076 68 1132 268
rect 1236 68 1292 268
rect 1524 68 1580 268
rect 1684 68 1740 268
rect 1844 68 1900 268
rect 2004 68 2060 268
rect 2164 68 2220 268
rect 2324 68 2380 268
rect 2484 68 2540 268
rect 2644 68 2700 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
rect 1076 440 1132 716
rect 1236 440 1292 716
rect 1524 440 1580 716
rect 1684 440 1740 716
rect 1844 440 1900 716
rect 2004 440 2060 716
rect 2164 440 2220 716
rect 2324 440 2380 716
rect 2484 440 2540 716
rect 2644 440 2700 716
<< ndiff >>
rect 28 178 116 268
rect 28 132 41 178
rect 87 132 116 178
rect 28 68 116 132
rect 172 127 276 268
rect 172 81 201 127
rect 247 81 276 127
rect 172 68 276 81
rect 332 230 436 268
rect 332 184 361 230
rect 407 184 436 230
rect 332 68 436 184
rect 492 127 596 268
rect 492 81 521 127
rect 567 81 596 127
rect 492 68 596 81
rect 652 230 756 268
rect 652 184 681 230
rect 727 184 756 230
rect 652 68 756 184
rect 812 152 916 268
rect 812 106 841 152
rect 887 106 916 152
rect 812 68 916 106
rect 972 244 1076 268
rect 972 198 1001 244
rect 1047 198 1076 244
rect 972 68 1076 198
rect 1132 152 1236 268
rect 1132 106 1161 152
rect 1207 106 1236 152
rect 1132 68 1236 106
rect 1292 244 1380 268
rect 1292 198 1321 244
rect 1367 198 1380 244
rect 1292 68 1380 198
rect 1436 244 1524 268
rect 1436 198 1449 244
rect 1495 198 1524 244
rect 1436 68 1524 198
rect 1580 152 1684 268
rect 1580 106 1609 152
rect 1655 106 1684 152
rect 1580 68 1684 106
rect 1740 244 1844 268
rect 1740 198 1769 244
rect 1815 198 1844 244
rect 1740 68 1844 198
rect 1900 152 2004 268
rect 1900 106 1929 152
rect 1975 106 2004 152
rect 1900 68 2004 106
rect 2060 244 2164 268
rect 2060 198 2089 244
rect 2135 198 2164 244
rect 2060 68 2164 198
rect 2220 127 2324 268
rect 2220 81 2249 127
rect 2295 81 2324 127
rect 2220 68 2324 81
rect 2380 244 2484 268
rect 2380 198 2409 244
rect 2455 198 2484 244
rect 2380 68 2484 198
rect 2540 127 2644 268
rect 2540 81 2569 127
rect 2615 81 2644 127
rect 2540 68 2644 81
rect 2700 244 2788 268
rect 2700 198 2729 244
rect 2775 198 2788 244
rect 2700 68 2788 198
<< pdiff >>
rect 28 667 116 716
rect 28 453 41 667
rect 87 453 116 667
rect 28 440 116 453
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 667 436 716
rect 332 453 361 667
rect 407 453 436 667
rect 332 440 436 453
rect 492 703 596 716
rect 492 657 521 703
rect 567 657 596 703
rect 492 440 596 657
rect 652 667 756 716
rect 652 453 681 667
rect 727 453 756 667
rect 652 440 756 453
rect 812 703 916 716
rect 812 657 841 703
rect 887 657 916 703
rect 812 440 916 657
rect 972 667 1076 716
rect 972 453 1001 667
rect 1047 453 1076 667
rect 972 440 1076 453
rect 1132 703 1236 716
rect 1132 657 1161 703
rect 1207 657 1236 703
rect 1132 440 1236 657
rect 1292 667 1524 716
rect 1292 453 1321 667
rect 1367 453 1524 667
rect 1292 440 1524 453
rect 1580 703 1684 716
rect 1580 657 1609 703
rect 1655 657 1684 703
rect 1580 440 1684 657
rect 1740 667 1844 716
rect 1740 453 1769 667
rect 1815 453 1844 667
rect 1740 440 1844 453
rect 1900 703 2004 716
rect 1900 657 1929 703
rect 1975 657 2004 703
rect 1900 440 2004 657
rect 2060 678 2164 716
rect 2060 632 2089 678
rect 2135 632 2164 678
rect 2060 440 2164 632
rect 2220 586 2324 716
rect 2220 540 2249 586
rect 2295 540 2324 586
rect 2220 440 2324 540
rect 2380 678 2484 716
rect 2380 632 2409 678
rect 2455 632 2484 678
rect 2380 440 2484 632
rect 2540 586 2644 716
rect 2540 540 2569 586
rect 2615 540 2644 586
rect 2540 440 2644 540
rect 2700 678 2884 716
rect 2700 632 2729 678
rect 2775 632 2884 678
rect 2700 440 2884 632
<< ndiffc >>
rect 41 132 87 178
rect 201 81 247 127
rect 361 184 407 230
rect 521 81 567 127
rect 681 184 727 230
rect 841 106 887 152
rect 1001 198 1047 244
rect 1161 106 1207 152
rect 1321 198 1367 244
rect 1449 198 1495 244
rect 1609 106 1655 152
rect 1769 198 1815 244
rect 1929 106 1975 152
rect 2089 198 2135 244
rect 2249 81 2295 127
rect 2409 198 2455 244
rect 2569 81 2615 127
rect 2729 198 2775 244
<< pdiffc >>
rect 41 453 87 667
rect 201 657 247 703
rect 361 453 407 667
rect 521 657 567 703
rect 681 453 727 667
rect 841 657 887 703
rect 1001 453 1047 667
rect 1161 657 1207 703
rect 1321 453 1367 667
rect 1609 657 1655 703
rect 1769 453 1815 667
rect 1929 657 1975 703
rect 2089 632 2135 678
rect 2249 540 2295 586
rect 2409 632 2455 678
rect 2569 540 2615 586
rect 2729 632 2775 678
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 1076 716 1132 760
rect 1236 716 1292 760
rect 1524 716 1580 760
rect 1684 716 1740 760
rect 1844 716 1900 760
rect 2004 716 2060 760
rect 2164 716 2220 760
rect 2324 716 2380 760
rect 2484 716 2540 760
rect 2644 716 2700 760
rect 116 390 172 440
rect 276 390 332 440
rect 436 390 492 440
rect 596 390 652 440
rect 756 390 812 440
rect 916 390 972 440
rect 1076 390 1132 440
rect 1236 390 1292 440
rect 94 377 653 390
rect 94 331 107 377
rect 640 331 653 377
rect 94 318 653 331
rect 756 377 1292 390
rect 756 331 769 377
rect 1279 331 1292 377
rect 756 318 1292 331
rect 116 268 172 318
rect 276 268 332 318
rect 436 268 492 318
rect 596 268 652 318
rect 756 268 812 318
rect 916 268 972 318
rect 1076 268 1132 318
rect 1236 268 1292 318
rect 1524 390 1580 440
rect 1684 390 1740 440
rect 1844 390 1900 440
rect 2004 390 2060 440
rect 1524 377 2060 390
rect 1524 331 1537 377
rect 2047 331 2060 377
rect 1524 318 2060 331
rect 1524 268 1580 318
rect 1684 268 1740 318
rect 1844 268 1900 318
rect 2004 268 2060 318
rect 2164 390 2220 440
rect 2324 390 2380 440
rect 2484 390 2540 440
rect 2644 390 2700 440
rect 2164 377 2700 390
rect 2164 331 2177 377
rect 2687 331 2700 377
rect 2164 318 2700 331
rect 2164 268 2220 318
rect 2324 268 2380 318
rect 2484 268 2540 318
rect 2644 268 2700 318
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
rect 1076 24 1132 68
rect 1236 24 1292 68
rect 1524 24 1580 68
rect 1684 24 1740 68
rect 1844 24 1900 68
rect 2004 24 2060 68
rect 2164 24 2220 68
rect 2324 24 2380 68
rect 2484 24 2540 68
rect 2644 24 2700 68
<< polycontact >>
rect 107 331 640 377
rect 769 331 1279 377
rect 1537 331 2047 377
rect 2177 331 2687 377
<< metal1 >>
rect 0 724 2912 844
rect 201 703 247 724
rect 41 667 87 678
rect 521 703 567 724
rect 201 646 247 657
rect 361 667 407 678
rect 87 542 361 588
rect 41 440 87 453
rect 841 703 887 724
rect 521 646 567 657
rect 681 667 727 678
rect 407 542 681 588
rect 361 440 407 453
rect 1161 703 1207 724
rect 841 646 887 657
rect 1001 667 1047 678
rect 727 542 1001 588
rect 681 440 727 453
rect 1609 703 1655 724
rect 1161 646 1207 657
rect 1321 667 1367 678
rect 1047 542 1321 588
rect 1001 440 1047 453
rect 1929 703 1975 724
rect 1609 646 1655 657
rect 1769 667 1815 678
rect 1367 542 1769 588
rect 1321 440 1367 453
rect 1929 646 1975 657
rect 2070 632 2089 678
rect 2135 632 2409 678
rect 2455 632 2729 678
rect 2775 632 2786 678
rect 2070 588 2116 632
rect 1815 542 2116 588
rect 2237 540 2249 586
rect 2295 540 2569 586
rect 2615 540 2814 586
rect 1769 440 1815 453
rect 94 377 653 385
rect 94 331 107 377
rect 640 331 653 377
rect 94 323 653 331
rect 756 377 1292 390
rect 756 331 769 377
rect 1279 331 1292 377
rect 756 318 1292 331
rect 1524 377 2060 390
rect 1524 331 1537 377
rect 2047 331 2060 377
rect 1524 318 2060 331
rect 2164 377 2699 390
rect 2164 331 2177 377
rect 2687 331 2699 377
rect 2164 318 2699 331
rect 2745 244 2814 540
rect 680 230 1001 244
rect 41 184 361 230
rect 407 184 681 230
rect 727 198 1001 230
rect 1047 198 1321 244
rect 1367 198 1378 244
rect 1431 198 1449 244
rect 1495 198 1769 244
rect 1815 198 2089 244
rect 2135 198 2409 244
rect 2455 198 2729 244
rect 2775 198 2814 244
rect 727 184 740 198
rect 41 178 87 184
rect 41 106 87 132
rect 201 127 247 138
rect 201 60 247 81
rect 521 127 567 138
rect 814 106 841 152
rect 887 106 1161 152
rect 1207 106 1609 152
rect 1655 106 1929 152
rect 1975 106 1986 152
rect 2249 127 2295 138
rect 521 60 567 81
rect 2249 60 2295 81
rect 2569 127 2615 138
rect 2569 60 2615 81
rect 0 -60 2912 60
<< labels >>
flabel metal1 s 0 724 2912 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 2912 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 94 323 653 385 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel metal1 756 318 1292 390 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel metal1 1524 318 2060 390 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel metal1 2164 318 2699 390 0 FreeSans 200 0 0 0 D
port 8 nsew signal input
flabel metal1 2745 198 2814 586 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2912 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
