magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 4566 1094
<< pwell >>
rect -86 -86 4566 453
<< mvnmos >>
rect 145 150 265 308
rect 369 150 489 308
rect 763 215 883 333
rect 987 215 1107 333
rect 1211 215 1331 333
rect 1379 215 1499 333
rect 1637 215 1757 333
rect 1925 215 2045 333
rect 2093 215 2213 333
rect 2317 215 2437 333
rect 2541 215 2661 333
rect 3041 175 3161 333
rect 3225 175 3345 333
rect 3449 175 3569 333
rect 3617 175 3737 333
rect 3985 69 4105 333
rect 4209 69 4329 333
<< mvpmos >>
rect 165 573 265 849
rect 369 573 469 849
rect 717 589 817 789
rect 921 589 1021 789
rect 1125 589 1225 789
rect 1379 589 1479 789
rect 1657 688 1757 888
rect 2005 591 2105 791
rect 2285 591 2385 791
rect 2489 591 2589 791
rect 2693 591 2793 791
rect 3041 575 3141 851
rect 3245 575 3345 851
rect 3449 575 3549 851
rect 3653 575 3753 851
rect 4005 573 4105 939
rect 4209 573 4309 939
<< mvndiff >>
rect 57 295 145 308
rect 57 249 70 295
rect 116 249 145 295
rect 57 150 145 249
rect 265 209 369 308
rect 265 163 294 209
rect 340 163 369 209
rect 265 150 369 163
rect 489 295 577 308
rect 489 249 518 295
rect 564 249 577 295
rect 489 150 577 249
rect 675 274 763 333
rect 675 228 688 274
rect 734 228 763 274
rect 675 215 763 228
rect 883 320 987 333
rect 883 274 912 320
rect 958 274 987 320
rect 883 215 987 274
rect 1107 320 1211 333
rect 1107 274 1136 320
rect 1182 274 1211 320
rect 1107 215 1211 274
rect 1331 215 1379 333
rect 1499 215 1637 333
rect 1757 274 1925 333
rect 1757 228 1786 274
rect 1832 228 1925 274
rect 1757 215 1925 228
rect 2045 215 2093 333
rect 2213 320 2317 333
rect 2213 274 2242 320
rect 2288 274 2317 320
rect 2213 215 2317 274
rect 2437 320 2541 333
rect 2437 274 2466 320
rect 2512 274 2541 320
rect 2437 215 2541 274
rect 2661 285 2749 333
rect 2661 239 2690 285
rect 2736 239 2749 285
rect 2661 215 2749 239
rect 2949 234 3041 333
rect 2949 188 2962 234
rect 3008 188 3041 234
rect 2949 175 3041 188
rect 3161 175 3225 333
rect 3345 234 3449 333
rect 3345 188 3374 234
rect 3420 188 3449 234
rect 3345 175 3449 188
rect 3569 175 3617 333
rect 3737 320 3825 333
rect 3737 274 3766 320
rect 3812 274 3825 320
rect 3737 175 3825 274
rect 3897 222 3985 333
rect 3897 82 3910 222
rect 3956 82 3985 222
rect 3897 69 3985 82
rect 4105 320 4209 333
rect 4105 180 4134 320
rect 4180 180 4209 320
rect 4105 69 4209 180
rect 4329 222 4417 333
rect 4329 82 4358 222
rect 4404 82 4417 222
rect 4329 69 4417 82
<< mvpdiff >>
rect 1525 953 1597 966
rect 77 726 165 849
rect 77 586 90 726
rect 136 586 165 726
rect 77 573 165 586
rect 265 836 369 849
rect 265 696 294 836
rect 340 696 369 836
rect 265 573 369 696
rect 469 632 557 849
rect 1525 907 1538 953
rect 1584 907 1597 953
rect 2153 953 2225 966
rect 1525 888 1597 907
rect 2153 907 2166 953
rect 2212 907 2225 953
rect 2153 894 2225 907
rect 1525 872 1657 888
rect 1539 789 1657 872
rect 469 586 498 632
rect 544 586 557 632
rect 629 776 717 789
rect 629 730 642 776
rect 688 730 717 776
rect 629 589 717 730
rect 817 742 921 789
rect 817 602 846 742
rect 892 602 921 742
rect 817 589 921 602
rect 1021 742 1125 789
rect 1021 602 1050 742
rect 1096 602 1125 742
rect 1021 589 1125 602
rect 1225 747 1379 789
rect 1225 607 1304 747
rect 1350 607 1379 747
rect 1225 589 1379 607
rect 1479 688 1657 789
rect 1757 747 1845 888
rect 2165 791 2225 894
rect 3917 926 4005 939
rect 2953 838 3041 851
rect 2953 792 2966 838
rect 3012 792 3041 838
rect 1757 701 1786 747
rect 1832 701 1845 747
rect 1757 688 1845 701
rect 1917 747 2005 791
rect 1479 589 1559 688
rect 469 573 557 586
rect 1917 607 1930 747
rect 1976 607 2005 747
rect 1917 591 2005 607
rect 2105 591 2285 791
rect 2385 744 2489 791
rect 2385 604 2414 744
rect 2460 604 2489 744
rect 2385 591 2489 604
rect 2589 744 2693 791
rect 2589 604 2618 744
rect 2664 604 2693 744
rect 2589 591 2693 604
rect 2793 650 2881 791
rect 2793 604 2822 650
rect 2868 604 2881 650
rect 2793 591 2881 604
rect 2953 575 3041 792
rect 3141 634 3245 851
rect 3141 588 3170 634
rect 3216 588 3245 634
rect 3141 575 3245 588
rect 3345 838 3449 851
rect 3345 792 3374 838
rect 3420 792 3449 838
rect 3345 575 3449 792
rect 3549 639 3653 851
rect 3549 593 3578 639
rect 3624 593 3653 639
rect 3549 575 3653 593
rect 3753 838 3841 851
rect 3753 792 3782 838
rect 3828 792 3841 838
rect 3753 575 3841 792
rect 3917 786 3930 926
rect 3976 786 4005 926
rect 3917 573 4005 786
rect 4105 726 4209 939
rect 4105 586 4134 726
rect 4180 586 4209 726
rect 4105 573 4209 586
rect 4309 926 4397 939
rect 4309 786 4338 926
rect 4384 786 4397 926
rect 4309 573 4397 786
<< mvndiffc >>
rect 70 249 116 295
rect 294 163 340 209
rect 518 249 564 295
rect 688 228 734 274
rect 912 274 958 320
rect 1136 274 1182 320
rect 1786 228 1832 274
rect 2242 274 2288 320
rect 2466 274 2512 320
rect 2690 239 2736 285
rect 2962 188 3008 234
rect 3374 188 3420 234
rect 3766 274 3812 320
rect 3910 82 3956 222
rect 4134 180 4180 320
rect 4358 82 4404 222
<< mvpdiffc >>
rect 90 586 136 726
rect 294 696 340 836
rect 1538 907 1584 953
rect 2166 907 2212 953
rect 498 586 544 632
rect 642 730 688 776
rect 846 602 892 742
rect 1050 602 1096 742
rect 1304 607 1350 747
rect 2966 792 3012 838
rect 1786 701 1832 747
rect 1930 607 1976 747
rect 2414 604 2460 744
rect 2618 604 2664 744
rect 2822 604 2868 650
rect 3170 588 3216 634
rect 3374 792 3420 838
rect 3578 593 3624 639
rect 3782 792 3828 838
rect 3930 786 3976 926
rect 4134 586 4180 726
rect 4338 786 4384 926
<< polysilicon >>
rect 369 909 1021 949
rect 165 849 265 893
rect 369 849 469 909
rect 717 789 817 833
rect 921 789 1021 909
rect 1657 888 1757 932
rect 1125 868 1225 881
rect 1125 822 1138 868
rect 1184 822 1225 868
rect 1125 789 1225 822
rect 1379 789 1479 833
rect 2005 791 2105 835
rect 2285 931 3141 971
rect 4005 939 4105 983
rect 4209 939 4309 983
rect 2285 791 2385 931
rect 2489 870 2589 883
rect 2489 824 2502 870
rect 2548 824 2589 870
rect 3041 851 3141 931
rect 3245 851 3345 895
rect 3449 851 3549 895
rect 3653 851 3753 895
rect 2489 791 2589 824
rect 2693 791 2793 835
rect 165 411 265 573
rect 165 365 178 411
rect 224 365 265 411
rect 165 352 265 365
rect 145 308 265 352
rect 369 387 469 573
rect 717 545 817 589
rect 921 545 1021 589
rect 369 341 382 387
rect 428 352 469 387
rect 763 425 817 545
rect 1125 529 1225 589
rect 1067 489 1225 529
rect 763 412 883 425
rect 763 366 809 412
rect 855 366 883 412
rect 1067 377 1107 489
rect 1379 447 1479 589
rect 428 341 489 352
rect 369 308 489 341
rect 763 333 883 366
rect 987 333 1107 377
rect 1211 412 1331 425
rect 1211 366 1272 412
rect 1318 366 1331 412
rect 1211 333 1331 366
rect 1379 401 1420 447
rect 1466 401 1479 447
rect 1379 377 1479 401
rect 1657 377 1757 688
rect 2005 558 2105 591
rect 2005 512 2018 558
rect 2064 512 2105 558
rect 2285 531 2385 591
rect 2489 547 2589 591
rect 2005 499 2105 512
rect 2005 377 2045 499
rect 2173 491 2385 531
rect 2173 377 2213 491
rect 2541 377 2589 547
rect 2693 531 2793 591
rect 2693 491 2878 531
rect 1379 333 1499 377
rect 1637 333 1757 377
rect 1925 333 2045 377
rect 2093 333 2213 377
rect 2317 333 2437 377
rect 2541 333 2661 377
rect 763 171 883 215
rect 987 171 1107 215
rect 145 106 265 150
rect 369 90 489 150
rect 1211 90 1331 215
rect 1379 171 1499 215
rect 369 50 1331 90
rect 1637 75 1757 215
rect 1925 171 2045 215
rect 2093 171 2213 215
rect 2317 182 2437 215
rect 2317 136 2330 182
rect 2376 136 2437 182
rect 2541 171 2661 215
rect 2809 190 2878 491
rect 3041 412 3141 575
rect 3041 366 3065 412
rect 3111 377 3141 412
rect 3245 418 3345 575
rect 3245 377 3286 418
rect 3111 366 3161 377
rect 3041 333 3161 366
rect 3225 372 3286 377
rect 3332 372 3345 418
rect 3225 333 3345 372
rect 3449 510 3549 575
rect 3449 464 3490 510
rect 3536 464 3549 510
rect 3449 377 3549 464
rect 3653 542 3753 575
rect 3653 496 3692 542
rect 3738 496 3753 542
rect 3653 483 3753 496
rect 3653 377 3737 483
rect 4005 465 4105 573
rect 4209 529 4309 573
rect 4209 465 4308 529
rect 4005 412 4308 465
rect 4005 377 4018 412
rect 3449 333 3569 377
rect 3617 333 3737 377
rect 3985 366 4018 377
rect 4064 393 4308 412
rect 4064 366 4105 393
rect 3985 333 4105 366
rect 4209 377 4308 393
rect 4209 333 4329 377
rect 2806 182 2878 190
rect 2317 123 2437 136
rect 2806 136 2819 182
rect 2865 136 2878 182
rect 2806 123 2878 136
rect 3041 131 3161 175
rect 3225 131 3345 175
rect 3449 131 3569 175
rect 3617 131 3737 175
rect 3449 75 3489 131
rect 1637 35 3489 75
rect 3985 25 4105 69
rect 4209 25 4329 69
<< polycontact >>
rect 1138 822 1184 868
rect 2502 824 2548 870
rect 178 365 224 411
rect 382 341 428 387
rect 809 366 855 412
rect 1272 366 1318 412
rect 1420 401 1466 447
rect 2018 512 2064 558
rect 2330 136 2376 182
rect 3065 366 3111 412
rect 3286 372 3332 418
rect 3490 464 3536 510
rect 3692 496 3738 542
rect 4018 366 4064 412
rect 2819 136 2865 182
<< metal1 >>
rect 0 953 4480 1098
rect 0 918 1538 953
rect 294 836 340 918
rect 90 726 136 737
rect 642 776 688 918
rect 1584 918 2166 953
rect 1538 896 1584 907
rect 2212 926 4480 953
rect 2212 918 3930 926
rect 2166 896 2212 907
rect 642 719 688 730
rect 734 822 1138 868
rect 1184 850 1195 868
rect 2491 850 2502 870
rect 1184 824 2502 850
rect 2548 824 2559 870
rect 1184 822 2559 824
rect 734 804 2559 822
rect 2955 838 3023 918
rect 294 685 340 696
rect 734 643 780 804
rect 2955 792 2966 838
rect 3012 792 3023 838
rect 3363 838 3431 918
rect 3363 792 3374 838
rect 3420 792 3431 838
rect 3782 838 3828 918
rect 3782 781 3828 792
rect 3976 918 4338 926
rect 3930 775 3976 786
rect 4384 918 4480 926
rect 4338 775 4384 786
rect 498 632 780 643
rect 136 586 428 621
rect 90 575 428 586
rect 142 411 316 430
rect 142 365 178 411
rect 224 365 316 411
rect 142 354 316 365
rect 382 387 428 575
rect 382 308 428 341
rect 70 295 428 308
rect 116 262 428 295
rect 544 597 780 632
rect 846 742 892 753
rect 1050 742 1096 753
rect 892 602 958 637
rect 544 586 564 597
rect 846 591 958 602
rect 498 295 564 586
rect 678 412 866 430
rect 678 366 809 412
rect 855 366 866 412
rect 678 354 866 366
rect 70 238 116 249
rect 498 249 518 295
rect 498 238 564 249
rect 688 274 734 285
rect 798 242 866 354
rect 912 320 958 591
rect 1050 550 1096 602
rect 1304 747 1832 758
rect 1350 701 1786 747
rect 1350 690 1832 701
rect 1930 747 1976 758
rect 1304 596 1350 607
rect 2414 744 2460 755
rect 1976 615 2156 661
rect 1930 596 1976 607
rect 2018 558 2064 569
rect 1050 512 2018 550
rect 1050 504 2064 512
rect 912 263 958 274
rect 1136 320 1182 504
rect 2018 501 2064 504
rect 2110 491 2156 615
rect 2414 491 2460 604
rect 1420 455 2001 458
rect 2110 455 2460 491
rect 1420 447 2460 455
rect 1272 412 1318 423
rect 1466 445 2460 447
rect 2618 746 2927 755
rect 2618 744 3738 746
rect 2664 709 3738 744
rect 2899 700 3738 709
rect 1466 412 2288 445
rect 1984 409 2288 412
rect 1420 390 1466 401
rect 1272 344 1318 366
rect 1506 344 1967 366
rect 1272 320 1967 344
rect 1272 298 1546 320
rect 1136 263 1182 274
rect 283 163 294 209
rect 340 163 351 209
rect 283 90 351 163
rect 688 90 734 228
rect 1775 228 1786 274
rect 1832 228 1843 274
rect 1775 90 1843 228
rect 1921 182 1967 320
rect 2242 320 2288 409
rect 2618 380 2664 604
rect 2242 263 2288 274
rect 2466 334 2664 380
rect 2822 650 2868 661
rect 2466 320 2512 334
rect 2822 296 2868 604
rect 3170 634 3216 645
rect 2466 263 2512 274
rect 2690 285 2868 296
rect 2736 274 2868 285
rect 3054 366 3065 412
rect 3111 366 3122 412
rect 2736 239 3008 274
rect 3054 242 3122 366
rect 2690 234 3008 239
rect 2690 228 2962 234
rect 3170 196 3216 588
rect 3578 639 3646 650
rect 3624 593 3646 639
rect 3578 582 3646 593
rect 3351 510 3554 542
rect 3351 464 3490 510
rect 3536 464 3554 510
rect 3600 423 3646 582
rect 3692 542 3738 700
rect 3692 485 3738 496
rect 4134 726 4226 766
rect 4180 586 4226 726
rect 3600 418 4064 423
rect 3275 372 3286 418
rect 3332 412 4064 418
rect 3332 372 4018 412
rect 3766 366 4018 372
rect 3766 355 4064 366
rect 3766 320 3812 355
rect 3766 263 3812 274
rect 4134 320 4226 586
rect 3008 188 3216 196
rect 1921 136 2330 182
rect 2376 136 2819 182
rect 2865 136 2876 182
rect 2962 150 3216 188
rect 3374 234 3420 245
rect 3374 90 3420 188
rect 3910 222 3956 233
rect 0 82 3910 90
rect 4180 180 4226 320
rect 4134 169 4226 180
rect 4358 222 4404 233
rect 3956 82 4358 90
rect 4404 82 4480 90
rect 0 -90 4480 82
<< labels >>
flabel metal1 s 142 354 316 430 0 FreeSans 200 0 0 0 CLKN
port 4 nsew clock input
flabel metal1 s 678 354 866 430 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4134 169 4226 766 0 FreeSans 200 0 0 0 Q
port 5 nsew default output
flabel metal1 s 3351 464 3554 542 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 3054 242 3122 412 0 FreeSans 200 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 0 918 4480 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 688 274 734 285 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 798 242 866 354 1 D
port 1 nsew default input
rlabel metal1 s 4338 896 4384 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3930 896 3976 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3782 896 3828 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3363 896 3431 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2955 896 3023 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2166 896 2212 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1538 896 1584 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 642 896 688 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 896 340 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4338 792 4384 896 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3930 792 3976 896 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3782 792 3828 896 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3363 792 3431 896 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2955 792 3023 896 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 642 792 688 896 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 792 340 896 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4338 781 4384 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3930 781 3976 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3782 781 3828 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 642 781 688 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 781 340 792 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4338 775 4384 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3930 775 3976 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 642 775 688 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 775 340 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 642 719 688 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 719 340 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 685 340 719 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1775 245 1843 274 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 688 245 734 274 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3374 233 3420 245 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1775 233 1843 245 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 688 233 734 245 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4358 209 4404 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3910 209 3956 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3374 209 3420 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1775 209 1843 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 688 209 734 233 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4358 90 4404 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3910 90 3956 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3374 90 3420 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1775 90 1843 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 688 90 734 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 283 90 351 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4480 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4480 1008
string GDS_END 541412
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 531184
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
