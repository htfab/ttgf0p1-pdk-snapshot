* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__nor2b_2.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__nor2b_2 VDD VNW VPW VSS Y B A
X0 VSS a_220_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X1 a_220_68# A VSS VPW nfet_03v3 ad=0.44p pd=2.88u as=0.445p ps=2.89u w=1u l=0.28u
X2 Y a_220_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X3 a_220_68# A VDD VNW pfet_03v3 ad=0.6072p pd=3.64u as=0.6141p ps=3.65u w=1.38u l=0.28u
X4 VDD a_220_68# a_364_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X5 a_364_440# B Y VNW pfet_03v3 ad=0.7176p pd=3.8u as=0.3588p ps=1.9u w=1.38u l=0.28u
X6 VSS B Y VPW nfet_03v3 ad=0.515p pd=3.03u as=0.26p ps=1.52u w=1u l=0.28u
X7 a_364_440# a_220_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X8 Y B VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X9 Y B a_364_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
.ends

