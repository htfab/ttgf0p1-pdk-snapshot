magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -519 25300 21677 30562
rect -519 18840 21684 21394
<< metal1 >>
rect 14862 17525 15251 17663
rect 15677 17525 16256 17663
<< metal2 >>
rect -996 31419 -896 32609
rect -996 31363 -970 31419
rect -914 31363 -896 31419
rect -996 31287 -896 31363
rect -996 31231 -970 31287
rect -914 31231 -896 31287
rect -996 31155 -896 31231
rect -996 31099 -970 31155
rect -914 31099 -896 31155
rect -996 31023 -896 31099
rect -996 30967 -970 31023
rect -914 30967 -896 31023
rect -996 28954 -896 30967
rect -636 30505 -536 32609
rect -636 30449 -613 30505
rect -557 30449 -536 30505
rect -636 30373 -536 30449
rect -636 30317 -613 30373
rect -557 30317 -536 30373
rect -636 30241 -536 30317
rect -636 30185 -613 30241
rect -557 30185 -536 30241
rect -636 30109 -536 30185
rect -636 30053 -613 30109
rect -557 30053 -536 30109
rect -636 29977 -536 30053
rect -636 29921 -613 29977
rect -557 29921 -536 29977
rect -636 29845 -536 29921
rect -636 29789 -613 29845
rect -557 29789 -536 29845
rect -636 29713 -536 29789
rect -636 29657 -613 29713
rect -557 29657 -536 29713
rect -636 29581 -536 29657
rect -636 29525 -613 29581
rect -557 29525 -536 29581
rect -636 29449 -536 29525
rect -636 29393 -613 29449
rect -557 29393 -536 29449
rect -636 29317 -536 29393
rect -636 29261 -613 29317
rect -557 29261 -536 29317
rect -636 29185 -536 29261
rect -636 29129 -613 29185
rect -557 29129 -536 29185
rect -636 29053 -536 29129
rect -636 28997 -613 29053
rect -557 28997 -536 29053
rect -636 28949 -536 28997
rect 9804 31419 9904 32609
rect 9804 31363 9827 31419
rect 9883 31363 9904 31419
rect 9804 31287 9904 31363
rect 9804 31231 9827 31287
rect 9883 31231 9904 31287
rect 9804 31155 9904 31231
rect 9804 31099 9827 31155
rect 9883 31099 9904 31155
rect 9804 31023 9904 31099
rect 9804 30967 9827 31023
rect 9883 30967 9904 31023
rect 9804 28973 9904 30967
rect 10164 30505 10264 32609
rect 10164 30449 10190 30505
rect 10246 30449 10264 30505
rect 10164 30373 10264 30449
rect 10164 30317 10190 30373
rect 10246 30317 10264 30373
rect 10164 30241 10264 30317
rect 10164 30185 10190 30241
rect 10246 30185 10264 30241
rect 10164 30109 10264 30185
rect 10164 30053 10190 30109
rect 10246 30053 10264 30109
rect 10164 29977 10264 30053
rect 10164 29921 10190 29977
rect 10246 29921 10264 29977
rect 10164 29845 10264 29921
rect 10164 29789 10190 29845
rect 10246 29789 10264 29845
rect 10164 29713 10264 29789
rect 10164 29657 10190 29713
rect 10246 29657 10264 29713
rect 10164 29581 10264 29657
rect 10164 29525 10190 29581
rect 10246 29525 10264 29581
rect 10164 29449 10264 29525
rect 10164 29393 10190 29449
rect 10246 29393 10264 29449
rect 10164 29317 10264 29393
rect 10164 29261 10190 29317
rect 10246 29261 10264 29317
rect 10164 29185 10264 29261
rect 10164 29129 10190 29185
rect 10246 29129 10264 29185
rect 10164 29053 10264 29129
rect 10164 28997 10190 29053
rect 10246 28997 10264 29053
rect 10164 28972 10264 28997
rect 20604 30505 20704 32609
rect 20604 30449 20625 30505
rect 20681 30449 20704 30505
rect 20604 30373 20704 30449
rect 20604 30317 20625 30373
rect 20681 30317 20704 30373
rect 20604 30241 20704 30317
rect 20604 30185 20625 30241
rect 20681 30185 20704 30241
rect 20604 30109 20704 30185
rect 20604 30053 20625 30109
rect 20681 30053 20704 30109
rect 20604 29977 20704 30053
rect 20604 29921 20625 29977
rect 20681 29921 20704 29977
rect 20604 29845 20704 29921
rect 20604 29789 20625 29845
rect 20681 29789 20704 29845
rect 20604 29713 20704 29789
rect 20604 29657 20625 29713
rect 20681 29657 20704 29713
rect 20604 29581 20704 29657
rect 20604 29525 20625 29581
rect 20681 29525 20704 29581
rect 20604 29449 20704 29525
rect 20604 29393 20625 29449
rect 20681 29393 20704 29449
rect 20604 29317 20704 29393
rect 20604 29261 20625 29317
rect 20681 29261 20704 29317
rect 20604 29185 20704 29261
rect 20604 29129 20625 29185
rect 20681 29129 20704 29185
rect 20604 29053 20704 29129
rect 20604 28997 20625 29053
rect 20681 28997 20704 29053
rect 20604 28957 20704 28997
rect 20964 31419 21064 32609
rect 20964 31363 20988 31419
rect 21044 31363 21064 31419
rect 20964 31287 21064 31363
rect 20964 31231 20988 31287
rect 21044 31231 21064 31287
rect 20964 31155 21064 31231
rect 20964 31099 20988 31155
rect 21044 31099 21064 31155
rect 20964 31023 21064 31099
rect 20964 30967 20988 31023
rect 21044 30967 21064 31023
rect 20964 28960 21064 30967
<< via2 >>
rect -970 31363 -914 31419
rect -970 31231 -914 31287
rect -970 31099 -914 31155
rect -970 30967 -914 31023
rect -613 30449 -557 30505
rect -613 30317 -557 30373
rect -613 30185 -557 30241
rect -613 30053 -557 30109
rect -613 29921 -557 29977
rect -613 29789 -557 29845
rect -613 29657 -557 29713
rect -613 29525 -557 29581
rect -613 29393 -557 29449
rect -613 29261 -557 29317
rect -613 29129 -557 29185
rect -613 28997 -557 29053
rect 9827 31363 9883 31419
rect 9827 31231 9883 31287
rect 9827 31099 9883 31155
rect 9827 30967 9883 31023
rect 10190 30449 10246 30505
rect 10190 30317 10246 30373
rect 10190 30185 10246 30241
rect 10190 30053 10246 30109
rect 10190 29921 10246 29977
rect 10190 29789 10246 29845
rect 10190 29657 10246 29713
rect 10190 29525 10246 29581
rect 10190 29393 10246 29449
rect 10190 29261 10246 29317
rect 10190 29129 10246 29185
rect 10190 28997 10246 29053
rect 20625 30449 20681 30505
rect 20625 30317 20681 30373
rect 20625 30185 20681 30241
rect 20625 30053 20681 30109
rect 20625 29921 20681 29977
rect 20625 29789 20681 29845
rect 20625 29657 20681 29713
rect 20625 29525 20681 29581
rect 20625 29393 20681 29449
rect 20625 29261 20681 29317
rect 20625 29129 20681 29185
rect 20625 28997 20681 29053
rect 20988 31363 21044 31419
rect 20988 31231 21044 31287
rect 20988 31099 21044 31155
rect 20988 30967 21044 31023
<< metal3 >>
rect -1102 60770 21770 61130
rect -1102 59750 21770 60110
rect -1102 58970 21770 59330
rect -1102 57950 21770 58310
rect -1102 57170 21770 57530
rect -1102 56150 21770 56510
rect -1102 55370 21770 55730
rect -1102 54350 21770 54710
rect -1102 53570 21770 53930
rect -1102 52550 21770 52910
rect -1102 51770 21770 52130
rect -1102 50750 21770 51110
rect -1102 49970 21770 50330
rect -1102 48950 21770 49310
rect -1102 48170 21770 48530
rect -1102 47150 21770 47510
rect -1102 46370 21770 46730
rect -1102 45350 21770 45710
rect -1102 44570 21770 44930
rect -1102 43550 21770 43910
rect -1102 42770 21770 43130
rect -1102 41750 21770 42110
rect -1102 40970 21770 41330
rect -1102 39950 21770 40310
rect -1102 39170 21770 39530
rect -1102 38150 21770 38510
rect -1102 37370 21770 37730
rect -1102 36350 21770 36710
rect -1102 35570 21770 35930
rect -1102 34550 21770 34910
rect -1102 33770 21770 34130
rect -1102 32750 21770 33110
rect -1102 31970 21770 32330
rect -1173 31419 22177 31430
rect -1173 31363 -970 31419
rect -914 31363 9827 31419
rect 9883 31363 20988 31419
rect 21044 31363 22177 31419
rect -1173 31287 22177 31363
rect -1173 31231 -970 31287
rect -914 31231 9827 31287
rect 9883 31231 20988 31287
rect 21044 31231 22177 31287
rect -1173 31155 22177 31231
rect -1173 31099 -970 31155
rect -914 31099 9827 31155
rect 9883 31099 20988 31155
rect 21044 31099 22177 31155
rect -1173 31023 22177 31099
rect -1173 30967 -970 31023
rect -914 30967 9827 31023
rect 9883 30967 20988 31023
rect 21044 30967 22177 31023
rect -1173 30950 22177 30967
rect -1173 30505 22177 30539
rect -1173 30449 -613 30505
rect -557 30449 10190 30505
rect 10246 30449 20625 30505
rect 20681 30449 22177 30505
rect -1173 30373 22177 30449
rect -1173 30317 -613 30373
rect -557 30317 10190 30373
rect 10246 30317 20625 30373
rect 20681 30317 22177 30373
rect -1173 30241 22177 30317
rect -1173 30185 -613 30241
rect -557 30185 10190 30241
rect 10246 30185 20625 30241
rect 20681 30185 22177 30241
rect -1173 30109 22177 30185
rect -1173 30053 -613 30109
rect -557 30053 10190 30109
rect 10246 30053 20625 30109
rect 20681 30053 22177 30109
rect -1173 29977 22177 30053
rect -1173 29921 -613 29977
rect -557 29921 10190 29977
rect 10246 29921 20625 29977
rect 20681 29921 22177 29977
rect -1173 29845 22177 29921
rect -1173 29789 -613 29845
rect -557 29789 10190 29845
rect 10246 29789 20625 29845
rect 20681 29789 22177 29845
rect -1173 29713 22177 29789
rect -1173 29657 -613 29713
rect -557 29657 10190 29713
rect 10246 29657 20625 29713
rect 20681 29657 22177 29713
rect -1173 29581 22177 29657
rect -1173 29525 -613 29581
rect -557 29525 10190 29581
rect 10246 29525 20625 29581
rect 20681 29525 22177 29581
rect -1173 29449 22177 29525
rect -1173 29393 -613 29449
rect -557 29393 10190 29449
rect 10246 29393 20625 29449
rect 20681 29393 22177 29449
rect -1173 29317 22177 29393
rect -1173 29261 -613 29317
rect -557 29261 10190 29317
rect 10246 29261 20625 29317
rect 20681 29261 22177 29317
rect -1173 29185 22177 29261
rect -1173 29129 -613 29185
rect -557 29129 10190 29185
rect 10246 29129 20625 29185
rect 20681 29129 22177 29185
rect -1173 29053 22177 29129
rect -1173 28997 -613 29053
rect -557 28997 10190 29053
rect 10246 28997 20625 29053
rect 20681 28997 22177 29053
rect -1173 28730 22177 28997
rect -659 22523 21342 22738
rect -659 22201 21342 22416
rect -659 21880 21342 22095
rect -659 21558 21342 21773
rect -659 20866 21342 21081
rect -659 20544 21342 20759
rect -659 20223 21342 20438
rect -659 19901 21342 20116
rect -659 19352 21342 19794
rect -659 18241 21342 18696
rect -659 14430 21342 17153
rect -659 13011 20770 14144
rect -659 10742 21342 13011
rect -688 9875 21342 10592
rect 20913 9260 21342 9261
rect -688 8450 21342 9260
rect -659 6588 21342 7905
rect -659 6356 20885 6444
rect -659 4567 21342 5929
rect -659 3394 21342 4009
rect -659 2718 21342 3287
rect -659 2180 21342 2612
rect -659 1588 21342 2043
rect -696 474 21433 929
rect -696 -165 21433 186
rect -696 -377 21433 -289
rect -696 -608 21433 -520
rect -696 -1084 21433 -733
rect -696 -1809 21433 -1354
use Cell_array8x8x4_256x8m81  Cell_array8x8x4_256x8m81_0
timestamp 1755005639
transform 1 0 -1066 0 1 32540
box -68 -68 22268 28868
use M3_M24310590878117_256x8m81  M3_M24310590878117_256x8m81_0
timestamp 1755005639
transform 1 0 9855 0 1 31193
box 0 0 1 1
use M3_M24310590878117_256x8m81  M3_M24310590878117_256x8m81_1
timestamp 1755005639
transform 1 0 -942 0 1 31193
box 0 0 1 1
use M3_M24310590878117_256x8m81  M3_M24310590878117_256x8m81_2
timestamp 1755005639
transform 1 0 21016 0 1 31193
box 0 0 1 1
use M3_M24310590878118_256x8m81  M3_M24310590878118_256x8m81_0
timestamp 1755005639
transform 1 0 20653 0 1 29751
box 0 0 1 1
use M3_M24310590878118_256x8m81  M3_M24310590878118_256x8m81_1
timestamp 1755005639
transform 1 0 -585 0 1 29751
box 0 0 1 1
use M3_M24310590878118_256x8m81  M3_M24310590878118_256x8m81_2
timestamp 1755005639
transform 1 0 10218 0 1 29751
box 0 0 1 1
use saout_m2_256x8m81  saout_m2_256x8m81_0
timestamp 1755005639
transform 1 0 -953 0 1 1432
box -269 -3393 7633 31140
use saout_m2_256x8m81  saout_m2_256x8m81_1
timestamp 1755005639
transform 1 0 9847 0 1 1432
box -269 -3393 7633 31140
use saout_R_m2_256x8m81  saout_R_m2_256x8m81_0
timestamp 1755005639
transform -1 0 21021 0 1 1439
box -269 -3400 7633 31133
use saout_R_m2_256x8m81  saout_R_m2_256x8m81_1
timestamp 1755005639
transform -1 0 10221 0 1 1439
box -269 -3400 7633 31133
<< labels >>
rlabel metal1 s 16450 17361 16450 17361 4 pcb[0]
port 1 nsew
rlabel metal1 s 14237 17361 14237 17361 4 pcb[1]
port 2 nsew
rlabel metal1 s 3685 17361 3685 17361 4 pcb[3]
port 3 nsew
rlabel metal1 s 5628 17361 5628 17361 4 pcb[2]
port 4 nsew
flabel metal1 s -354 -1922 -354 -1922 0 FreeSans 600 0 0 0 WEN[3]
port 5 nsew
flabel metal1 s 9753 -1896 9753 -1896 0 FreeSans 600 0 0 0 WEN[2]
port 6 nsew
flabel metal1 s 10407 -1896 10407 -1896 0 FreeSans 600 0 0 0 WEN[1]
port 7 nsew
flabel metal1 s 20475 -1896 20475 -1896 0 FreeSans 600 0 0 0 WEN[0]
port 8 nsew
rlabel metal3 s -715 35703 -715 35703 4 WL[3]
port 9 nsew
rlabel metal3 s 810 20024 810 20024 4 ypass[0]
port 10 nsew
rlabel metal3 s 810 20346 810 20346 4 ypass[1]
port 11 nsew
rlabel metal3 s 810 20981 810 20981 4 ypass[3]
port 12 nsew
rlabel metal3 s 810 21636 810 21636 4 ypass[4]
port 13 nsew
rlabel metal3 s 810 21960 810 21960 4 ypass[5]
port 14 nsew
rlabel metal3 s 810 22595 810 22595 4 ypass[7]
port 15 nsew
rlabel metal3 s 881 2899 881 2899 4 men
port 16 nsew
flabel metal3 s -314 6410 -314 6410 0 FreeSans 448 0 0 0 GWE
port 17 nsew
flabel metal3 s -314 -1619 -314 -1619 0 FreeSans 448 0 0 0 VDD
port 18 nsew
flabel metal3 s -314 695 -314 695 0 FreeSans 448 0 0 0 VDD
port 18 nsew
rlabel metal3 s -715 34803 -715 34803 4 WL[2]
port 19 nsew
rlabel metal3 s -715 33903 -715 33903 4 WL[1]
port 20 nsew
rlabel metal3 s -715 60903 -715 60903 4 WL[31]
port 21 nsew
flabel metal3 s -314 1823 -314 1823 0 FreeSans 448 0 0 0 VDD
port 18 nsew
rlabel metal3 s -715 60003 -715 60003 4 WL[30]
port 22 nsew
rlabel metal3 s -715 59103 -715 59103 4 WL[29]
port 23 nsew
rlabel metal3 s -715 54603 -715 54603 4 WL[24]
port 24 nsew
rlabel metal3 s -715 53703 -715 53703 4 WL[23]
port 25 nsew
rlabel metal3 s -715 52803 -715 52803 4 WL[22]
port 26 nsew
rlabel metal3 s -715 51903 -715 51903 4 WL[21]
port 27 nsew
rlabel metal3 s -715 51003 -715 51003 4 WL[20]
port 28 nsew
rlabel metal3 s -715 50103 -715 50103 4 WL[19]
port 29 nsew
rlabel metal3 s -715 43803 -715 43803 4 WL[12]
port 30 nsew
rlabel metal3 s -715 42903 -715 42903 4 WL[11]
port 31 nsew
rlabel metal3 s -715 42003 -715 42003 4 WL[10]
port 32 nsew
rlabel metal3 s -715 41103 -715 41103 4 WL[9]
port 33 nsew
rlabel metal3 s -715 40203 -715 40203 4 WL[8]
port 34 nsew
rlabel metal3 s -715 39303 -715 39303 4 WL[7]
port 35 nsew
rlabel metal3 s -715 38403 -715 38403 4 WL[6]
port 36 nsew
rlabel metal3 s -715 37503 -715 37503 4 WL[5]
port 37 nsew
rlabel metal3 s -715 36603 -715 36603 4 WL[4]
port 38 nsew
rlabel metal3 s -715 49203 -715 49203 4 WL[18]
port 39 nsew
rlabel metal3 s -715 48303 -715 48303 4 WL[17]
port 40 nsew
rlabel metal3 s -715 47403 -715 47403 4 WL[16]
port 41 nsew
rlabel metal3 s -715 46503 -715 46503 4 WL[15]
port 42 nsew
rlabel metal3 s -715 45603 -715 45603 4 WL[14]
port 43 nsew
rlabel metal3 s -715 44703 -715 44703 4 WL[13]
port 44 nsew
rlabel metal3 s -715 58203 -715 58203 4 WL[28]
port 45 nsew
rlabel metal3 s -715 57303 -715 57303 4 WL[27]
port 46 nsew
rlabel metal3 s -715 56403 -715 56403 4 WL[26]
port 47 nsew
rlabel metal3 s -715 33003 -715 33003 4 WL[0]
port 48 nsew
rlabel metal3 s 811 22277 811 22277 4 ypass[6]
port 49 nsew
rlabel metal3 s 811 20663 811 20663 4 ypass[2]
port 50 nsew
rlabel metal3 s -715 55503 -715 55503 4 WL[25]
port 51 nsew
flabel metal3 s -314 2431 -314 2431 0 FreeSans 448 0 0 0 VSS
port 52 nsew
flabel metal3 s -314 3758 -314 3758 0 FreeSans 448 0 0 0 VSS
port 52 nsew
flabel metal3 s -314 5292 -314 5292 0 FreeSans 448 0 0 0 VDD
port 18 nsew
flabel metal3 s -314 9015 -314 9015 0 FreeSans 448 0 0 0 VDD
port 18 nsew
flabel metal3 s -314 15443 -314 15443 0 FreeSans 448 0 0 0 VDD
port 18 nsew
flabel metal3 s -314 19570 -314 19570 0 FreeSans 448 0 0 0 VDD
port 18 nsew
flabel metal3 s -314 29359 -314 29359 0 FreeSans 448 0 0 0 VDD
port 18 nsew
flabel metal3 s -314 31204 -314 31204 0 FreeSans 448 0 0 0 VSS
port 52 nsew
flabel metal3 s -314 24403 -314 24403 0 FreeSans 448 0 0 0 VSS
port 52 nsew
flabel metal3 s -314 18534 -314 18534 0 FreeSans 448 0 0 0 VSS
port 52 nsew
flabel metal3 s -314 12897 -314 12897 0 FreeSans 448 0 0 0 VSS
port 52 nsew
flabel metal3 s -314 7357 -314 7357 0 FreeSans 448 0 0 0 VSS
port 52 nsew
rlabel metal2 s 19247 30448 19247 30448 4 b[1]
port 53 nsew
rlabel metal2 s 17806 30448 17806 30448 4 b[4]
port 54 nsew
rlabel metal2 s 15531 30448 15531 30448 4 b[7]
port 55 nsew
rlabel metal2 s 14090 30448 14090 30448 4 b[10]
port 56 nsew
rlabel metal2 s 11815 30448 11815 30448 4 b[13]
port 57 nsew
rlabel metal2 s 9479 30448 9479 30448 4 b[16]
port 58 nsew
rlabel metal2 s 7203 30448 7203 30448 4 b[19]
port 59 nsew
rlabel metal2 s 5763 30448 5763 30448 4 b[22]
port 60 nsew
rlabel metal2 s 3488 30448 3488 30448 4 b[25]
port 61 nsew
rlabel metal2 s 2047 30448 2047 30448 4 b[28]
port 62 nsew
rlabel metal2 s -228 30448 -228 30448 4 b[31]
port 63 nsew
rlabel metal2 s 9710 1537 9710 1537 4 din[1]
port 64 nsew
rlabel metal2 s 20498 1537 20498 1537 4 din[3]
port 65 nsew
rlabel metal2 s 10349 1537 10349 1537 4 din[2]
port 66 nsew
rlabel metal2 s -447 1537 -447 1537 4 din[0]
port 67 nsew
rlabel metal2 s 402 1537 402 1537 4 q[0]
port 68 nsew
rlabel metal2 s 8866 1537 8866 1537 4 q[1]
port 69 nsew
rlabel metal2 s 11183 1537 11183 1537 4 q[2]
port 70 nsew
rlabel metal2 s 19659 1537 19659 1537 4 q[3]
port 71 nsew
rlabel metal2 s 1011 30448 1011 30448 4 b[29]
port 72 nsew
rlabel metal2 s 3286 30448 3286 30448 4 b[26]
port 73 nsew
rlabel metal2 s 4726 30448 4726 30448 4 b[23]
port 74 nsew
rlabel metal2 s 7001 30448 7001 30448 4 b[20]
port 75 nsew
rlabel metal2 s 8442 30448 8442 30448 4 b[17]
port 76 nsew
rlabel metal2 s 11613 30448 11613 30448 4 b[14]
port 77 nsew
rlabel metal2 s 13054 30448 13054 30448 4 b[11]
port 78 nsew
rlabel metal2 s 15329 30448 15329 30448 4 b[8]
port 79 nsew
rlabel metal2 s 16770 30448 16770 30448 4 b[5]
port 80 nsew
rlabel metal2 s 19045 30448 19045 30448 4 b[2]
port 81 nsew
rlabel metal2 s 19866 30448 19866 30448 4 bb[0]
port 82 nsew
rlabel metal2 s 19664 30448 19664 30448 4 bb[1]
port 83 nsew
rlabel metal2 s 18627 30448 18627 30448 4 bb[2]
port 84 nsew
rlabel metal2 s 18425 30448 18425 30448 4 bb[3]
port 85 nsew
rlabel metal2 s 17389 30448 17389 30448 4 bb[4]
port 86 nsew
rlabel metal2 s 17187 30448 17187 30448 4 bb[5]
port 87 nsew
rlabel metal2 s 16150 30448 16150 30448 4 bb[6]
port 88 nsew
rlabel metal2 s 15948 30448 15948 30448 4 bb[7]
port 89 nsew
rlabel metal2 s 14912 30448 14912 30448 4 bb[8]
port 90 nsew
rlabel metal2 s 14710 30448 14710 30448 4 bb[9]
port 91 nsew
rlabel metal2 s 13673 30448 13673 30448 4 bb[10]
port 92 nsew
rlabel metal2 s 13471 30448 13471 30448 4 bb[11]
port 93 nsew
rlabel metal2 s 12435 30448 12435 30448 4 bb[12]
port 94 nsew
rlabel metal2 s 12233 30448 12233 30448 4 bb[13]
port 95 nsew
rlabel metal2 s 11196 30448 11196 30448 4 bb[14]
port 96 nsew
rlabel metal2 s 10994 30448 10994 30448 4 bb[15]
port 97 nsew
rlabel metal2 s 9061 30448 9061 30448 4 bb[16]
port 98 nsew
rlabel metal2 s 8859 30448 8859 30448 4 bb[17]
port 99 nsew
rlabel metal2 s 7823 30448 7823 30448 4 bb[18]
port 100 nsew
rlabel metal2 s 7621 30448 7621 30448 4 bb[19]
port 101 nsew
rlabel metal2 s 6584 30448 6584 30448 4 bb[20]
port 102 nsew
rlabel metal2 s 6382 30448 6382 30448 4 bb[21]
port 103 nsew
rlabel metal2 s 5346 30448 5346 30448 4 bb[22]
port 104 nsew
rlabel metal2 s 5144 30448 5144 30448 4 bb[23]
port 105 nsew
rlabel metal2 s 4107 30448 4107 30448 4 bb[24]
port 106 nsew
rlabel metal2 s 3905 30448 3905 30448 4 bb[25]
port 107 nsew
rlabel metal2 s 2869 30448 2869 30448 4 bb[26]
port 108 nsew
rlabel metal2 s 2667 30448 2667 30448 4 bb[27]
port 109 nsew
rlabel metal2 s 1630 30448 1630 30448 4 bb[28]
port 110 nsew
rlabel metal2 s 1428 30448 1428 30448 4 bb[29]
port 111 nsew
rlabel metal2 s 391 30448 391 30448 4 bb[30]
port 112 nsew
rlabel metal2 s 189 30448 189 30448 4 bb[31]
port 113 nsew
rlabel metal2 s 809 30448 809 30448 4 b[30]
port 114 nsew
rlabel metal2 s 2249 30448 2249 30448 4 b[27]
port 115 nsew
rlabel metal2 s 4524 30448 4524 30448 4 b[24]
port 116 nsew
rlabel metal2 s 10577 30448 10577 30448 4 b[15]
port 117 nsew
rlabel metal2 s 12852 30448 12852 30448 4 b[12]
port 118 nsew
rlabel metal2 s 14292 30448 14292 30448 4 b[9]
port 119 nsew
rlabel metal2 s 5965 30448 5965 30448 4 b[21]
port 120 nsew
rlabel metal2 s 20283 30448 20283 30448 4 b[0]
port 121 nsew
rlabel metal2 s 18008 30448 18008 30448 4 b[3]
port 122 nsew
rlabel metal2 s 16568 30448 16568 30448 4 b[6]
port 123 nsew
rlabel metal2 s 8240 30448 8240 30448 4 b[18]
port 124 nsew
<< properties >>
string FIXED_BBOX 15379 30068 15489 32635
string GDS_END 1916604
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1903660
string path 50.175 142.140 50.175 307.040 
<< end >>
