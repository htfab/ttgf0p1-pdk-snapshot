* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__clkbuff_8.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__clkbuff_8 VDD VNW VPW VSS A Y
X0 VSS a_172_68# Y VPW nfet_03v3 ad=0.1872p pd=1.24u as=0.1872p ps=1.24u w=0.72u l=0.28u
X1 VDD A a_172_68# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X2 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X3 a_172_68# A VSS VPW nfet_03v3 ad=0.1872p pd=1.24u as=0.3168p ps=2.32u w=0.72u l=0.28u
X4 VSS a_172_68# Y VPW nfet_03v3 ad=0.1872p pd=1.24u as=0.1872p ps=1.24u w=0.72u l=0.28u
X5 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X6 Y a_172_68# VDD VNW pfet_03v3 ad=1.4904p pd=4.92u as=0.3588p ps=1.9u w=1.38u l=0.28u
X7 Y a_172_68# VSS VPW nfet_03v3 ad=0.1872p pd=1.24u as=0.1872p ps=1.24u w=0.72u l=0.28u
X8 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X9 Y a_172_68# VSS VPW nfet_03v3 ad=0.1872p pd=1.24u as=0.1872p ps=1.24u w=0.72u l=0.28u
X10 a_172_68# A VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X11 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X12 VSS a_172_68# a_172_68# VPW nfet_03v3 ad=0.1872p pd=1.24u as=0.1872p ps=1.24u w=0.72u l=0.28u
X13 VSS a_172_68# Y VPW nfet_03v3 ad=0.1872p pd=1.24u as=0.1872p ps=1.24u w=0.72u l=0.28u
X14 VDD a_172_68# a_172_68# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X15 a_172_68# A VSS VPW nfet_03v3 ad=0.1872p pd=1.24u as=0.1872p ps=1.24u w=0.72u l=0.28u
X16 Y a_172_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X17 VDD a_172_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X18 Y a_172_68# VSS VPW nfet_03v3 ad=0.1872p pd=1.24u as=0.1872p ps=1.24u w=0.72u l=0.28u
X19 a_172_68# A VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X20 VSS A a_172_68# VPW nfet_03v3 ad=0.1872p pd=1.24u as=0.1872p ps=1.24u w=0.72u l=0.28u
X21 Y a_172_68# VSS VPW nfet_03v3 ad=0.7776p pd=3.6u as=0.1872p ps=1.24u w=0.72u l=0.28u
.ends

