VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO nor3_x1
  CLASS BLOCK ;
  FOREIGN nor3_x1 ;
  ORIGIN 0.430 0.000 ;
  SIZE 4.280 BY 7.430 ;
  PIN vss
    ANTENNADIFFAREA 2.930400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 3.420 1.340 ;
    END
  END vss
  PIN vdd
    ANTENNADIFFAREA 2.043400 ;
    PORT
      LAYER Nwell ;
        RECT -0.430 3.400 3.850 7.430 ;
      LAYER Metal1 ;
        RECT 0.000 5.660 3.420 7.000 ;
    END
  END vdd
  PIN nq
    ANTENNADIFFAREA 2.713000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.610 2.910 2.870 5.430 ;
        RECT 1.025 1.570 2.870 2.910 ;
    END
  END nq
  PIN i0
    ANTENNAGATEAREA 1.106000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.210 1.570 0.470 5.430 ;
    END
  END i0
  PIN i1
    ANTENNAGATEAREA 1.106000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.170 3.140 1.430 5.430 ;
    END
  END i1
  PIN i2
    ANTENNAGATEAREA 1.106000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.970 3.140 2.230 5.430 ;
    END
  END i2
END nor3_x1
END LIBRARY

