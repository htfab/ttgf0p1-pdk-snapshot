magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 2366 1486
<< nmos >>
rect 120 209 176 385
rect 280 209 336 385
rect 600 209 656 385
rect 760 209 816 385
rect 920 209 976 385
rect 1080 209 1136 385
rect 1240 209 1296 385
rect 1400 209 1456 385
rect 1560 209 1616 385
rect 1720 209 1776 385
rect 1880 209 1936 385
rect 2084 209 2140 386
<< pmos >>
rect 120 1015 176 1191
rect 280 1015 336 1191
rect 600 1015 656 1191
rect 760 1015 816 1191
rect 920 1015 976 1191
rect 1080 1015 1136 1191
rect 1240 1015 1296 1191
rect 1400 1015 1456 1191
rect 1560 1015 1616 1191
rect 1720 1015 1776 1191
rect 1880 1015 1936 1191
rect 2084 974 2140 1191
<< ndiff >>
rect 1996 385 2084 386
rect 32 371 120 385
rect 32 325 45 371
rect 91 325 120 371
rect 32 209 120 325
rect 176 268 280 385
rect 176 222 205 268
rect 251 222 280 268
rect 176 209 280 222
rect 336 371 424 385
rect 336 325 365 371
rect 411 325 424 371
rect 336 209 424 325
rect 512 371 600 385
rect 512 325 525 371
rect 571 325 600 371
rect 512 209 600 325
rect 656 268 760 385
rect 656 222 685 268
rect 731 222 760 268
rect 656 209 760 222
rect 816 209 920 385
rect 976 371 1080 385
rect 976 325 1005 371
rect 1051 325 1080 371
rect 976 209 1080 325
rect 1136 209 1240 385
rect 1296 268 1400 385
rect 1296 222 1325 268
rect 1371 222 1400 268
rect 1296 209 1400 222
rect 1456 371 1560 385
rect 1456 325 1485 371
rect 1531 325 1560 371
rect 1456 209 1560 325
rect 1616 371 1720 385
rect 1616 325 1645 371
rect 1691 325 1720 371
rect 1616 209 1720 325
rect 1776 209 1880 385
rect 1936 268 2084 385
rect 1936 222 2009 268
rect 2055 222 2084 268
rect 1936 209 2084 222
rect 2140 372 2228 386
rect 2140 326 2169 372
rect 2215 326 2228 372
rect 2140 209 2228 326
<< pdiff >>
rect 32 1075 120 1191
rect 32 1029 45 1075
rect 91 1029 120 1075
rect 32 1015 120 1029
rect 176 1178 280 1191
rect 176 1132 205 1178
rect 251 1132 280 1178
rect 176 1015 280 1132
rect 336 1075 424 1191
rect 336 1029 365 1075
rect 411 1029 424 1075
rect 336 1015 424 1029
rect 512 1075 600 1191
rect 512 1029 525 1075
rect 571 1029 600 1075
rect 512 1015 600 1029
rect 656 1178 760 1191
rect 656 1132 685 1178
rect 731 1132 760 1178
rect 656 1015 760 1132
rect 816 1015 920 1191
rect 976 1075 1080 1191
rect 976 1029 1005 1075
rect 1051 1029 1080 1075
rect 976 1015 1080 1029
rect 1136 1015 1240 1191
rect 1296 1178 1400 1191
rect 1296 1132 1325 1178
rect 1371 1132 1400 1178
rect 1296 1015 1400 1132
rect 1456 1075 1560 1191
rect 1456 1029 1485 1075
rect 1531 1029 1560 1075
rect 1456 1015 1560 1029
rect 1616 1075 1720 1191
rect 1616 1029 1645 1075
rect 1691 1029 1720 1075
rect 1616 1015 1720 1029
rect 1776 1015 1880 1191
rect 1936 1178 2084 1191
rect 1936 1132 2009 1178
rect 2055 1132 2084 1178
rect 1936 1015 2084 1132
rect 1996 974 2084 1015
rect 2140 1054 2228 1191
rect 2140 1008 2169 1054
rect 2215 1008 2228 1054
rect 2140 974 2228 1008
<< ndiffc >>
rect 45 325 91 371
rect 205 222 251 268
rect 365 325 411 371
rect 525 325 571 371
rect 685 222 731 268
rect 1005 325 1051 371
rect 1325 222 1371 268
rect 1485 325 1531 371
rect 1645 325 1691 371
rect 2009 222 2055 268
rect 2169 326 2215 372
<< pdiffc >>
rect 45 1029 91 1075
rect 205 1132 251 1178
rect 365 1029 411 1075
rect 525 1029 571 1075
rect 685 1132 731 1178
rect 1005 1029 1051 1075
rect 1325 1132 1371 1178
rect 1485 1029 1531 1075
rect 1645 1029 1691 1075
rect 2009 1132 2055 1178
rect 2169 1008 2215 1054
<< psubdiff >>
rect 28 87 2252 100
rect 28 41 67 87
rect 2213 41 2252 87
rect 28 28 2252 41
<< nsubdiff >>
rect 28 1359 2252 1372
rect 28 1313 67 1359
rect 2213 1313 2252 1359
rect 28 1300 2252 1313
<< psubdiffcont >>
rect 67 41 2213 87
<< nsubdiffcont >>
rect 67 1313 2213 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 600 1191 656 1235
rect 760 1191 816 1235
rect 920 1191 976 1235
rect 1080 1191 1136 1235
rect 1240 1191 1296 1235
rect 1400 1191 1456 1235
rect 1560 1191 1616 1235
rect 1720 1191 1776 1235
rect 1880 1191 1936 1235
rect 2084 1191 2140 1235
rect 120 914 176 1015
rect 120 901 202 914
rect 120 855 143 901
rect 189 855 202 901
rect 120 842 202 855
rect 280 782 336 1015
rect 600 914 656 1015
rect 760 914 816 1015
rect 920 914 976 1015
rect 482 901 656 914
rect 482 855 495 901
rect 541 855 656 901
rect 482 842 656 855
rect 704 901 816 914
rect 704 855 717 901
rect 763 855 816 901
rect 704 842 816 855
rect 864 901 976 914
rect 864 855 877 901
rect 923 855 976 901
rect 864 842 976 855
rect 1080 782 1136 1015
rect 1240 914 1296 1015
rect 1400 914 1456 1015
rect 1184 901 1296 914
rect 1184 855 1197 901
rect 1243 855 1296 901
rect 1184 842 1296 855
rect 1344 901 1456 914
rect 1344 855 1357 901
rect 1403 855 1456 901
rect 1344 842 1456 855
rect 1560 782 1616 1015
rect 1720 914 1776 1015
rect 1664 901 1776 914
rect 1664 855 1677 901
rect 1723 855 1776 901
rect 1664 842 1776 855
rect 1880 782 1936 1015
rect 32 769 1740 782
rect 32 723 45 769
rect 91 723 877 769
rect 923 723 1681 769
rect 1727 723 1740 769
rect 32 710 1740 723
rect 1864 769 1936 782
rect 1864 723 1877 769
rect 1923 723 1936 769
rect 1864 710 1936 723
rect 120 637 202 650
rect 120 591 143 637
rect 189 591 202 637
rect 120 578 202 591
rect 120 385 176 578
rect 280 385 336 710
rect 2084 650 2140 974
rect 384 637 1642 650
rect 384 591 397 637
rect 443 591 975 637
rect 1021 591 1583 637
rect 1629 591 1642 637
rect 384 578 1642 591
rect 1766 637 2140 650
rect 1766 591 1779 637
rect 1825 591 2140 637
rect 1766 578 2140 591
rect 482 505 656 518
rect 482 459 495 505
rect 541 459 656 505
rect 482 446 656 459
rect 704 505 816 518
rect 704 459 717 505
rect 763 459 816 505
rect 704 446 816 459
rect 864 505 976 518
rect 864 459 877 505
rect 923 459 976 505
rect 864 446 976 459
rect 600 385 656 446
rect 760 385 816 446
rect 920 385 976 446
rect 1080 385 1136 578
rect 1184 505 1296 518
rect 1184 459 1197 505
rect 1243 459 1296 505
rect 1184 446 1296 459
rect 1344 505 1456 518
rect 1344 459 1357 505
rect 1403 459 1456 505
rect 1344 446 1456 459
rect 1240 385 1296 446
rect 1400 385 1456 446
rect 1560 385 1616 578
rect 1668 505 1776 518
rect 1668 459 1681 505
rect 1727 459 1776 505
rect 1668 446 1776 459
rect 1864 505 1936 518
rect 1864 459 1877 505
rect 1923 459 1936 505
rect 1864 446 1936 459
rect 1720 385 1776 446
rect 1880 385 1936 446
rect 2084 386 2140 578
rect 120 165 176 209
rect 280 165 336 209
rect 600 165 656 209
rect 760 165 816 209
rect 920 165 976 209
rect 1080 165 1136 209
rect 1240 165 1296 209
rect 1400 165 1456 209
rect 1560 165 1616 209
rect 1720 165 1776 209
rect 1880 165 1936 209
rect 2084 165 2140 209
<< polycontact >>
rect 143 855 189 901
rect 495 855 541 901
rect 717 855 763 901
rect 877 855 923 901
rect 1197 855 1243 901
rect 1357 855 1403 901
rect 1677 855 1723 901
rect 45 723 91 769
rect 877 723 923 769
rect 1681 723 1727 769
rect 1877 723 1923 769
rect 143 591 189 637
rect 397 591 443 637
rect 975 591 1021 637
rect 1583 591 1629 637
rect 1779 591 1825 637
rect 495 459 541 505
rect 717 459 763 505
rect 877 459 923 505
rect 1197 459 1243 505
rect 1357 459 1403 505
rect 1681 459 1727 505
rect 1877 459 1923 505
<< metal1 >>
rect 0 1359 2280 1400
rect 0 1313 67 1359
rect 2213 1313 2280 1359
rect 0 1178 2280 1313
rect 0 1132 205 1178
rect 251 1132 685 1178
rect 731 1132 1325 1178
rect 1371 1132 2009 1178
rect 2055 1132 2280 1178
rect 42 1075 94 1086
rect 42 1029 45 1075
rect 91 1029 94 1075
rect 42 769 94 1029
rect 42 723 45 769
rect 91 723 94 769
rect 42 371 94 723
rect 42 325 45 371
rect 91 325 94 371
rect 42 314 94 325
rect 140 901 192 1086
rect 140 855 143 901
rect 189 855 192 901
rect 140 637 192 855
rect 140 591 143 637
rect 189 591 192 637
rect 140 314 192 591
rect 362 1075 414 1086
rect 362 1029 365 1075
rect 411 1029 414 1075
rect 362 648 414 1029
rect 525 1075 766 1086
rect 571 1029 766 1075
rect 525 1018 766 1029
rect 1005 1075 1406 1086
rect 1051 1029 1406 1075
rect 1005 1018 1406 1029
rect 492 901 544 972
rect 492 855 495 901
rect 541 855 544 901
rect 362 637 443 648
rect 362 591 397 637
rect 362 580 443 591
rect 362 371 414 580
rect 492 505 544 855
rect 492 459 495 505
rect 541 459 544 505
rect 492 428 544 459
rect 714 901 766 1018
rect 714 855 717 901
rect 763 855 766 901
rect 714 505 766 855
rect 877 901 1024 912
rect 923 855 1024 901
rect 877 844 1024 855
rect 714 459 717 505
rect 763 459 766 505
rect 714 382 766 459
rect 874 769 926 780
rect 874 723 877 769
rect 923 723 926 769
rect 874 505 926 723
rect 972 637 1024 844
rect 972 591 975 637
rect 1021 591 1024 637
rect 972 580 1024 591
rect 874 459 877 505
rect 923 459 926 505
rect 874 448 926 459
rect 1070 382 1122 1018
rect 362 325 365 371
rect 411 325 414 371
rect 362 314 414 325
rect 525 371 766 382
rect 571 325 766 371
rect 525 314 766 325
rect 1005 371 1122 382
rect 1051 325 1122 371
rect 1005 314 1122 325
rect 1194 901 1246 912
rect 1194 855 1197 901
rect 1243 855 1246 901
rect 1194 505 1246 855
rect 1194 459 1197 505
rect 1243 459 1246 505
rect 1194 382 1246 459
rect 1354 901 1406 1018
rect 1354 855 1357 901
rect 1403 855 1406 901
rect 1354 505 1406 855
rect 1354 459 1357 505
rect 1403 459 1406 505
rect 1354 448 1406 459
rect 1482 1075 1534 1086
rect 1482 1029 1485 1075
rect 1531 1029 1534 1075
rect 1482 382 1534 1029
rect 1645 1075 1828 1086
rect 1691 1029 1828 1075
rect 1645 1018 1828 1029
rect 1580 901 1723 912
rect 1580 855 1677 901
rect 1580 844 1723 855
rect 1580 637 1632 844
rect 1580 591 1583 637
rect 1629 591 1632 637
rect 1580 580 1632 591
rect 1678 769 1730 780
rect 1678 723 1681 769
rect 1727 723 1730 769
rect 1678 505 1730 723
rect 1678 459 1681 505
rect 1727 459 1730 505
rect 1678 448 1730 459
rect 1776 637 1828 1018
rect 1776 591 1779 637
rect 1825 591 1828 637
rect 1776 382 1828 591
rect 1194 371 1534 382
rect 1194 325 1485 371
rect 1531 325 1534 371
rect 1194 314 1534 325
rect 1645 371 1828 382
rect 1691 325 1828 371
rect 1645 314 1828 325
rect 1874 1054 2215 1086
rect 1874 1008 2169 1054
rect 1874 997 2215 1008
rect 1874 769 1926 997
rect 1874 723 1877 769
rect 1923 723 1926 769
rect 1874 505 1926 723
rect 1874 459 1877 505
rect 1923 459 1926 505
rect 1874 383 1926 459
rect 1874 372 2215 383
rect 1874 326 2169 372
rect 1874 314 2215 326
rect 0 222 205 268
rect 251 222 685 268
rect 731 222 1325 268
rect 1371 222 2009 268
rect 2055 222 2280 268
rect 0 87 2280 222
rect 0 41 67 87
rect 2213 41 2280 87
rect 0 0 2280 41
<< labels >>
rlabel metal1 s 0 1132 2280 1400 4 vdd
port 3 nsew
rlabel metal1 s 0 0 2280 268 4 vss
port 5 nsew
rlabel metal1 s 140 314 192 1086 4 clk
port 7 nsew
rlabel metal1 s 492 428 544 972 4 i
port 9 nsew
rlabel metal1 s 1874 314 1926 1086 4 q
port 11 nsew
<< end >>
