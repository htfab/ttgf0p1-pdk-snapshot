module gf180mcu_ht_io__brk5_vss (VSS);
	inout	VSS;
endmodule

module gf180mcu_ht_io__brk5_vss_vdd (VSS, VDD);
	inout	VSS;
	inout	VDD;
endmodule

module gf180mcu_ht_io__brk5_vss_dvss (VSS, DVSS);
	inout	VSS;
	inout	DVSS;
endmodule

module gf180mcu_ht_io__brk5_vss_vdd_dvss (VSS, VDD, DVSS);
	inout	VSS;
	inout	VDD;
	inout	DVSS;
endmodule

module gf180mcu_ht_io__brk5_vss_dvdd (VSS, DVDD);
	inout	VSS;
	inout	DVDD;
endmodule

module gf180mcu_ht_io__brk5_vss_vdd_dvdd (VSS, VDD, DVDD);
	inout	VSS;
	inout	VDD;
	inout	DVDD;
endmodule

module gf180mcu_ht_io__brk5_vss_dvss_dvdd (VSS, DVSS, DVDD);
	inout	VSS;
	inout	DVSS;
	inout	DVDD;
endmodule

module gf180mcu_ht_io__brk5_vss_vdd_dvss_dvdd (VSS, VDD, DVSS, DVDD);
	inout	VSS;
	inout	VDD;
	inout	DVSS;
	inout	DVDD;
endmodule

