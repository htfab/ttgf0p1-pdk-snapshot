VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO or2_x1
  CLASS BLOCK ;
  FOREIGN or2_x1 ;
  ORIGIN 0.430 0.000 ;
  SIZE 4.280 BY 7.430 ;
  PIN vss
    ANTENNADIFFAREA 2.606600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 3.420 1.340 ;
    END
  END vss
  PIN vdd
    ANTENNADIFFAREA 2.307400 ;
    PORT
      LAYER Nwell ;
        RECT -0.430 3.400 3.850 7.430 ;
      LAYER Metal1 ;
        RECT 0.000 5.660 3.420 7.000 ;
    END
  END vdd
  PIN i0
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.210 1.570 0.470 4.860 ;
    END
  END i0
  PIN i1
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.170 2.140 1.430 4.860 ;
    END
  END i1
  PIN q
    ANTENNADIFFAREA 1.738000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.830 1.570 3.090 5.430 ;
    END
  END q
  OBS
      LAYER Metal1 ;
        RECT 0.225 5.090 2.230 5.430 ;
        RECT 1.970 1.910 2.230 5.090 ;
        RECT 1.025 1.570 2.230 1.910 ;
  END
END or2_x1
END LIBRARY

