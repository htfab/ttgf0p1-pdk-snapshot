magic
tech gf180mcuD
timestamp 1755005639
<< properties >>
string GDS_END 5346506
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 5342534
<< end >>
