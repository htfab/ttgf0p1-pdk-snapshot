magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 377 5126 870
rect -86 352 645 377
rect 2851 352 5126 377
<< pwell >>
rect 645 352 2851 377
rect -86 -86 5126 352
<< metal1 >>
rect 0 724 5040 844
rect 241 586 311 724
rect 602 601 670 724
rect 1506 689 1574 724
rect 2146 689 2214 724
rect 141 120 214 430
rect 273 60 319 232
rect 570 330 792 430
rect 702 60 770 230
rect 1770 60 1838 183
rect 3025 586 3093 724
rect 3454 586 3522 724
rect 2913 334 3191 445
rect 3343 357 3623 426
rect 3873 546 3919 724
rect 4017 506 4063 724
rect 4209 472 4267 676
rect 4414 524 4482 724
rect 4612 472 4684 676
rect 4833 506 4879 724
rect 4209 456 4684 472
rect 4209 425 4801 456
rect 3434 60 3502 215
rect 4628 263 4801 425
rect 4209 217 4801 263
rect 3985 60 4031 181
rect 4209 131 4255 217
rect 4433 60 4479 153
rect 4628 120 4801 217
rect 4881 60 4927 181
rect 0 -60 5040 60
<< obsm1 >>
rect 49 540 95 645
rect 457 545 503 645
rect 730 632 999 678
rect 1156 643 1460 678
rect 1636 643 2096 678
rect 2260 643 2550 659
rect 1156 632 2550 643
rect 730 545 776 632
rect 49 476 407 540
rect 49 162 95 476
rect 361 256 407 476
rect 457 498 776 545
rect 457 221 503 498
rect 861 241 907 586
rect 953 379 999 632
rect 1414 597 1682 632
rect 2049 613 2550 632
rect 2609 624 2963 671
rect 2049 597 2306 613
rect 1065 459 1111 588
rect 1258 551 1326 577
rect 1754 551 1822 586
rect 1258 505 1822 551
rect 1898 551 1966 586
rect 2394 551 2462 567
rect 1898 505 2462 551
rect 1065 413 2072 459
rect 1065 408 1207 413
rect 457 153 543 221
rect 861 173 983 241
rect 1161 173 1207 408
rect 2256 367 2302 505
rect 2609 459 2655 624
rect 1253 275 1299 337
rect 1406 321 2302 367
rect 2480 412 2655 459
rect 1253 229 2176 275
rect 2130 152 2176 229
rect 2234 198 2302 321
rect 2349 152 2400 347
rect 2480 244 2526 412
rect 2701 366 2747 486
rect 2458 198 2526 244
rect 2579 320 2747 366
rect 2579 152 2625 320
rect 2813 244 2859 578
rect 2917 540 2963 624
rect 3139 618 3407 665
rect 3139 540 3185 618
rect 2917 493 3185 540
rect 3237 493 3307 561
rect 3361 540 3407 618
rect 3577 607 3807 654
rect 3577 540 3623 607
rect 3361 493 3623 540
rect 2682 215 2859 244
rect 3237 215 3283 493
rect 3669 311 3715 561
rect 3761 401 3807 607
rect 4061 311 4578 357
rect 3329 265 4119 311
rect 2682 198 3283 215
rect 2813 169 3283 198
rect 2130 106 2625 152
rect 3841 158 3887 265
<< labels >>
rlabel metal1 s 570 330 792 430 6 D
port 1 nsew default input
rlabel metal1 s 3343 357 3623 426 6 RN
port 2 nsew default input
rlabel metal1 s 2913 334 3191 445 6 SETN
port 3 nsew default input
rlabel metal1 s 141 120 214 430 6 CLK
port 4 nsew clock input
rlabel metal1 s 4628 120 4801 217 6 Q
port 5 nsew default output
rlabel metal1 s 4209 131 4255 217 6 Q
port 5 nsew default output
rlabel metal1 s 4209 217 4801 263 6 Q
port 5 nsew default output
rlabel metal1 s 4628 263 4801 425 6 Q
port 5 nsew default output
rlabel metal1 s 4209 425 4801 456 6 Q
port 5 nsew default output
rlabel metal1 s 4209 456 4684 472 6 Q
port 5 nsew default output
rlabel metal1 s 4612 472 4684 676 6 Q
port 5 nsew default output
rlabel metal1 s 4209 472 4267 676 6 Q
port 5 nsew default output
rlabel metal1 s 4833 506 4879 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4414 524 4482 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4017 506 4063 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3873 546 3919 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3454 586 3522 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3025 586 3093 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2146 689 2214 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1506 689 1574 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 602 601 670 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 241 586 311 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 724 5040 844 6 VDD
port 6 nsew power bidirectional abutment
rlabel nwell s 2851 352 5126 377 6 VNW
port 7 nsew power bidirectional
rlabel nwell s -86 352 645 377 6 VNW
port 7 nsew power bidirectional
rlabel nwell s -86 377 5126 870 6 VNW
port 7 nsew power bidirectional
rlabel pwell s -86 -86 5126 352 6 VPW
port 8 nsew ground bidirectional
rlabel pwell s 645 352 2851 377 6 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 0 -60 5040 60 8 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4881 60 4927 181 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4433 60 4479 153 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3985 60 4031 181 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3434 60 3502 215 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1770 60 1838 183 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 702 60 770 230 6 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 232 6 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5040 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1049066
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1038088
<< end >>
