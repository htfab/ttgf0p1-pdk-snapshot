magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
use pnp_10p00x10p00_0  pnp_10p00x10p00_0_0
timestamp 1755005639
transform 1 0 1360 0 1 1360
box -1296 -1296 1296 1296
<< labels >>
flabel metal1 s 365 365 365 365 0 FreeSans 200 0 0 0 I1_default_E
port 3 nsew
flabel metal1 s 69 69 69 69 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 69 69 69 69 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 2577 69 2577 69 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 69 2577 69 2577 0 FreeSans 200 0 0 0 I1_default_C
port 1 nsew
flabel metal1 s 217 217 217 217 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
flabel metal1 s 217 217 217 217 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
flabel metal1 s 2429 217 2429 217 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
flabel metal1 s 217 2429 217 2429 0 FreeSans 200 0 0 0 I1_default_B
port 2 nsew
<< properties >>
string GDS_END 41064
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_pr/gds/pnp_10p00x10p00.gds
string GDS_START 40370
string device primitive
<< end >>
