magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 3782 1094
<< pwell >>
rect -86 -86 3782 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 978 68 1098 332
rect 1202 68 1322 332
rect 1426 68 1546 332
rect 1650 68 1770 332
rect 1874 68 1994 332
rect 2098 68 2218 332
rect 2322 68 2442 332
rect 2546 68 2666 332
rect 2770 68 2890 332
rect 2994 68 3114 332
rect 3218 68 3338 332
rect 3442 68 3562 332
<< mvpmos >>
rect 124 573 224 933
rect 328 573 428 933
rect 660 573 760 933
rect 1058 580 1158 940
rect 1262 580 1362 940
rect 1466 580 1566 940
rect 1670 580 1770 940
rect 1874 580 1974 940
rect 2078 580 2178 940
rect 2282 580 2382 940
rect 2486 580 2586 940
rect 2690 580 2790 940
rect 2894 580 2994 940
rect 3098 580 3198 940
rect 3302 580 3402 940
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 69 124 274
rect 244 128 348 333
rect 244 82 273 128
rect 319 82 348 128
rect 244 69 348 82
rect 468 287 572 333
rect 468 147 497 287
rect 543 147 572 287
rect 468 69 572 147
rect 692 320 780 333
rect 692 274 721 320
rect 767 274 780 320
rect 692 69 780 274
rect 852 125 978 332
rect 852 79 865 125
rect 911 79 978 125
rect 852 68 978 79
rect 1098 228 1202 332
rect 1098 182 1127 228
rect 1173 182 1202 228
rect 1098 68 1202 182
rect 1322 127 1426 332
rect 1322 81 1351 127
rect 1397 81 1426 127
rect 1322 68 1426 81
rect 1546 287 1650 332
rect 1546 147 1575 287
rect 1621 147 1650 287
rect 1546 68 1650 147
rect 1770 127 1874 332
rect 1770 81 1799 127
rect 1845 81 1874 127
rect 1770 68 1874 81
rect 1994 273 2098 332
rect 1994 227 2023 273
rect 2069 227 2098 273
rect 1994 68 2098 227
rect 2218 127 2322 332
rect 2218 81 2247 127
rect 2293 81 2322 127
rect 2218 68 2322 81
rect 2442 319 2546 332
rect 2442 179 2471 319
rect 2517 179 2546 319
rect 2442 68 2546 179
rect 2666 127 2770 332
rect 2666 81 2695 127
rect 2741 81 2770 127
rect 2666 68 2770 81
rect 2890 319 2994 332
rect 2890 179 2919 319
rect 2965 179 2994 319
rect 2890 68 2994 179
rect 3114 127 3218 332
rect 3114 81 3143 127
rect 3189 81 3218 127
rect 3114 68 3218 81
rect 3338 319 3442 332
rect 3338 179 3367 319
rect 3413 179 3442 319
rect 3338 68 3442 179
rect 3562 221 3650 332
rect 3562 81 3591 221
rect 3637 81 3650 221
rect 3562 68 3650 81
rect 852 66 918 68
<< mvpdiff >>
rect 36 726 124 933
rect 36 586 49 726
rect 95 586 124 726
rect 36 573 124 586
rect 224 920 328 933
rect 224 780 253 920
rect 299 780 328 920
rect 224 573 328 780
rect 428 818 660 933
rect 428 678 585 818
rect 631 678 660 818
rect 428 573 660 678
rect 760 726 848 933
rect 760 586 789 726
rect 835 586 848 726
rect 760 573 848 586
rect 970 927 1058 940
rect 970 787 983 927
rect 1029 787 1058 927
rect 970 580 1058 787
rect 1158 639 1262 940
rect 1158 593 1187 639
rect 1233 593 1262 639
rect 1158 580 1262 593
rect 1362 927 1466 940
rect 1362 787 1391 927
rect 1437 787 1466 927
rect 1362 580 1466 787
rect 1566 755 1670 940
rect 1566 615 1595 755
rect 1641 615 1670 755
rect 1566 580 1670 615
rect 1770 927 1874 940
rect 1770 787 1799 927
rect 1845 787 1874 927
rect 1770 580 1874 787
rect 1974 709 2078 940
rect 1974 663 2003 709
rect 2049 663 2078 709
rect 1974 580 2078 663
rect 2178 927 2282 940
rect 2178 881 2207 927
rect 2253 881 2282 927
rect 2178 580 2282 881
rect 2382 756 2486 940
rect 2382 616 2411 756
rect 2457 616 2486 756
rect 2382 580 2486 616
rect 2586 927 2690 940
rect 2586 881 2615 927
rect 2661 881 2690 927
rect 2586 580 2690 881
rect 2790 756 2894 940
rect 2790 616 2819 756
rect 2865 616 2894 756
rect 2790 580 2894 616
rect 2994 927 3098 940
rect 2994 881 3023 927
rect 3069 881 3098 927
rect 2994 580 3098 881
rect 3198 756 3302 940
rect 3198 616 3227 756
rect 3273 616 3302 756
rect 3198 580 3302 616
rect 3402 927 3490 940
rect 3402 787 3431 927
rect 3477 787 3490 927
rect 3402 580 3490 787
<< mvndiffc >>
rect 49 274 95 320
rect 273 82 319 128
rect 497 147 543 287
rect 721 274 767 320
rect 865 79 911 125
rect 1127 182 1173 228
rect 1351 81 1397 127
rect 1575 147 1621 287
rect 1799 81 1845 127
rect 2023 227 2069 273
rect 2247 81 2293 127
rect 2471 179 2517 319
rect 2695 81 2741 127
rect 2919 179 2965 319
rect 3143 81 3189 127
rect 3367 179 3413 319
rect 3591 81 3637 221
<< mvpdiffc >>
rect 49 586 95 726
rect 253 780 299 920
rect 585 678 631 818
rect 789 586 835 726
rect 983 787 1029 927
rect 1187 593 1233 639
rect 1391 787 1437 927
rect 1595 615 1641 755
rect 1799 787 1845 927
rect 2003 663 2049 709
rect 2207 881 2253 927
rect 2411 616 2457 756
rect 2615 881 2661 927
rect 2819 616 2865 756
rect 3023 881 3069 927
rect 3227 616 3273 756
rect 3431 787 3477 927
<< polysilicon >>
rect 124 933 224 977
rect 328 933 428 977
rect 660 933 760 977
rect 1058 940 1158 984
rect 1262 940 1362 984
rect 1466 940 1566 984
rect 1670 940 1770 984
rect 1874 940 1974 984
rect 2078 940 2178 984
rect 2282 940 2382 984
rect 2486 940 2586 984
rect 2690 940 2790 984
rect 2894 940 2994 984
rect 3098 940 3198 984
rect 3302 940 3402 984
rect 124 513 224 573
rect 328 513 428 573
rect 660 540 760 573
rect 124 487 612 513
rect 124 441 142 487
rect 188 473 612 487
rect 660 494 673 540
rect 719 494 760 540
rect 660 481 760 494
rect 1058 520 1158 580
rect 1262 520 1362 580
rect 1466 520 1566 580
rect 1670 520 1770 580
rect 188 441 244 473
rect 124 333 244 441
rect 348 412 468 425
rect 348 366 361 412
rect 407 366 468 412
rect 348 333 468 366
rect 572 377 612 473
rect 1058 480 1770 520
rect 1874 539 1974 580
rect 1874 493 1887 539
rect 1933 520 1974 539
rect 2078 539 2178 580
rect 2078 520 2105 539
rect 1933 493 2105 520
rect 2151 520 2178 539
rect 2282 539 2382 580
rect 2282 520 2309 539
rect 2151 493 2309 520
rect 2355 520 2382 539
rect 2486 539 2586 580
rect 2486 520 2513 539
rect 2355 493 2513 520
rect 2559 520 2586 539
rect 2690 539 2790 580
rect 2690 520 2718 539
rect 2559 493 2718 520
rect 2764 520 2790 539
rect 2894 539 2994 580
rect 2894 520 2922 539
rect 2764 493 2922 520
rect 2968 520 2994 539
rect 3098 520 3198 580
rect 3302 520 3402 580
rect 2968 493 3402 520
rect 1874 480 3402 493
rect 572 333 692 377
rect 1058 376 1098 480
rect 978 332 1098 376
rect 1202 332 1322 480
rect 1426 411 1546 480
rect 1426 365 1446 411
rect 1492 365 1546 411
rect 1426 332 1546 365
rect 1650 411 1770 480
rect 1650 365 1686 411
rect 1732 365 1770 411
rect 1650 332 1770 365
rect 1874 419 3562 432
rect 1874 373 1887 419
rect 1933 392 2134 419
rect 1933 373 1994 392
rect 1874 332 1994 373
rect 2098 373 2134 392
rect 2180 392 2361 419
rect 2180 373 2218 392
rect 2098 332 2218 373
rect 2322 373 2361 392
rect 2407 392 2582 419
rect 2407 373 2442 392
rect 2322 332 2442 373
rect 2546 373 2582 392
rect 2628 392 2808 419
rect 2628 373 2666 392
rect 2546 332 2666 373
rect 2770 373 2808 392
rect 2854 392 3562 419
rect 2854 373 2890 392
rect 2770 332 2890 373
rect 2994 332 3114 392
rect 3218 332 3338 392
rect 3442 332 3562 392
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 978 24 1098 68
rect 1202 24 1322 68
rect 1426 24 1546 68
rect 1650 24 1770 68
rect 1874 24 1994 68
rect 2098 24 2218 68
rect 2322 24 2442 68
rect 2546 24 2666 68
rect 2770 24 2890 68
rect 2994 24 3114 68
rect 3218 24 3338 68
rect 3442 24 3562 68
<< polycontact >>
rect 142 441 188 487
rect 673 494 719 540
rect 361 366 407 412
rect 1887 493 1933 539
rect 2105 493 2151 539
rect 2309 493 2355 539
rect 2513 493 2559 539
rect 2718 493 2764 539
rect 2922 493 2968 539
rect 1446 365 1492 411
rect 1686 365 1732 411
rect 1887 373 1933 419
rect 2134 373 2180 419
rect 2361 373 2407 419
rect 2582 373 2628 419
rect 2808 373 2854 419
<< metal1 >>
rect 0 927 3696 1098
rect 0 920 983 927
rect 0 918 253 920
rect 299 918 983 920
rect 253 769 299 780
rect 585 818 927 829
rect 49 726 95 737
rect 631 783 927 818
rect 585 667 631 678
rect 789 726 835 737
rect 49 320 95 586
rect 142 487 306 542
rect 188 441 306 487
rect 142 430 306 441
rect 361 494 673 540
rect 719 494 730 540
rect 361 412 407 494
rect 789 448 835 586
rect 361 309 407 366
rect 95 274 407 309
rect 629 402 835 448
rect 881 650 927 783
rect 1029 918 1391 927
rect 983 776 1029 787
rect 1437 918 1799 927
rect 1391 776 1437 787
rect 1845 918 2207 927
rect 2253 918 2615 927
rect 2207 870 2253 881
rect 2661 918 3023 927
rect 2615 870 2661 881
rect 3069 918 3431 927
rect 3023 870 3069 881
rect 1799 776 1845 787
rect 3477 918 3696 927
rect 3431 776 3477 787
rect 1595 755 1641 766
rect 881 639 1595 650
rect 881 593 1187 639
rect 1233 615 1595 639
rect 2003 756 3273 767
rect 2003 709 2411 756
rect 2049 663 2411 709
rect 1641 615 1933 628
rect 2003 616 2411 663
rect 2457 616 2819 756
rect 2865 616 3227 756
rect 1233 593 1933 615
rect 881 582 1933 593
rect 629 298 675 402
rect 881 356 927 582
rect 1887 550 1933 582
rect 1887 539 2979 550
rect 1933 493 2105 539
rect 2151 493 2309 539
rect 2355 493 2513 539
rect 2559 493 2718 539
rect 2764 493 2922 539
rect 2968 493 2979 539
rect 1887 482 2979 493
rect 49 263 407 274
rect 497 287 675 298
rect 543 217 675 287
rect 721 320 927 356
rect 1435 411 1762 430
rect 1435 365 1446 411
rect 1492 365 1686 411
rect 1732 365 1762 411
rect 1435 354 1762 365
rect 1887 419 2865 430
rect 1933 373 2134 419
rect 2180 373 2361 419
rect 2407 373 2582 419
rect 2628 373 2808 419
rect 2854 373 2865 419
rect 1887 365 2865 373
rect 767 310 927 320
rect 1887 298 1933 365
rect 3152 330 3273 616
rect 3152 319 3413 330
rect 721 263 767 274
rect 1127 287 1933 298
rect 1127 252 1575 287
rect 1127 228 1173 252
rect 543 182 1127 217
rect 543 171 1173 182
rect 273 128 319 139
rect 497 136 543 147
rect 1621 252 1933 287
rect 2023 273 2471 319
rect 2069 227 2471 273
rect 2023 179 2471 227
rect 2517 179 2919 319
rect 2965 179 3367 319
rect 2023 173 3413 179
rect 3367 168 3413 173
rect 3591 221 3637 232
rect 0 82 273 90
rect 1351 127 1397 138
rect 1575 136 1621 147
rect 854 90 865 125
rect 319 82 865 90
rect 0 79 865 82
rect 911 90 922 125
rect 911 81 1351 90
rect 1799 127 1845 138
rect 1397 81 1799 90
rect 2236 90 2247 127
rect 1845 81 2247 90
rect 2293 90 2304 127
rect 2684 90 2695 127
rect 2293 81 2695 90
rect 2741 90 2752 127
rect 3132 90 3143 127
rect 2741 81 3143 90
rect 3189 90 3200 127
rect 3189 81 3591 90
rect 3637 81 3696 90
rect 911 79 3696 81
rect 0 -90 3696 79
<< labels >>
flabel metal1 s 142 430 306 542 0 FreeSans 200 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1435 354 1762 430 0 FreeSans 200 0 0 0 I
port 2 nsew default input
flabel metal1 s 0 918 3696 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 3591 139 3637 232 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 2003 616 3273 767 0 FreeSans 200 0 0 0 Z
port 3 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 3152 330 3273 616 1 Z
port 3 nsew default output
rlabel metal1 s 3152 319 3413 330 1 Z
port 3 nsew default output
rlabel metal1 s 2023 173 3413 319 1 Z
port 3 nsew default output
rlabel metal1 s 3367 168 3413 173 1 Z
port 3 nsew default output
rlabel metal1 s 3431 870 3477 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3023 870 3069 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2615 870 2661 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2207 870 2253 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1799 870 1845 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1391 870 1437 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 983 870 1029 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 253 870 299 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3431 776 3477 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1799 776 1845 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1391 776 1437 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 983 776 1029 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 253 776 299 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 253 769 299 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3591 138 3637 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 138 319 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3591 127 3637 138 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1799 127 1845 138 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1351 127 1397 138 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 127 319 138 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3591 125 3637 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3132 125 3200 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2684 125 2752 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2236 125 2304 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1799 125 1845 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1351 125 1397 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 125 319 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3591 90 3637 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3132 90 3200 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2684 90 2752 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2236 90 2304 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1799 90 1845 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1351 90 1397 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 854 90 922 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 125 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3696 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3696 1008
string GDS_END 1356718
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1348266
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
