magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
use M1_NACTIVE$$203393068_64x8m81  M1_NACTIVE$$203393068_64x8m81_0
timestamp 1755005639
transform 1 0 14063 0 1 8159
box 0 0 1 1
use M1_NWELL$$204218412_64x8m81  M1_NWELL$$204218412_64x8m81_0
timestamp 1755005639
transform -1 0 25568 0 1 8086
box 0 0 1 1
use M1_NWELL$$204218412_64x8m81  M1_NWELL$$204218412_64x8m81_1
timestamp 1755005639
transform 1 0 2200 0 1 8086
box 0 0 1 1
use M1_PACTIVE$$204148780_64x8m81  M1_PACTIVE$$204148780_64x8m81_0
timestamp 1755005639
transform 1 0 11463 0 1 8159
box 0 0 1 1
use M1_PACTIVE$$204148780_64x8m81  M1_PACTIVE$$204148780_64x8m81_1
timestamp 1755005639
transform 1 0 21475 0 1 8159
box 0 0 1 1
use M1_PACTIVE$$204148780_64x8m81  M1_PACTIVE$$204148780_64x8m81_2
timestamp 1755005639
transform 1 0 4390 0 1 8159
box 0 0 1 1
use M1_PACTIVE$$204149804_64x8m81  M1_PACTIVE$$204149804_64x8m81_0
timestamp 1755005639
transform 1 0 15860 0 1 8159
box 0 0 1 1
use M1_POLY2$$204150828_64x8m81  M1_POLY2$$204150828_64x8m81_0
timestamp 1755005639
transform 1 0 9381 0 1 7848
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_0
timestamp 1755005639
transform 1 0 15413 0 1 8141
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_0
timestamp 1755005639
transform 0 -1 13712 1 0 8093
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_1
timestamp 1755005639
transform 1 0 15625 0 1 7801
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_2
timestamp 1755005639
transform 1 0 18313 0 1 7836
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_3
timestamp 1755005639
transform 1 0 12040 0 1 7761
box 0 0 1 1
use M2_M1$$201262124_64x8m81  M2_M1$$201262124_64x8m81_0
timestamp 1755005639
transform 1 0 13701 0 1 8091
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_0
timestamp 1755005639
transform 1 0 13284 0 1 3362
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_1
timestamp 1755005639
transform 1 0 13284 0 1 5162
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_2
timestamp 1755005639
transform 1 0 13284 0 1 6962
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_3
timestamp 1755005639
transform 1 0 14794 0 1 5869
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_4
timestamp 1755005639
transform 1 0 14794 0 1 4931
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_5
timestamp 1755005639
transform 1 0 14794 0 1 4069
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_6
timestamp 1755005639
transform 1 0 14794 0 1 3131
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_7
timestamp 1755005639
transform 1 0 14794 0 1 2269
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_8
timestamp 1755005639
transform 1 0 14794 0 1 1331
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_9
timestamp 1755005639
transform 1 0 14794 0 1 469
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_10
timestamp 1755005639
transform 1 0 13284 0 1 2038
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_11
timestamp 1755005639
transform 1 0 13284 0 1 1562
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_12
timestamp 1755005639
transform 1 0 13284 0 1 238
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_13
timestamp 1755005639
transform 1 0 13284 0 1 5638
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_14
timestamp 1755005639
transform 1 0 13284 0 1 3838
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_15
timestamp 1755005639
transform 1 0 19590 0 1 578
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_16
timestamp 1755005639
transform 1 0 19213 0 1 1222
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_17
timestamp 1755005639
transform 1 0 18835 0 1 2378
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_18
timestamp 1755005639
transform 1 0 18457 0 1 3022
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_19
timestamp 1755005639
transform 1 0 18080 0 1 4178
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_20
timestamp 1755005639
transform 1 0 17702 0 1 4822
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_21
timestamp 1755005639
transform 1 0 17324 0 1 5978
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_22
timestamp 1755005639
transform 1 0 16946 0 1 6622
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_23
timestamp 1755005639
transform 1 0 14794 0 1 6731
box 0 0 1 1
use M2_M1$$204138540_64x8m81  M2_M1$$204138540_64x8m81_0
timestamp 1755005639
transform 1 0 10402 0 1 7848
box 0 0 1 1
use M2_M1$$204138540_64x8m81  M2_M1$$204138540_64x8m81_1
timestamp 1755005639
transform 1 0 14059 0 1 8152
box 0 0 1 1
use M2_M1$$204139564_64x8m81  M2_M1$$204139564_64x8m81_0
timestamp 1755005639
transform 1 0 11601 0 1 8105
box 0 0 1 1
use M2_M1$$204140588_64x8m81  M2_M1$$204140588_64x8m81_0
timestamp 1755005639
transform 1 0 12359 0 1 7617
box 0 0 1 1
use M2_M1$$204141612_64x8m81  M2_M1$$204141612_64x8m81_0
timestamp 1755005639
transform 1 0 15126 0 1 8152
box 0 0 1 1
use M2_M1$$204141612_64x8m81  M2_M1$$204141612_64x8m81_1
timestamp 1755005639
transform 1 0 20177 0 1 8080
box 0 0 1 1
use M2_M1$$204141612_64x8m81  M2_M1$$204141612_64x8m81_2
timestamp 1755005639
transform 1 0 20177 0 1 7617
box 0 0 1 1
use M2_M1$$204220460_64x8m81  M2_M1$$204220460_64x8m81_0
timestamp 1755005639
transform 1 0 6792 0 1 7617
box 0 0 1 1
use M2_M1$$204220460_64x8m81  M2_M1$$204220460_64x8m81_1
timestamp 1755005639
transform 1 0 22430 0 1 7617
box 0 0 1 1
use M2_M1$$204220460_64x8m81  M2_M1$$204220460_64x8m81_2
timestamp 1755005639
transform 1 0 4399 0 1 7619
box 0 0 1 1
use M2_M1$$204220460_64x8m81  M2_M1$$204220460_64x8m81_3
timestamp 1755005639
transform 1 0 6792 0 1 8080
box 0 0 1 1
use M2_M1$$204221484_64x8m81  M2_M1$$204221484_64x8m81_0
timestamp 1755005639
transform -1 0 25612 0 1 8100
box 0 0 1 1
use M2_M1$$204221484_64x8m81  M2_M1$$204221484_64x8m81_1
timestamp 1755005639
transform 1 0 2156 0 1 8100
box 0 0 1 1
use M2_M1$$204222508_64x8m81  M2_M1$$204222508_64x8m81_0
timestamp 1755005639
transform 1 0 21486 0 1 8100
box 0 0 1 1
use M2_M1$$204222508_64x8m81  M2_M1$$204222508_64x8m81_1
timestamp 1755005639
transform 1 0 5639 0 1 8100
box 0 0 1 1
use M3_M2$$204142636_64x8m81  M3_M2$$204142636_64x8m81_0
timestamp 1755005639
transform 1 0 5639 0 1 8100
box 0 0 1 1
use M3_M2$$204142636_64x8m81  M3_M2$$204142636_64x8m81_1
timestamp 1755005639
transform 1 0 8250 0 1 7617
box 0 0 1 1
use M3_M2$$204142636_64x8m81  M3_M2$$204142636_64x8m81_2
timestamp 1755005639
transform 1 0 21486 0 1 8100
box 0 0 1 1
use M3_M2$$204143660_64x8m81  M3_M2$$204143660_64x8m81_0
timestamp 1755005639
transform 1 0 11601 0 1 8100
box 0 0 1 1
use M3_M2$$204144684_64x8m81  M3_M2$$204144684_64x8m81_0
timestamp 1755005639
transform 1 0 22430 0 1 7617
box 0 0 1 1
use M3_M2$$204144684_64x8m81  M3_M2$$204144684_64x8m81_1
timestamp 1755005639
transform 1 0 4399 0 1 7619
box 0 0 1 1
use M3_M2$$204145708_64x8m81  M3_M2$$204145708_64x8m81_0
timestamp 1755005639
transform 1 0 12359 0 1 7617
box 0 0 1 1
use M3_M2$$204146732_64x8m81  M3_M2$$204146732_64x8m81_0
timestamp 1755005639
transform 1 0 14059 0 1 7610
box 0 0 1 1
use M3_M2$$204147756_64x8m81  M3_M2$$204147756_64x8m81_0
timestamp 1755005639
transform 1 0 12339 0 1 7200
box 0 0 1 1
use nmos_1p2$$204215_R270_64x8m81  nmos_1p2$$204215_R270_64x8m81_0
timestamp 1755005639
transform 0 -1 13604 -1 0 7762
box -31 0 -30 1
use nmos_1p2$$204213292_R90_64x8m81  nmos_1p2$$204213292_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 6346 1 0 7703
box -31 0 -30 1
use nmos_5p04310589983299_64x8m81  nmos_5p04310589983299_64x8m81_0
timestamp 1755005639
transform 0 -1 23346 1 0 7672
box 0 0 1 1
use nmos_5p043105899832103_64x8m81  nmos_5p043105899832103_64x8m81_0
timestamp 1755005639
transform 0 -1 16283 1 0 7672
box 0 0 1 1
use nmos_5p043105899832103_64x8m81  nmos_5p043105899832103_64x8m81_1
timestamp 1755005639
transform 0 -1 11913 1 0 7672
box 0 0 1 1
use pmos_1p2$$204216364_R90_64x8m81  pmos_1p2$$204216364_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 20950 1 0 7703
box -31 0 -30 1
use pmos_1p2$$204216364_R90_64x8m81  pmos_1p2$$204216364_R90_64x8m81_1
timestamp 1755005639
transform 0 -1 9245 1 0 7703
box -31 0 -30 1
use pmos_1p2$$204217388_R90_64x8m81  pmos_1p2$$204217388_R90_64x8m81_0
timestamp 1755005639
transform 0 -1 11004 1 0 7703
box -31 0 -30 1
use pmos_5p043105899832101_64x8m81  pmos_5p043105899832101_64x8m81_0
timestamp 1755005639
transform 0 -1 15304 1 0 7672
box 0 0 1 1
use pmos_5p043105899832101_64x8m81  pmos_5p043105899832101_64x8m81_1
timestamp 1755005639
transform 0 -1 17974 1 0 7672
box 0 0 1 1
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_0
timestamp 1755005639
transform 0 -1 2203 -1 0 7350
box 0 0 1 1
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_1
timestamp 1755005639
transform 0 -1 2203 -1 0 5550
box 0 0 1 1
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_2
timestamp 1755005639
transform 0 -1 2203 -1 0 3750
box 0 0 1 1
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_3
timestamp 1755005639
transform 0 -1 2203 -1 0 1950
box 0 0 1 1
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_4
timestamp 1755005639
transform 0 1 25566 -1 0 7350
box 0 0 1 1
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_5
timestamp 1755005639
transform 0 1 25566 -1 0 5550
box 0 0 1 1
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_6
timestamp 1755005639
transform 0 1 25566 -1 0 3750
box 0 0 1 1
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_7
timestamp 1755005639
transform 0 1 25566 -1 0 1950
box 0 0 1 1
use pmoscap_W2_5_R270_64x8m81  pmoscap_W2_5_R270_64x8m81_0
timestamp 1755005639
transform 0 -1 2203 -1 0 8250
box 150 220 1051 2048
use pmoscap_W2_5_R270_64x8m81  pmoscap_W2_5_R270_64x8m81_1
timestamp 1755005639
transform 0 1 25566 -1 0 8250
box 150 220 1051 2048
use xdec8_64x8m81  xdec8_64x8m81_0
timestamp 1755005639
transform 1 0 1726 0 1 0
box 1426 -1 22889 7201
<< properties >>
string GDS_END 1864818
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1849418
<< end >>
