magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 542 1486
<< nmos >>
rect 120 209 176 385
rect 280 209 336 385
<< pmos >>
rect 120 1015 176 1191
rect 280 1015 336 1191
<< ndiff >>
rect 32 268 120 385
rect 32 222 45 268
rect 91 222 120 268
rect 32 209 120 222
rect 176 371 280 385
rect 176 325 205 371
rect 251 325 280 371
rect 176 209 280 325
rect 336 268 424 385
rect 336 222 365 268
rect 411 222 424 268
rect 336 209 424 222
<< pdiff >>
rect 32 1178 120 1191
rect 32 1132 45 1178
rect 91 1132 120 1178
rect 32 1015 120 1132
rect 176 1015 280 1191
rect 336 1075 424 1191
rect 336 1029 365 1075
rect 411 1029 424 1075
rect 336 1015 424 1029
<< ndiffc >>
rect 45 222 91 268
rect 205 325 251 371
rect 365 222 411 268
<< pdiffc >>
rect 45 1132 91 1178
rect 365 1029 411 1075
<< psubdiff >>
rect 28 87 428 100
rect 28 41 55 87
rect 401 41 428 87
rect 28 28 428 41
<< nsubdiff >>
rect 28 1359 428 1372
rect 28 1313 55 1359
rect 401 1313 428 1359
rect 28 1300 428 1313
<< psubdiffcont >>
rect 55 41 401 87
<< nsubdiffcont >>
rect 55 1313 401 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 120 716 176 1015
rect 280 716 336 1015
rect 32 703 176 716
rect 32 657 45 703
rect 91 657 176 703
rect 32 644 176 657
rect 224 703 336 716
rect 224 657 237 703
rect 283 657 336 703
rect 224 644 336 657
rect 120 385 176 644
rect 280 385 336 644
rect 120 165 176 209
rect 280 165 336 209
<< polycontact >>
rect 45 657 91 703
rect 237 657 283 703
<< metal1 >>
rect 0 1359 456 1400
rect 0 1313 55 1359
rect 401 1313 456 1359
rect 0 1178 456 1313
rect 0 1132 45 1178
rect 91 1132 456 1178
rect 42 703 94 1086
rect 42 657 45 703
rect 91 657 94 703
rect 42 314 94 657
rect 234 703 286 1086
rect 234 657 237 703
rect 283 657 286 703
rect 234 428 286 657
rect 362 1075 414 1086
rect 362 1029 365 1075
rect 411 1029 414 1075
rect 362 382 414 1029
rect 205 371 414 382
rect 251 325 414 371
rect 205 314 414 325
rect 0 222 45 268
rect 91 222 365 268
rect 411 222 456 268
rect 0 87 456 222
rect 0 41 55 87
rect 401 41 456 87
rect 0 0 456 41
<< labels >>
rlabel metal1 s 0 0 456 268 4 vss
port 3 nsew
rlabel metal1 s 0 1132 456 1400 4 vdd
port 5 nsew
rlabel metal1 s 362 314 414 1086 4 nq
port 7 nsew
rlabel metal1 s 42 314 94 1086 4 i0
port 9 nsew
rlabel metal1 s 234 428 286 1086 4 i1
port 11 nsew
<< end >>
