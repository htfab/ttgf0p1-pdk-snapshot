* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__ao21_4.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__ao21_4 VDD VNW VPW VSS Y A B C
X0 VSS a_332_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.3025p ps=1.605u w=1u l=0.28u
X1 a_28_440# B VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X2 Y a_332_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X3 a_172_68# A VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X4 a_332_68# C a_28_440# VNW pfet_03v3 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.28u
X5 Y a_332_68# VDD VNW pfet_03v3 ad=0.41745p pd=1.985u as=0.6072p ps=3.64u w=1.38u l=0.28u
X6 VDD a_332_68# Y VNW pfet_03v3 ad=0.6279p pd=3.67u as=0.3588p ps=1.9u w=1.38u l=0.28u
X7 VSS a_332_68# Y VPW nfet_03v3 ad=0.455p pd=2.91u as=0.26p ps=1.52u w=1u l=0.28u
X8 VSS C a_332_68# VPW nfet_03v3 ad=0.58p pd=2.16u as=0.26p ps=1.52u w=1u l=0.28u
X9 Y a_332_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X10 Y a_332_68# VSS VPW nfet_03v3 ad=0.3025p pd=1.605u as=0.58p ps=2.16u w=1u l=0.28u
X11 VDD a_332_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.41745p ps=1.985u w=1.38u l=0.28u
X12 VDD A a_28_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X13 a_332_68# B a_172_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

