VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO nor2_x1
  CLASS BLOCK ;
  FOREIGN nor2_x1 ;
  ORIGIN 0.430 0.000 ;
  SIZE 3.140 BY 7.430 ;
  PIN vss
    ANTENNADIFFAREA 2.370000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 2.280 1.340 ;
    END
  END vss
  PIN vdd
    ANTENNADIFFAREA 1.633000 ;
    PORT
      LAYER Nwell ;
        RECT -0.430 3.400 2.710 7.430 ;
      LAYER Metal1 ;
        RECT 0.000 5.660 2.280 7.000 ;
    END
  END vdd
  PIN nq
    ANTENNADIFFAREA 1.888000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.810 2.910 2.070 5.430 ;
        RECT 1.025 1.570 2.070 2.910 ;
    END
  END nq
  PIN i0
    ANTENNAGATEAREA 1.106000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.210 1.570 0.470 5.430 ;
    END
  END i0
  PIN i1
    ANTENNAGATEAREA 1.106000 ;
    PORT
      LAYER Metal1 ;
        RECT 1.170 3.140 1.430 5.430 ;
    END
  END i1
END nor2_x1
END LIBRARY

