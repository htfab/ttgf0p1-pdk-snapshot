magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 998 1486
<< nmos >>
rect 120 209 176 385
rect 280 209 336 385
rect 440 209 496 385
rect 644 209 700 584
<< pmos >>
rect 120 1015 176 1191
rect 280 1015 336 1191
rect 440 1015 496 1191
rect 644 776 700 1191
<< ndiff >>
rect 556 385 644 584
rect 32 371 120 385
rect 32 325 45 371
rect 91 325 120 371
rect 32 209 120 325
rect 176 268 280 385
rect 176 222 205 268
rect 251 222 280 268
rect 176 209 280 222
rect 336 371 440 385
rect 336 325 365 371
rect 411 325 440 371
rect 336 209 440 325
rect 496 268 644 385
rect 496 222 569 268
rect 615 222 644 268
rect 496 209 644 222
rect 700 571 788 584
rect 700 325 729 571
rect 775 325 788 571
rect 700 209 788 325
<< pdiff >>
rect 32 1075 120 1191
rect 32 1029 45 1075
rect 91 1029 120 1075
rect 32 1015 120 1029
rect 176 1015 280 1191
rect 336 1015 440 1191
rect 496 1178 644 1191
rect 496 1132 569 1178
rect 615 1132 644 1178
rect 496 1015 644 1132
rect 556 776 644 1015
rect 700 1055 788 1191
rect 700 809 729 1055
rect 775 809 788 1055
rect 700 776 788 809
<< ndiffc >>
rect 45 325 91 371
rect 205 222 251 268
rect 365 325 411 371
rect 569 222 615 268
rect 729 325 775 571
<< pdiffc >>
rect 45 1029 91 1075
rect 569 1132 615 1178
rect 729 809 775 1055
<< psubdiff >>
rect 28 87 884 100
rect 28 41 83 87
rect 829 41 884 87
rect 28 28 884 41
<< nsubdiff >>
rect 28 1359 884 1372
rect 28 1313 83 1359
rect 829 1313 884 1359
rect 28 1300 884 1313
<< psubdiffcont >>
rect 83 41 829 87
<< nsubdiffcont >>
rect 83 1313 829 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 644 1191 700 1235
rect 120 716 176 1015
rect 280 716 336 1015
rect 440 716 496 1015
rect 644 716 700 776
rect 32 703 176 716
rect 32 657 45 703
rect 91 657 176 703
rect 32 644 176 657
rect 224 703 336 716
rect 224 657 237 703
rect 283 657 336 703
rect 224 644 336 657
rect 384 703 496 716
rect 384 657 397 703
rect 443 657 496 703
rect 384 644 496 657
rect 544 703 700 716
rect 544 657 557 703
rect 603 657 700 703
rect 544 644 700 657
rect 120 385 176 644
rect 280 385 336 644
rect 440 385 496 644
rect 644 584 700 644
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
rect 644 165 700 209
<< polycontact >>
rect 45 657 91 703
rect 237 657 283 703
rect 397 657 443 703
rect 557 657 603 703
<< metal1 >>
rect 0 1359 912 1400
rect 0 1313 83 1359
rect 829 1313 912 1359
rect 0 1178 912 1313
rect 0 1132 569 1178
rect 615 1132 912 1178
rect 45 1075 606 1086
rect 91 1029 606 1075
rect 45 1018 606 1029
rect 42 703 94 972
rect 42 657 45 703
rect 91 657 94 703
rect 42 428 94 657
rect 234 703 286 972
rect 234 657 237 703
rect 283 657 286 703
rect 234 428 286 657
rect 394 703 446 972
rect 394 657 397 703
rect 443 657 446 703
rect 394 428 446 657
rect 554 703 606 1018
rect 554 657 557 703
rect 603 657 606 703
rect 554 382 606 657
rect 45 371 606 382
rect 91 325 365 371
rect 411 325 606 371
rect 45 314 606 325
rect 726 1055 778 1086
rect 726 809 729 1055
rect 775 809 778 1055
rect 726 571 778 809
rect 726 325 729 571
rect 775 325 778 571
rect 726 314 778 325
rect 0 222 205 268
rect 251 222 569 268
rect 615 222 912 268
rect 0 87 912 222
rect 0 41 83 87
rect 829 41 912 87
rect 0 0 912 41
<< labels >>
rlabel metal1 s 0 1132 912 1400 4 vdd
port 3 nsew
rlabel metal1 s 0 0 912 268 4 vss
port 5 nsew
rlabel metal1 s 42 428 94 972 4 i0
port 7 nsew
rlabel metal1 s 234 428 286 972 4 i1
port 9 nsew
rlabel metal1 s 394 428 446 972 4 i2
port 11 nsew
rlabel metal1 s 726 314 778 1086 4 q
port 13 nsew
<< end >>
