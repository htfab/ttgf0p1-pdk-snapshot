magic
tech gf180mcuD
magscale 1 5
timestamp 1755005639
use 018SRAM_strap1_64x8m81  018SRAM_strap1_64x8m81_0
timestamp 1755005639
transform 1 0 0 0 -1 0
box -34 -34 334 484
use 018SRAM_strap1_64x8m81  018SRAM_strap1_64x8m81_1
timestamp 1755005639
transform 1 0 0 0 1 0
box -34 -34 334 484
<< properties >>
string GDS_END 536842
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 536740
<< end >>
