magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 352 1094 870
<< pwell >>
rect -86 -86 1094 352
<< mvnmos >>
rect 137 69 257 232
rect 321 69 441 232
rect 545 69 665 232
rect 729 69 849 232
<< mvpmos >>
rect 137 472 237 715
rect 341 472 441 715
rect 545 472 645 715
rect 749 472 849 715
<< mvndiff >>
rect 49 134 137 232
rect 49 88 62 134
rect 108 88 137 134
rect 49 69 137 88
rect 257 69 321 232
rect 441 174 545 232
rect 441 128 470 174
rect 516 128 545 174
rect 441 69 545 128
rect 665 69 729 232
rect 849 142 937 232
rect 849 96 878 142
rect 924 96 937 142
rect 849 69 937 96
<< mvpdiff >>
rect 49 665 137 715
rect 49 525 62 665
rect 108 525 137 665
rect 49 472 137 525
rect 237 665 341 715
rect 237 619 266 665
rect 312 619 341 665
rect 237 472 341 619
rect 441 676 545 715
rect 441 630 470 676
rect 516 630 545 676
rect 441 472 545 630
rect 645 531 749 715
rect 645 485 674 531
rect 720 485 749 531
rect 645 472 749 485
rect 849 665 937 715
rect 849 525 878 665
rect 924 525 937 665
rect 849 472 937 525
<< mvndiffc >>
rect 62 88 108 134
rect 470 128 516 174
rect 878 96 924 142
<< mvpdiffc >>
rect 62 525 108 665
rect 266 619 312 665
rect 470 630 516 676
rect 674 485 720 531
rect 878 525 924 665
<< polysilicon >>
rect 137 715 237 760
rect 341 715 441 760
rect 545 715 645 760
rect 749 715 849 760
rect 137 415 237 472
rect 137 369 162 415
rect 208 369 237 415
rect 137 276 237 369
rect 341 366 441 472
rect 341 320 368 366
rect 414 320 441 366
rect 341 276 441 320
rect 137 232 257 276
rect 321 232 441 276
rect 545 351 645 472
rect 545 305 586 351
rect 632 305 645 351
rect 545 276 645 305
rect 749 412 849 472
rect 749 366 790 412
rect 836 366 849 412
rect 749 276 849 366
rect 545 232 665 276
rect 729 232 849 276
rect 137 24 257 69
rect 321 24 441 69
rect 545 24 665 69
rect 729 24 849 69
<< polycontact >>
rect 162 369 208 415
rect 368 320 414 366
rect 586 305 632 351
rect 790 366 836 412
<< metal1 >>
rect 0 724 1008 844
rect 51 665 119 676
rect 51 525 62 665
rect 108 552 119 665
rect 266 665 312 724
rect 266 608 312 619
rect 364 630 470 676
rect 516 665 935 676
rect 516 630 878 665
rect 364 629 878 630
rect 364 552 410 629
rect 108 525 410 552
rect 51 506 410 525
rect 470 531 778 542
rect 470 485 674 531
rect 720 485 778 531
rect 867 525 878 629
rect 924 525 935 665
rect 867 506 935 525
rect 470 476 778 485
rect 122 415 314 430
rect 122 369 162 415
rect 208 369 314 415
rect 122 354 314 369
rect 360 366 424 430
rect 122 217 201 354
rect 360 320 368 366
rect 414 320 424 366
rect 62 134 108 145
rect 360 110 424 320
rect 470 174 536 476
rect 516 128 536 174
rect 470 117 536 128
rect 584 351 648 430
rect 584 305 586 351
rect 632 305 648 351
rect 584 110 648 305
rect 696 412 909 430
rect 696 366 790 412
rect 836 366 909 412
rect 696 360 909 366
rect 696 110 760 360
rect 878 142 924 181
rect 62 60 108 88
rect 878 60 924 96
rect 0 -60 1008 60
<< labels >>
flabel metal1 s 360 110 424 430 0 FreeSans 400 0 0 0 B1
port 3 nsew default input
flabel metal1 s 122 354 314 430 0 FreeSans 400 0 0 0 B2
port 4 nsew default input
flabel metal1 s 0 724 1008 844 0 FreeSans 400 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 878 145 924 181 0 FreeSans 400 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 470 476 778 542 0 FreeSans 400 0 0 0 ZN
port 5 nsew default output
flabel metal1 s 584 110 648 430 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 696 360 909 430 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 696 110 760 360 1 A2
port 2 nsew default input
rlabel metal1 s 122 217 201 354 1 B2
port 4 nsew default input
rlabel metal1 s 470 117 536 476 1 ZN
port 5 nsew default output
rlabel metal1 s 266 608 312 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 878 60 924 145 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 62 60 108 145 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1008 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1008 784
string GDS_END 1264640
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1261234
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
