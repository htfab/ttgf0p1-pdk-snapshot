magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 2102 1094
<< pwell >>
rect -86 -86 2102 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1048 69 1168 333
rect 1272 69 1392 333
rect 1496 69 1616 333
rect 1720 69 1840 333
<< mvpmos >>
rect 144 573 244 939
rect 358 573 458 939
rect 582 573 682 939
rect 796 573 896 939
rect 1068 573 1168 939
rect 1292 573 1392 939
rect 1506 573 1606 939
rect 1720 573 1820 939
<< mvndiff >>
rect 36 287 124 333
rect 36 147 49 287
rect 95 147 124 287
rect 36 69 124 147
rect 244 287 348 333
rect 244 147 273 287
rect 319 147 348 287
rect 244 69 348 147
rect 468 287 572 333
rect 468 147 497 287
rect 543 147 572 287
rect 468 69 572 147
rect 692 287 796 333
rect 692 147 721 287
rect 767 147 796 287
rect 692 69 796 147
rect 916 287 1048 333
rect 916 147 945 287
rect 991 147 1048 287
rect 916 69 1048 147
rect 1168 287 1272 333
rect 1168 147 1197 287
rect 1243 147 1272 287
rect 1168 69 1272 147
rect 1392 185 1496 333
rect 1392 139 1421 185
rect 1467 139 1496 185
rect 1392 69 1496 139
rect 1616 287 1720 333
rect 1616 147 1645 287
rect 1691 147 1720 287
rect 1616 69 1720 147
rect 1840 287 1928 333
rect 1840 147 1869 287
rect 1915 147 1928 287
rect 1840 69 1928 147
<< mvpdiff >>
rect 56 861 144 939
rect 56 721 69 861
rect 115 721 144 861
rect 56 573 144 721
rect 244 573 358 939
rect 458 861 582 939
rect 458 721 507 861
rect 553 721 582 861
rect 458 573 582 721
rect 682 573 796 939
rect 896 861 1068 939
rect 896 721 993 861
rect 1039 721 1068 861
rect 896 573 1068 721
rect 1168 861 1292 939
rect 1168 721 1217 861
rect 1263 721 1292 861
rect 1168 573 1292 721
rect 1392 861 1506 939
rect 1392 721 1421 861
rect 1467 721 1506 861
rect 1392 573 1506 721
rect 1606 861 1720 939
rect 1606 721 1635 861
rect 1681 721 1720 861
rect 1606 573 1720 721
rect 1820 861 1908 939
rect 1820 721 1849 861
rect 1895 721 1908 861
rect 1820 573 1908 721
<< mvndiffc >>
rect 49 147 95 287
rect 273 147 319 287
rect 497 147 543 287
rect 721 147 767 287
rect 945 147 991 287
rect 1197 147 1243 287
rect 1421 139 1467 185
rect 1645 147 1691 287
rect 1869 147 1915 287
<< mvpdiffc >>
rect 69 721 115 861
rect 507 721 553 861
rect 993 721 1039 861
rect 1217 721 1263 861
rect 1421 721 1467 861
rect 1635 721 1681 861
rect 1849 721 1895 861
<< polysilicon >>
rect 144 939 244 983
rect 358 939 458 983
rect 582 939 682 983
rect 796 939 896 983
rect 1068 939 1168 983
rect 1292 939 1392 983
rect 1506 939 1606 983
rect 1720 939 1820 983
rect 144 500 244 573
rect 144 454 185 500
rect 231 454 244 500
rect 144 377 244 454
rect 358 513 458 573
rect 582 513 682 573
rect 358 500 682 513
rect 358 454 371 500
rect 417 454 682 500
rect 358 441 682 454
rect 358 377 468 441
rect 124 333 244 377
rect 348 333 468 377
rect 572 377 682 441
rect 796 500 896 573
rect 796 454 809 500
rect 855 454 896 500
rect 796 377 896 454
rect 1068 513 1168 573
rect 1292 513 1392 573
rect 1506 513 1606 573
rect 1720 513 1820 573
rect 1068 500 1820 513
rect 1068 454 1197 500
rect 1243 454 1421 500
rect 1467 454 1820 500
rect 1068 441 1820 454
rect 1068 377 1168 441
rect 572 333 692 377
rect 796 333 916 377
rect 1048 333 1168 377
rect 1272 333 1392 441
rect 1496 333 1616 441
rect 1720 377 1820 441
rect 1720 333 1840 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1048 25 1168 69
rect 1272 25 1392 69
rect 1496 25 1616 69
rect 1720 25 1840 69
<< polycontact >>
rect 185 454 231 500
rect 371 454 417 500
rect 809 454 855 500
rect 1197 454 1243 500
rect 1421 454 1467 500
<< metal1 >>
rect 0 918 2016 1098
rect 69 861 115 918
rect 69 710 115 721
rect 507 861 553 872
rect 993 861 1039 918
rect 553 721 947 726
rect 507 680 947 721
rect 993 710 1039 721
rect 1217 861 1263 872
rect 174 588 855 634
rect 174 500 242 588
rect 174 454 185 500
rect 231 454 242 500
rect 360 500 428 542
rect 360 454 371 500
rect 417 454 428 500
rect 478 500 855 588
rect 478 454 809 500
rect 478 443 855 454
rect 901 500 947 680
rect 1217 664 1263 721
rect 1421 861 1467 918
rect 1421 710 1467 721
rect 1635 861 1681 872
rect 1635 664 1681 721
rect 1849 861 1895 918
rect 1849 710 1895 721
rect 1217 618 1681 664
rect 901 454 1197 500
rect 1243 454 1421 500
rect 1467 454 1478 500
rect 901 394 947 454
rect 273 348 947 394
rect 49 287 95 298
rect 49 90 95 147
rect 273 287 319 348
rect 273 136 319 147
rect 497 287 543 298
rect 497 90 543 147
rect 721 287 767 348
rect 1524 318 1570 618
rect 1197 298 1570 318
rect 721 136 767 147
rect 945 287 991 298
rect 945 90 991 147
rect 1197 287 1691 298
rect 1243 242 1645 287
rect 1197 136 1243 147
rect 1421 185 1467 196
rect 1421 90 1467 139
rect 1645 136 1691 147
rect 1869 287 1915 298
rect 1869 90 1915 147
rect 0 -90 2016 90
<< labels >>
flabel metal1 s 360 454 428 542 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 174 588 855 634 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 0 918 2016 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 1869 196 1915 298 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 1635 664 1681 872 0 FreeSans 200 0 0 0 Z
port 3 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 478 454 855 588 1 A2
port 2 nsew default input
rlabel metal1 s 174 454 242 588 1 A2
port 2 nsew default input
rlabel metal1 s 478 443 855 454 1 A2
port 2 nsew default input
rlabel metal1 s 1217 664 1263 872 1 Z
port 3 nsew default output
rlabel metal1 s 1217 618 1681 664 1 Z
port 3 nsew default output
rlabel metal1 s 1524 318 1570 618 1 Z
port 3 nsew default output
rlabel metal1 s 1197 298 1570 318 1 Z
port 3 nsew default output
rlabel metal1 s 1197 242 1691 298 1 Z
port 3 nsew default output
rlabel metal1 s 1645 136 1691 242 1 Z
port 3 nsew default output
rlabel metal1 s 1197 136 1243 242 1 Z
port 3 nsew default output
rlabel metal1 s 1849 710 1895 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1421 710 1467 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 993 710 1039 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 69 710 115 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 945 196 991 298 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 497 196 543 298 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 49 196 95 298 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1869 90 1915 196 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1421 90 1467 196 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 196 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 196 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 196 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2016 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2016 1008
string GDS_END 275158
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 269938
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
