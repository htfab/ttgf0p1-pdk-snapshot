VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fill_w2
  CLASS BLOCK ;
  FOREIGN fill_w2 ;
  ORIGIN 0.430 0.000 ;
  SIZE 3.140 BY 7.430 ;
  PIN vdd
    PORT
      LAYER Metal1 ;
        RECT 0.000 5.660 2.280 7.000 ;
    END
  END vdd
  PIN vss
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 2.280 1.340 ;
    END
  END vss
  OBS
      LAYER Nwell ;
        RECT -0.430 3.400 2.710 7.430 ;
  END
END fill_w2
END LIBRARY

