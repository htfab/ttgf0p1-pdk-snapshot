VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO diode_w1
  CLASS BLOCK ;
  FOREIGN diode_w1 ;
  ORIGIN 0.430 0.000 ;
  SIZE 2.000 BY 7.430 ;
  PIN vdd
    ANTENNADIFFAREA 0.309600 ;
    PORT
      LAYER Nwell ;
        RECT -0.430 3.400 1.570 7.430 ;
      LAYER Metal1 ;
        RECT 0.000 5.660 1.140 7.000 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 0.309600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 1.140 1.340 ;
    END
  END vss
  PIN i
    ANTENNADIFFAREA 1.080000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.400 3.830 0.740 5.430 ;
        RECT 0.440 2.970 0.700 3.830 ;
        RECT 0.400 1.570 0.740 2.970 ;
    END
  END i
END diode_w1
END LIBRARY

