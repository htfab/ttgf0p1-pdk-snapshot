VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ht_io__brk5_vss_vdd_dvss_dvdd
  CLASS PAD ;
  FOREIGN gf180mcu_ht_io__brk5_vss_vdd_dvss_dvdd ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal5 ;
        RECT 4.000 246.000 5.000 253.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 4.000 318.000 5.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.000 246.000 5.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 4.000 318.000 5.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 4.000 246.000 5.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 4.000 318.000 5.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 318.000 1.000 325.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 1.000 253.000 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal5 ;
        RECT 0.000 254.000 5.000 261.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 310.000 5.000 317.000 ;
    END
  END VDD
  PIN DVSS
    PORT
      LAYER Metal5 ;
        RECT 0.000 70.000 5.000 85.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 86.000 5.000 101.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 102.000 5.000 117.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 126.000 5.000 133.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 198.000 5.000 205.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 230.000 5.000 245.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 286.000 5.000 293.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 302.000 5.000 309.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 342.000 5.000 348.390 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 326.000 5.000 333.000 ;
    END
  END DVSS
  PIN DVDD
    PORT
      LAYER Metal5 ;
        RECT 0.000 334.000 5.000 341.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 118.000 5.000 125.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 134.000 5.000 149.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 150.000 5.000 165.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 166.000 5.000 181.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 182.000 5.000 197.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 206.000 5.000 213.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 214.000 5.000 229.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 294.000 5.000 301.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 262.000 5.000 269.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 270.000 5.000 277.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 0.000 278.000 5.000 285.000 ;
    END
  END DVDD
  OBS
      LAYER Metal1 ;
        RECT -0.160 65.540 5.160 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 68.110 5.000 348.080 ;
      LAYER Metal3 ;
        RECT 1.300 317.700 3.700 325.000 ;
        RECT 1.000 253.300 4.000 317.700 ;
        RECT 1.300 246.000 3.700 253.300 ;
      LAYER Metal4 ;
        RECT 1.300 317.700 3.700 325.000 ;
        RECT 1.000 253.300 4.000 317.700 ;
        RECT 1.300 246.000 3.700 253.300 ;
      LAYER Metal5 ;
        RECT 1.500 317.500 3.500 325.000 ;
        RECT 1.000 253.500 4.000 317.500 ;
        RECT 1.500 246.000 3.500 253.500 ;
  END
END gf180mcu_ht_io__brk5_vss_vdd_dvss_dvdd
END LIBRARY

