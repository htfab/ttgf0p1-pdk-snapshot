magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 998 1486
<< nmos >>
rect 120 209 176 518
rect 280 209 336 518
rect 440 209 496 518
rect 600 209 656 518
<< pmos >>
rect 120 842 176 1191
rect 280 842 336 1191
rect 440 842 496 1191
rect 600 842 656 1191
<< ndiff >>
rect 32 488 120 518
rect 32 342 45 488
rect 91 342 120 488
rect 32 209 120 342
rect 176 209 280 518
rect 336 268 440 518
rect 336 222 365 268
rect 411 222 440 268
rect 336 209 440 222
rect 496 209 600 518
rect 656 488 744 518
rect 656 342 685 488
rect 731 342 744 488
rect 656 209 744 342
<< pdiff >>
rect 32 1178 120 1191
rect 32 1132 45 1178
rect 91 1132 120 1178
rect 32 842 120 1132
rect 176 1038 280 1191
rect 176 892 205 1038
rect 251 892 280 1038
rect 176 842 280 892
rect 336 1178 440 1191
rect 336 1132 365 1178
rect 411 1132 440 1178
rect 336 842 440 1132
rect 496 1038 600 1191
rect 496 892 525 1038
rect 571 892 600 1038
rect 496 842 600 892
rect 656 1178 744 1191
rect 656 1132 685 1178
rect 731 1132 744 1178
rect 656 842 744 1132
<< ndiffc >>
rect 45 342 91 488
rect 365 222 411 268
rect 685 342 731 488
<< pdiffc >>
rect 45 1132 91 1178
rect 205 892 251 1038
rect 365 1132 411 1178
rect 525 892 571 1038
rect 685 1132 731 1178
<< psubdiff >>
rect 28 87 884 100
rect 28 41 83 87
rect 829 41 884 87
rect 28 28 884 41
<< nsubdiff >>
rect 28 1359 884 1372
rect 28 1313 83 1359
rect 829 1313 884 1359
rect 28 1300 884 1313
<< psubdiffcont >>
rect 83 41 829 87
<< nsubdiffcont >>
rect 83 1313 829 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 600 1191 656 1235
rect 120 782 176 842
rect 32 769 176 782
rect 32 723 45 769
rect 91 723 176 769
rect 32 710 176 723
rect 120 518 176 710
rect 280 650 336 842
rect 440 782 496 842
rect 384 769 496 782
rect 384 723 397 769
rect 443 723 496 769
rect 384 710 496 723
rect 228 637 336 650
rect 228 591 241 637
rect 287 591 336 637
rect 228 578 336 591
rect 280 518 336 578
rect 440 518 496 710
rect 600 650 656 842
rect 600 637 682 650
rect 600 591 623 637
rect 669 591 682 637
rect 600 578 682 591
rect 600 518 656 578
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
rect 600 165 656 209
<< polycontact >>
rect 45 723 91 769
rect 397 723 443 769
rect 241 591 287 637
rect 623 591 669 637
<< metal1 >>
rect 0 1359 912 1400
rect 0 1313 83 1359
rect 829 1313 912 1359
rect 0 1178 912 1313
rect 0 1132 45 1178
rect 91 1132 365 1178
rect 411 1132 685 1178
rect 731 1132 912 1178
rect 42 769 94 1086
rect 42 723 45 769
rect 91 723 94 769
rect 42 545 94 723
rect 140 1038 251 1086
rect 140 892 205 1038
rect 140 881 251 892
rect 522 1038 574 1086
rect 522 892 525 1038
rect 571 892 574 1038
rect 140 780 192 881
rect 140 769 443 780
rect 140 723 397 769
rect 140 712 443 723
rect 140 499 192 712
rect 522 648 574 892
rect 241 637 574 648
rect 287 591 574 637
rect 241 580 574 591
rect 45 488 192 499
rect 91 342 192 488
rect 45 314 192 342
rect 522 499 574 580
rect 620 637 672 1086
rect 620 591 623 637
rect 669 591 672 637
rect 620 545 672 591
rect 522 488 731 499
rect 522 342 685 488
rect 522 314 731 342
rect 0 222 365 268
rect 411 222 912 268
rect 0 87 912 222
rect 0 41 83 87
rect 829 41 912 87
rect 0 0 912 41
<< labels >>
rlabel metal1 s 140 314 192 1086 4 q
port 3 nsew
rlabel metal1 s 0 1132 912 1400 4 vdd
port 5 nsew
rlabel metal1 s 0 0 912 268 4 vss
port 7 nsew
rlabel metal1 s 42 545 94 1086 4 nset
port 9 nsew
rlabel metal1 s 522 314 574 1086 4 nq
port 11 nsew
rlabel metal1 s 620 545 672 1086 4 nrst
port 13 nsew
<< end >>
