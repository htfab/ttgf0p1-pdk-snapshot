magic
tech gf180mcuD
magscale 1 5
timestamp 1751546430
<< nwell >>
rect -43 177 1051 435
<< pwell >>
rect -43 -43 1051 177
<< ndiff >>
rect 14 34 994 134
<< pdiff >>
rect 14 220 994 358
<< metal1 >>
rect 0 362 1008 422
rect 0 -30 1008 30
<< labels >>
flabel metal1 s 0 362 1008 422 0 FreeSans 200 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -30 1008 30 0 FreeSans 200 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 5 367 55 417 0 FreeSans 200 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 5 -25 55 25 0 FreeSans 200 0 0 0 VPW
port 3 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1008 392
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
