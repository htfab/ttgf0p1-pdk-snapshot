magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 352 2102 870
<< pwell >>
rect -86 -86 2102 352
<< metal1 >>
rect 0 724 2016 844
rect 49 510 95 724
rect 253 546 299 676
rect 466 593 534 724
rect 701 546 747 676
rect 914 593 982 724
rect 253 545 747 546
rect 1149 545 1195 676
rect 1362 593 1430 724
rect 1597 545 1643 676
rect 253 482 1643 545
rect 1821 510 1867 724
rect 126 353 758 430
rect 914 307 990 482
rect 1066 353 1792 430
rect 273 243 1663 307
rect 49 60 95 208
rect 273 140 319 243
rect 486 60 554 197
rect 721 140 767 243
rect 934 60 1002 197
rect 1169 140 1215 243
rect 1382 60 1450 197
rect 1617 140 1663 243
rect 1841 60 1887 208
rect 0 -60 2016 60
<< labels >>
rlabel metal1 s 1066 353 1792 430 6 I
port 1 nsew default input
rlabel metal1 s 126 353 758 430 6 I
port 1 nsew default input
rlabel metal1 s 1617 140 1663 243 6 ZN
port 2 nsew default output
rlabel metal1 s 1169 140 1215 243 6 ZN
port 2 nsew default output
rlabel metal1 s 721 140 767 243 6 ZN
port 2 nsew default output
rlabel metal1 s 273 140 319 243 6 ZN
port 2 nsew default output
rlabel metal1 s 273 243 1663 307 6 ZN
port 2 nsew default output
rlabel metal1 s 914 307 990 482 6 ZN
port 2 nsew default output
rlabel metal1 s 253 482 1643 545 6 ZN
port 2 nsew default output
rlabel metal1 s 1597 545 1643 676 6 ZN
port 2 nsew default output
rlabel metal1 s 1149 545 1195 676 6 ZN
port 2 nsew default output
rlabel metal1 s 253 545 747 546 6 ZN
port 2 nsew default output
rlabel metal1 s 701 546 747 676 6 ZN
port 2 nsew default output
rlabel metal1 s 253 546 299 676 6 ZN
port 2 nsew default output
rlabel metal1 s 1821 510 1867 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1362 593 1430 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 914 593 982 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 466 593 534 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 510 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 724 2016 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 352 2102 870 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 2102 352 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -60 2016 60 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1841 60 1887 208 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 197 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 197 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 197 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 208 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2016 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 831608
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 826404
<< end >>
