magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 998 1486
<< nmos >>
rect 120 209 176 584
rect 280 209 336 584
rect 440 209 496 584
rect 600 209 656 584
<< pmos >>
rect 120 776 176 1191
rect 280 776 336 1191
rect 440 776 496 1191
rect 600 776 656 1191
<< ndiff >>
rect 32 268 120 584
rect 32 222 45 268
rect 91 222 120 268
rect 32 209 120 222
rect 176 571 280 584
rect 176 325 205 571
rect 251 325 280 571
rect 176 209 280 325
rect 336 268 440 584
rect 336 222 365 268
rect 411 222 440 268
rect 336 209 440 222
rect 496 571 600 584
rect 496 325 525 571
rect 571 325 600 571
rect 496 209 600 325
rect 656 268 744 584
rect 656 222 685 268
rect 731 222 744 268
rect 656 209 744 222
<< pdiff >>
rect 32 1178 120 1191
rect 32 1132 45 1178
rect 91 1132 120 1178
rect 32 776 120 1132
rect 176 1055 280 1191
rect 176 809 205 1055
rect 251 809 280 1055
rect 176 776 280 809
rect 336 1178 440 1191
rect 336 1132 365 1178
rect 411 1132 440 1178
rect 336 776 440 1132
rect 496 1055 600 1191
rect 496 809 525 1055
rect 571 809 600 1055
rect 496 776 600 809
rect 656 1178 744 1191
rect 656 1132 685 1178
rect 731 1132 744 1178
rect 656 776 744 1132
<< ndiffc >>
rect 45 222 91 268
rect 205 325 251 571
rect 365 222 411 268
rect 525 325 571 571
rect 685 222 731 268
<< pdiffc >>
rect 45 1132 91 1178
rect 205 809 251 1055
rect 365 1132 411 1178
rect 525 809 571 1055
rect 685 1132 731 1178
<< psubdiff >>
rect 28 87 884 100
rect 28 41 83 87
rect 829 41 884 87
rect 28 28 884 41
<< nsubdiff >>
rect 28 1359 884 1372
rect 28 1313 83 1359
rect 829 1313 884 1359
rect 28 1300 884 1313
<< psubdiffcont >>
rect 83 41 829 87
<< nsubdiffcont >>
rect 83 1313 829 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 600 1191 656 1235
rect 120 716 176 776
rect 280 716 336 776
rect 440 716 496 776
rect 600 716 656 776
rect 32 703 656 716
rect 32 657 45 703
rect 91 657 656 703
rect 32 644 656 657
rect 120 584 176 644
rect 280 584 336 644
rect 440 584 496 644
rect 600 584 656 644
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
rect 600 165 656 209
<< polycontact >>
rect 45 657 91 703
<< metal1 >>
rect 0 1359 912 1400
rect 0 1313 83 1359
rect 829 1313 912 1359
rect 0 1178 912 1313
rect 0 1132 45 1178
rect 91 1132 365 1178
rect 411 1132 685 1178
rect 731 1132 912 1178
rect 42 703 94 1086
rect 42 657 45 703
rect 91 657 94 703
rect 42 314 94 657
rect 202 1055 254 1086
rect 202 809 205 1055
rect 251 809 254 1055
rect 525 1055 571 1086
rect 202 714 254 809
rect 522 809 525 866
rect 571 809 574 866
rect 522 714 574 809
rect 202 646 574 714
rect 202 571 254 646
rect 202 325 205 571
rect 251 325 254 571
rect 522 571 574 646
rect 522 514 525 571
rect 202 314 254 325
rect 571 514 574 571
rect 525 314 571 325
rect 0 222 45 268
rect 91 222 365 268
rect 411 222 685 268
rect 731 222 912 268
rect 0 87 912 222
rect 0 41 83 87
rect 829 41 912 87
rect 0 0 912 41
<< labels >>
rlabel metal1 s 0 0 912 268 4 vss
port 3 nsew
rlabel metal1 s 0 1132 912 1400 4 vdd
port 5 nsew
rlabel metal1 s 202 314 254 1086 4 nq
port 7 nsew
rlabel metal1 s 42 314 94 1086 4 i
port 9 nsew
<< end >>
