magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 7478 1094
<< pwell >>
rect -86 -86 7478 453
<< mvnmos >>
rect 124 68 244 332
rect 348 68 468 332
rect 572 68 692 332
rect 1008 69 1128 333
rect 1232 69 1352 333
rect 1456 69 1576 333
rect 1680 69 1800 333
rect 1904 69 2024 333
rect 2128 69 2248 333
rect 2352 69 2472 333
rect 2576 69 2696 333
rect 2800 69 2920 333
rect 3024 69 3144 333
rect 3284 68 3404 332
rect 3508 68 3628 332
rect 3732 68 3852 332
rect 3956 68 4076 332
rect 4180 68 4300 332
rect 4404 68 4524 332
rect 4628 68 4748 332
rect 4852 68 4972 332
rect 5076 68 5196 332
rect 5300 68 5420 332
rect 5524 68 5644 332
rect 5748 68 5868 332
rect 5972 68 6092 332
rect 6196 68 6316 332
rect 6420 68 6540 332
rect 6644 68 6764 332
rect 6868 68 6988 332
rect 7092 68 7212 332
<< mvpmos >>
rect 252 580 352 940
rect 456 580 556 940
rect 660 580 760 940
rect 1008 580 1108 940
rect 1232 580 1332 940
rect 1456 580 1556 940
rect 1680 580 1780 940
rect 1904 580 2004 940
rect 2128 580 2228 940
rect 2352 580 2452 940
rect 2576 580 2676 940
rect 2800 580 2900 940
rect 3024 580 3124 940
rect 3284 580 3384 940
rect 3508 580 3608 940
rect 3742 580 3842 940
rect 3956 580 4056 940
rect 4180 580 4280 940
rect 4404 580 4504 940
rect 4628 580 4728 940
rect 4852 580 4952 940
rect 5076 580 5176 940
rect 5300 580 5400 940
rect 5524 580 5624 940
rect 5748 580 5848 940
rect 5972 580 6072 940
rect 6196 580 6296 940
rect 6420 580 6520 940
rect 6644 580 6744 940
rect 6868 580 6968 940
rect 7092 580 7192 940
<< mvndiff >>
rect 36 287 124 332
rect 36 147 49 287
rect 95 147 124 287
rect 36 68 124 147
rect 244 221 348 332
rect 244 81 273 221
rect 319 81 348 221
rect 244 68 348 81
rect 468 287 572 332
rect 468 147 497 287
rect 543 147 572 287
rect 468 68 572 147
rect 692 319 780 332
rect 692 273 721 319
rect 767 273 780 319
rect 692 68 780 273
rect 920 128 1008 333
rect 920 82 933 128
rect 979 82 1008 128
rect 920 69 1008 82
rect 1128 320 1232 333
rect 1128 274 1157 320
rect 1203 274 1232 320
rect 1128 69 1232 274
rect 1352 128 1456 333
rect 1352 82 1381 128
rect 1427 82 1456 128
rect 1352 69 1456 82
rect 1576 320 1680 333
rect 1576 274 1605 320
rect 1651 274 1680 320
rect 1576 69 1680 274
rect 1800 128 1904 333
rect 1800 82 1829 128
rect 1875 82 1904 128
rect 1800 69 1904 82
rect 2024 193 2128 333
rect 2024 147 2053 193
rect 2099 147 2128 193
rect 2024 69 2128 147
rect 2248 280 2352 333
rect 2248 140 2277 280
rect 2323 140 2352 280
rect 2248 69 2352 140
rect 2472 287 2576 333
rect 2472 147 2501 287
rect 2547 147 2576 287
rect 2472 69 2576 147
rect 2696 287 2800 333
rect 2696 147 2725 287
rect 2771 147 2800 287
rect 2696 69 2800 147
rect 2920 287 3024 333
rect 2920 147 2949 287
rect 2995 147 3024 287
rect 2920 69 3024 147
rect 3144 332 3224 333
rect 3144 287 3284 332
rect 3144 147 3173 287
rect 3219 147 3284 287
rect 3144 69 3284 147
rect 3204 68 3284 69
rect 3404 287 3508 332
rect 3404 147 3433 287
rect 3479 147 3508 287
rect 3404 68 3508 147
rect 3628 287 3732 332
rect 3628 147 3657 287
rect 3703 147 3732 287
rect 3628 68 3732 147
rect 3852 273 3956 332
rect 3852 227 3881 273
rect 3927 227 3956 273
rect 3852 68 3956 227
rect 4076 133 4180 332
rect 4076 87 4105 133
rect 4151 87 4180 133
rect 4076 68 4180 87
rect 4300 319 4404 332
rect 4300 179 4329 319
rect 4375 179 4404 319
rect 4300 68 4404 179
rect 4524 133 4628 332
rect 4524 87 4553 133
rect 4599 87 4628 133
rect 4524 68 4628 87
rect 4748 319 4852 332
rect 4748 179 4777 319
rect 4823 179 4852 319
rect 4748 68 4852 179
rect 4972 133 5076 332
rect 4972 87 5001 133
rect 5047 87 5076 133
rect 4972 68 5076 87
rect 5196 319 5300 332
rect 5196 179 5225 319
rect 5271 179 5300 319
rect 5196 68 5300 179
rect 5420 133 5524 332
rect 5420 87 5449 133
rect 5495 87 5524 133
rect 5420 68 5524 87
rect 5644 319 5748 332
rect 5644 179 5673 319
rect 5719 179 5748 319
rect 5644 68 5748 179
rect 5868 133 5972 332
rect 5868 87 5897 133
rect 5943 87 5972 133
rect 5868 68 5972 87
rect 6092 319 6196 332
rect 6092 179 6121 319
rect 6167 179 6196 319
rect 6092 68 6196 179
rect 6316 133 6420 332
rect 6316 87 6345 133
rect 6391 87 6420 133
rect 6316 68 6420 87
rect 6540 319 6644 332
rect 6540 179 6569 319
rect 6615 179 6644 319
rect 6540 68 6644 179
rect 6764 133 6868 332
rect 6764 87 6793 133
rect 6839 87 6868 133
rect 6764 68 6868 87
rect 6988 272 7092 332
rect 6988 226 7017 272
rect 7063 226 7092 272
rect 6988 68 7092 226
rect 7212 287 7300 332
rect 7212 147 7241 287
rect 7287 147 7300 287
rect 7212 68 7300 147
<< mvpdiff >>
rect 164 813 252 940
rect 164 673 177 813
rect 223 673 252 813
rect 164 580 252 673
rect 352 813 456 940
rect 352 673 381 813
rect 427 673 456 813
rect 352 580 456 673
rect 556 813 660 940
rect 556 673 585 813
rect 631 673 660 813
rect 556 580 660 673
rect 760 719 848 940
rect 760 673 789 719
rect 835 673 848 719
rect 760 580 848 673
rect 920 927 1008 940
rect 920 881 933 927
rect 979 881 1008 927
rect 920 580 1008 881
rect 1108 719 1232 940
rect 1108 673 1157 719
rect 1203 673 1232 719
rect 1108 580 1232 673
rect 1332 927 1456 940
rect 1332 881 1361 927
rect 1407 881 1456 927
rect 1332 580 1456 881
rect 1556 719 1680 940
rect 1556 673 1605 719
rect 1651 673 1680 719
rect 1556 580 1680 673
rect 1780 813 1904 940
rect 1780 673 1809 813
rect 1855 673 1904 813
rect 1780 580 1904 673
rect 2004 813 2128 940
rect 2004 673 2033 813
rect 2079 673 2128 813
rect 2004 580 2128 673
rect 2228 813 2352 940
rect 2228 673 2257 813
rect 2303 673 2352 813
rect 2228 580 2352 673
rect 2452 813 2576 940
rect 2452 673 2481 813
rect 2527 673 2576 813
rect 2452 580 2576 673
rect 2676 813 2800 940
rect 2676 673 2705 813
rect 2751 673 2800 813
rect 2676 580 2800 673
rect 2900 813 3024 940
rect 2900 673 2929 813
rect 2975 673 3024 813
rect 2900 580 3024 673
rect 3124 813 3284 940
rect 3124 673 3153 813
rect 3199 673 3284 813
rect 3124 580 3284 673
rect 3384 813 3508 940
rect 3384 673 3413 813
rect 3459 673 3508 813
rect 3384 580 3508 673
rect 3608 927 3742 940
rect 3608 787 3637 927
rect 3683 787 3742 927
rect 3608 580 3742 787
rect 3842 813 3956 940
rect 3842 673 3881 813
rect 3927 673 3956 813
rect 3842 580 3956 673
rect 4056 900 4180 940
rect 4056 760 4085 900
rect 4131 760 4180 900
rect 4056 580 4180 760
rect 4280 813 4404 940
rect 4280 673 4309 813
rect 4355 673 4404 813
rect 4280 580 4404 673
rect 4504 900 4628 940
rect 4504 760 4533 900
rect 4579 760 4628 900
rect 4504 580 4628 760
rect 4728 813 4852 940
rect 4728 673 4757 813
rect 4803 673 4852 813
rect 4728 580 4852 673
rect 4952 900 5076 940
rect 4952 760 4981 900
rect 5027 760 5076 900
rect 4952 580 5076 760
rect 5176 813 5300 940
rect 5176 673 5205 813
rect 5251 673 5300 813
rect 5176 580 5300 673
rect 5400 900 5524 940
rect 5400 760 5429 900
rect 5475 760 5524 900
rect 5400 580 5524 760
rect 5624 813 5748 940
rect 5624 673 5653 813
rect 5699 673 5748 813
rect 5624 580 5748 673
rect 5848 900 5972 940
rect 5848 760 5877 900
rect 5923 760 5972 900
rect 5848 580 5972 760
rect 6072 813 6196 940
rect 6072 673 6101 813
rect 6147 673 6196 813
rect 6072 580 6196 673
rect 6296 900 6420 940
rect 6296 760 6325 900
rect 6371 760 6420 900
rect 6296 580 6420 760
rect 6520 813 6644 940
rect 6520 673 6549 813
rect 6595 673 6644 813
rect 6520 580 6644 673
rect 6744 900 6868 940
rect 6744 760 6773 900
rect 6819 760 6868 900
rect 6744 580 6868 760
rect 6968 813 7092 940
rect 6968 673 7017 813
rect 7063 673 7092 813
rect 6968 580 7092 673
rect 7192 813 7280 940
rect 7192 673 7221 813
rect 7267 673 7280 813
rect 7192 580 7280 673
<< mvndiffc >>
rect 49 147 95 287
rect 273 81 319 221
rect 497 147 543 287
rect 721 273 767 319
rect 933 82 979 128
rect 1157 274 1203 320
rect 1381 82 1427 128
rect 1605 274 1651 320
rect 1829 82 1875 128
rect 2053 147 2099 193
rect 2277 140 2323 280
rect 2501 147 2547 287
rect 2725 147 2771 287
rect 2949 147 2995 287
rect 3173 147 3219 287
rect 3433 147 3479 287
rect 3657 147 3703 287
rect 3881 227 3927 273
rect 4105 87 4151 133
rect 4329 179 4375 319
rect 4553 87 4599 133
rect 4777 179 4823 319
rect 5001 87 5047 133
rect 5225 179 5271 319
rect 5449 87 5495 133
rect 5673 179 5719 319
rect 5897 87 5943 133
rect 6121 179 6167 319
rect 6345 87 6391 133
rect 6569 179 6615 319
rect 6793 87 6839 133
rect 7017 226 7063 272
rect 7241 147 7287 287
<< mvpdiffc >>
rect 177 673 223 813
rect 381 673 427 813
rect 585 673 631 813
rect 789 673 835 719
rect 933 881 979 927
rect 1157 673 1203 719
rect 1361 881 1407 927
rect 1605 673 1651 719
rect 1809 673 1855 813
rect 2033 673 2079 813
rect 2257 673 2303 813
rect 2481 673 2527 813
rect 2705 673 2751 813
rect 2929 673 2975 813
rect 3153 673 3199 813
rect 3413 673 3459 813
rect 3637 787 3683 927
rect 3881 673 3927 813
rect 4085 760 4131 900
rect 4309 673 4355 813
rect 4533 760 4579 900
rect 4757 673 4803 813
rect 4981 760 5027 900
rect 5205 673 5251 813
rect 5429 760 5475 900
rect 5653 673 5699 813
rect 5877 760 5923 900
rect 6101 673 6147 813
rect 6325 760 6371 900
rect 6549 673 6595 813
rect 6773 760 6819 900
rect 7017 673 7063 813
rect 7221 673 7267 813
<< polysilicon >>
rect 252 940 352 984
rect 456 940 556 984
rect 660 940 760 984
rect 1008 940 1108 984
rect 1232 940 1332 984
rect 1456 940 1556 984
rect 1680 940 1780 984
rect 1904 940 2004 984
rect 2128 940 2228 984
rect 2352 940 2452 984
rect 2576 940 2676 984
rect 2800 940 2900 984
rect 3024 940 3124 984
rect 3284 940 3384 984
rect 3508 940 3608 984
rect 3742 940 3842 984
rect 3956 940 4056 984
rect 4180 940 4280 984
rect 4404 940 4504 984
rect 4628 940 4728 984
rect 4852 940 4952 984
rect 5076 940 5176 984
rect 5300 940 5400 984
rect 5524 940 5624 984
rect 5748 940 5848 984
rect 5972 940 6072 984
rect 6196 940 6296 984
rect 6420 940 6520 984
rect 6644 940 6744 984
rect 6868 940 6968 984
rect 7092 940 7192 984
rect 252 520 352 580
rect 456 520 556 580
rect 660 547 760 580
rect 252 480 612 520
rect 660 501 673 547
rect 719 501 760 547
rect 660 488 760 501
rect 1008 520 1108 580
rect 1232 520 1332 580
rect 1456 520 1556 580
rect 1680 520 1780 580
rect 1008 507 1780 520
rect 252 440 292 480
rect 124 427 292 440
rect 124 381 185 427
rect 231 400 292 427
rect 348 419 468 432
rect 231 381 244 400
rect 124 332 244 381
rect 348 373 361 419
rect 407 373 468 419
rect 348 332 468 373
rect 572 376 612 480
rect 1008 461 1026 507
rect 1542 461 1780 507
rect 1008 448 1780 461
rect 572 332 692 376
rect 1008 333 1128 448
rect 1232 447 1780 448
rect 1232 333 1352 447
rect 1456 377 1575 447
rect 1680 377 1780 447
rect 1904 520 2004 580
rect 2128 520 2228 580
rect 2352 520 2452 580
rect 2576 520 2676 580
rect 2800 520 2900 580
rect 3024 520 3124 580
rect 3284 520 3384 580
rect 3508 520 3608 580
rect 1904 507 3608 520
rect 1904 461 1917 507
rect 3279 461 3608 507
rect 3742 547 3842 580
rect 3742 501 3766 547
rect 3812 520 3842 547
rect 3956 547 4056 580
rect 3956 520 3984 547
rect 3812 501 3984 520
rect 4030 520 4056 547
rect 4180 547 4280 580
rect 4180 520 4209 547
rect 4030 501 4209 520
rect 4255 520 4280 547
rect 4404 547 4504 580
rect 4404 520 4431 547
rect 4255 501 4431 520
rect 4477 520 4504 547
rect 4628 547 4728 580
rect 4628 520 4656 547
rect 4477 501 4656 520
rect 4702 520 4728 547
rect 4852 547 4952 580
rect 4852 520 4881 547
rect 4702 501 4881 520
rect 4927 520 4952 547
rect 5076 547 5176 580
rect 5076 520 5105 547
rect 4927 501 5105 520
rect 5151 520 5176 547
rect 5300 547 5400 580
rect 5300 520 5325 547
rect 5151 501 5325 520
rect 5371 520 5400 547
rect 5524 547 5624 580
rect 5524 520 5549 547
rect 5371 501 5549 520
rect 5595 520 5624 547
rect 5748 547 5848 580
rect 5748 520 5776 547
rect 5595 501 5776 520
rect 5822 520 5848 547
rect 5972 547 6072 580
rect 5972 520 5999 547
rect 5822 501 5999 520
rect 6045 520 6072 547
rect 6196 547 6296 580
rect 6196 520 6223 547
rect 6045 501 6223 520
rect 6269 520 6296 547
rect 6420 547 6520 580
rect 6420 520 6447 547
rect 6269 501 6447 520
rect 6493 520 6520 547
rect 6644 547 6744 580
rect 6644 520 6670 547
rect 6493 501 6670 520
rect 6716 520 6744 547
rect 6868 520 6968 580
rect 7092 520 7192 580
rect 6716 501 7192 520
rect 3742 480 7192 501
rect 1904 448 3608 461
rect 1456 333 1576 377
rect 1680 333 1800 377
rect 1904 333 2024 448
rect 2128 333 2248 448
rect 2352 333 2472 448
rect 2576 333 2696 448
rect 2800 333 2920 448
rect 3024 333 3144 448
rect 3284 332 3404 448
rect 3508 376 3608 448
rect 3732 419 7212 432
rect 3508 332 3628 376
rect 3732 373 3768 419
rect 3814 392 3996 419
rect 3814 373 3852 392
rect 3732 332 3852 373
rect 3956 373 3996 392
rect 4042 392 4219 419
rect 4042 373 4076 392
rect 3956 332 4076 373
rect 4180 373 4219 392
rect 4265 392 4442 419
rect 4265 373 4300 392
rect 4180 332 4300 373
rect 4404 373 4442 392
rect 4488 392 4665 419
rect 4488 373 4524 392
rect 4404 332 4524 373
rect 4628 373 4665 392
rect 4711 392 4888 419
rect 4711 373 4748 392
rect 4628 332 4748 373
rect 4852 373 4888 392
rect 4934 392 5112 419
rect 4934 373 4972 392
rect 4852 332 4972 373
rect 5076 373 5112 392
rect 5158 392 5337 419
rect 5158 373 5196 392
rect 5076 332 5196 373
rect 5300 373 5337 392
rect 5383 392 5561 419
rect 5383 373 5420 392
rect 5300 332 5420 373
rect 5524 373 5561 392
rect 5607 392 5785 419
rect 5607 373 5644 392
rect 5524 332 5644 373
rect 5748 373 5785 392
rect 5831 392 6007 419
rect 5831 373 5868 392
rect 5748 332 5868 373
rect 5972 373 6007 392
rect 6053 392 6234 419
rect 6053 373 6092 392
rect 5972 332 6092 373
rect 6196 373 6234 392
rect 6280 392 6457 419
rect 6280 373 6316 392
rect 6196 332 6316 373
rect 6420 373 6457 392
rect 6503 392 6680 419
rect 6503 373 6540 392
rect 6420 332 6540 373
rect 6644 373 6680 392
rect 6726 392 7212 419
rect 6726 373 6764 392
rect 6644 332 6764 373
rect 6868 332 6988 392
rect 7092 332 7212 392
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 1008 25 1128 69
rect 1232 25 1352 69
rect 1456 25 1576 69
rect 1680 25 1800 69
rect 1904 25 2024 69
rect 2128 25 2248 69
rect 2352 25 2472 69
rect 2576 25 2696 69
rect 2800 25 2920 69
rect 3024 25 3144 69
rect 3284 24 3404 68
rect 3508 24 3628 68
rect 3732 24 3852 68
rect 3956 24 4076 68
rect 4180 24 4300 68
rect 4404 24 4524 68
rect 4628 24 4748 68
rect 4852 24 4972 68
rect 5076 24 5196 68
rect 5300 24 5420 68
rect 5524 24 5644 68
rect 5748 24 5868 68
rect 5972 24 6092 68
rect 6196 24 6316 68
rect 6420 24 6540 68
rect 6644 24 6764 68
rect 6868 24 6988 68
rect 7092 24 7212 68
<< polycontact >>
rect 673 501 719 547
rect 185 381 231 427
rect 361 373 407 419
rect 1026 461 1542 507
rect 1917 461 3279 507
rect 3766 501 3812 547
rect 3984 501 4030 547
rect 4209 501 4255 547
rect 4431 501 4477 547
rect 4656 501 4702 547
rect 4881 501 4927 547
rect 5105 501 5151 547
rect 5325 501 5371 547
rect 5549 501 5595 547
rect 5776 501 5822 547
rect 5999 501 6045 547
rect 6223 501 6269 547
rect 6447 501 6493 547
rect 6670 501 6716 547
rect 3768 373 3814 419
rect 3996 373 4042 419
rect 4219 373 4265 419
rect 4442 373 4488 419
rect 4665 373 4711 419
rect 4888 373 4934 419
rect 5112 373 5158 419
rect 5337 373 5383 419
rect 5561 373 5607 419
rect 5785 373 5831 419
rect 6007 373 6053 419
rect 6234 373 6280 419
rect 6457 373 6503 419
rect 6680 373 6726 419
<< metal1 >>
rect 0 927 7392 1098
rect 0 918 933 927
rect 177 813 223 824
rect 177 547 223 673
rect 381 813 427 918
rect 979 918 1361 927
rect 933 870 979 881
rect 1407 918 3637 927
rect 1361 870 1407 881
rect 381 662 427 673
rect 585 813 1763 824
rect 631 778 1763 813
rect 585 662 631 673
rect 789 719 835 730
rect 177 501 673 547
rect 719 501 730 547
rect 163 427 231 455
rect 163 381 185 427
rect 163 370 231 381
rect 361 419 407 501
rect 789 419 835 673
rect 361 324 407 373
rect 49 287 407 324
rect 618 373 835 419
rect 618 298 664 373
rect 881 319 927 778
rect 1146 719 1662 730
rect 1146 673 1157 719
rect 1203 673 1605 719
rect 1651 673 1662 719
rect 1146 662 1662 673
rect 1616 524 1662 662
rect 1717 616 1763 778
rect 1809 813 1855 918
rect 1809 662 1855 673
rect 2033 813 2079 824
rect 2033 616 2079 673
rect 2257 813 2303 918
rect 2257 662 2303 673
rect 2481 813 2527 824
rect 2481 616 2527 673
rect 2705 813 2751 918
rect 2705 662 2751 673
rect 2929 813 2975 824
rect 2929 616 2975 673
rect 3153 813 3199 918
rect 3153 662 3199 673
rect 3413 813 3459 824
rect 3683 918 7392 927
rect 4085 900 4131 918
rect 3637 776 3683 787
rect 3881 813 3927 824
rect 3413 616 3459 673
rect 1717 570 3459 616
rect 4533 900 4579 918
rect 4085 749 4131 760
rect 4309 813 4355 824
rect 4981 900 5027 918
rect 4533 749 4579 760
rect 4757 813 4803 824
rect 5429 900 5475 918
rect 4981 749 5027 760
rect 5205 813 5251 824
rect 5877 900 5923 918
rect 5429 749 5475 760
rect 5653 813 5699 824
rect 6325 900 6371 918
rect 5877 749 5923 760
rect 6101 813 6147 824
rect 6773 900 6819 918
rect 6325 749 6371 760
rect 6549 813 6595 824
rect 6773 749 6819 760
rect 7017 813 7063 824
rect 3881 593 7063 673
rect 7221 813 7267 918
rect 7221 662 7267 673
rect 3413 547 3459 570
rect 1013 507 1542 521
rect 1013 461 1026 507
rect 1013 406 1542 461
rect 1616 507 3290 524
rect 1616 461 1917 507
rect 3279 461 3290 507
rect 3413 501 3766 547
rect 3812 501 3984 547
rect 4030 501 4209 547
rect 4255 501 4431 547
rect 4477 501 4656 547
rect 4702 501 4881 547
rect 4927 501 5105 547
rect 5151 501 5325 547
rect 5371 501 5549 547
rect 5595 501 5776 547
rect 5822 501 5999 547
rect 6045 501 6223 547
rect 6269 501 6447 547
rect 6493 501 6670 547
rect 6716 501 6740 547
rect 1616 320 1662 461
rect 3722 415 3768 419
rect 95 278 407 287
rect 497 287 664 298
rect 49 136 95 147
rect 273 221 319 232
rect 0 81 273 90
rect 543 227 664 287
rect 710 273 721 319
rect 767 273 927 319
rect 1146 274 1157 320
rect 1203 274 1605 320
rect 1651 274 1662 320
rect 2054 373 3768 415
rect 3814 373 3996 419
rect 4042 373 4219 419
rect 4265 373 4442 419
rect 4488 373 4665 419
rect 4711 373 4888 419
rect 4934 373 5112 419
rect 5158 373 5337 419
rect 5383 373 5561 419
rect 5607 373 5785 419
rect 5831 373 6007 419
rect 6053 373 6234 419
rect 6280 373 6457 419
rect 6503 373 6680 419
rect 6726 373 6746 419
rect 2054 350 3760 373
rect 2054 227 2100 350
rect 543 193 2100 227
rect 543 181 2053 193
rect 497 136 543 147
rect 2099 147 2100 193
rect 2053 136 2100 147
rect 2277 280 2323 291
rect 922 90 933 128
rect 319 82 933 90
rect 979 90 990 128
rect 1370 90 1381 128
rect 979 82 1381 90
rect 1427 90 1438 128
rect 1818 90 1829 128
rect 1427 82 1829 90
rect 1875 90 1886 128
rect 2277 90 2323 140
rect 2501 287 2547 350
rect 2501 136 2547 147
rect 2725 287 2771 298
rect 2725 90 2771 147
rect 2949 287 2995 350
rect 2949 136 2995 147
rect 3173 287 3219 298
rect 3173 90 3219 147
rect 3433 287 3479 350
rect 6967 319 7063 593
rect 3433 136 3479 147
rect 3657 287 3703 298
rect 3881 273 4329 319
rect 3927 227 4329 273
rect 3881 179 4329 227
rect 4375 179 4777 319
rect 4823 179 5225 319
rect 5271 179 5673 319
rect 5719 179 6121 319
rect 6167 179 6569 319
rect 6615 272 7063 319
rect 6615 226 7017 272
rect 6615 179 7063 226
rect 7241 287 7287 298
rect 3657 90 3703 147
rect 4094 90 4105 133
rect 1875 87 4105 90
rect 4151 90 4162 133
rect 4542 90 4553 133
rect 4151 87 4553 90
rect 4599 90 4610 133
rect 4990 90 5001 133
rect 4599 87 5001 90
rect 5047 90 5058 133
rect 5438 90 5449 133
rect 5047 87 5449 90
rect 5495 90 5506 133
rect 5886 90 5897 133
rect 5495 87 5897 90
rect 5943 90 5954 133
rect 6334 90 6345 133
rect 5943 87 6345 90
rect 6391 90 6402 133
rect 6782 90 6793 133
rect 6391 87 6793 90
rect 6839 90 6850 133
rect 7241 90 7287 147
rect 6839 87 7392 90
rect 1875 82 7392 87
rect 319 81 7392 82
rect 0 -90 7392 81
<< labels >>
flabel metal1 s 163 370 231 455 0 FreeSans 200 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1013 406 1542 521 0 FreeSans 200 0 0 0 I
port 2 nsew default input
flabel metal1 s 0 918 7392 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 7241 291 7287 298 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 7017 673 7063 824 0 FreeSans 200 0 0 0 ZN
port 3 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 6549 673 6595 824 1 ZN
port 3 nsew default output
rlabel metal1 s 6101 673 6147 824 1 ZN
port 3 nsew default output
rlabel metal1 s 5653 673 5699 824 1 ZN
port 3 nsew default output
rlabel metal1 s 5205 673 5251 824 1 ZN
port 3 nsew default output
rlabel metal1 s 4757 673 4803 824 1 ZN
port 3 nsew default output
rlabel metal1 s 4309 673 4355 824 1 ZN
port 3 nsew default output
rlabel metal1 s 3881 673 3927 824 1 ZN
port 3 nsew default output
rlabel metal1 s 3881 593 7063 673 1 ZN
port 3 nsew default output
rlabel metal1 s 6967 319 7063 593 1 ZN
port 3 nsew default output
rlabel metal1 s 3881 179 7063 319 1 ZN
port 3 nsew default output
rlabel metal1 s 7221 870 7267 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6773 870 6819 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6325 870 6371 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5877 870 5923 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5429 870 5475 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4981 870 5027 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4533 870 4579 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4085 870 4131 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3637 870 3683 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3153 870 3199 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2705 870 2751 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2257 870 2303 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1809 870 1855 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1361 870 1407 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 933 870 979 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 381 870 427 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 7221 776 7267 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6773 776 6819 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6325 776 6371 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5877 776 5923 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5429 776 5475 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4981 776 5027 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4533 776 4579 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4085 776 4131 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3637 776 3683 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3153 776 3199 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2705 776 2751 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2257 776 2303 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1809 776 1855 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 381 776 427 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 7221 749 7267 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6773 749 6819 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6325 749 6371 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5877 749 5923 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5429 749 5475 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4981 749 5027 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4533 749 4579 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4085 749 4131 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3153 749 3199 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2705 749 2751 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2257 749 2303 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1809 749 1855 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 381 749 427 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 7221 662 7267 749 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3153 662 3199 749 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2705 662 2751 749 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2257 662 2303 749 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1809 662 1855 749 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 381 662 427 749 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3657 291 3703 298 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3173 291 3219 298 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2725 291 2771 298 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 7241 232 7287 291 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3657 232 3703 291 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3173 232 3219 291 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2725 232 2771 291 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2277 232 2323 291 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 7241 133 7287 232 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3657 133 3703 232 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3173 133 3219 232 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2725 133 2771 232 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2277 133 2323 232 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 133 319 232 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 7241 128 7287 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 6782 128 6850 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 6334 128 6402 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5886 128 5954 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5438 128 5506 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4990 128 5058 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4542 128 4610 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4094 128 4162 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3657 128 3703 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3173 128 3219 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2725 128 2771 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2277 128 2323 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 128 319 133 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 7241 90 7287 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 6782 90 6850 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 6334 90 6402 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5886 90 5954 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5438 90 5506 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4990 90 5058 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4542 90 4610 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4094 90 4162 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3657 90 3703 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3173 90 3219 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2725 90 2771 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2277 90 2323 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1818 90 1886 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1370 90 1438 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 922 90 990 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 128 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 7392 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 7392 1008
string GDS_END 982694
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 966034
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
