magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 770 1486
<< nmos >>
rect 120 209 176 385
rect 280 209 336 385
rect 484 209 540 584
<< pmos >>
rect 120 1015 176 1191
rect 280 1015 336 1191
rect 484 776 540 1191
<< ndiff >>
rect 396 385 484 584
rect 32 268 120 385
rect 32 222 45 268
rect 91 222 120 268
rect 32 209 120 222
rect 176 371 280 385
rect 176 325 205 371
rect 251 325 280 371
rect 176 209 280 325
rect 336 268 484 385
rect 336 222 409 268
rect 455 222 484 268
rect 336 209 484 222
rect 540 571 628 584
rect 540 325 569 571
rect 615 325 628 571
rect 540 209 628 325
<< pdiff >>
rect 32 1075 120 1191
rect 32 1029 45 1075
rect 91 1029 120 1075
rect 32 1015 120 1029
rect 176 1015 280 1191
rect 336 1178 484 1191
rect 336 1132 409 1178
rect 455 1132 484 1178
rect 336 1015 484 1132
rect 396 776 484 1015
rect 540 1055 628 1191
rect 540 809 569 1055
rect 615 809 628 1055
rect 540 776 628 809
<< ndiffc >>
rect 45 222 91 268
rect 205 325 251 371
rect 409 222 455 268
rect 569 325 615 571
<< pdiffc >>
rect 45 1029 91 1075
rect 409 1132 455 1178
rect 569 809 615 1055
<< psubdiff >>
rect 28 87 656 100
rect 28 41 69 87
rect 615 41 656 87
rect 28 28 656 41
<< nsubdiff >>
rect 28 1359 656 1372
rect 28 1313 69 1359
rect 615 1313 656 1359
rect 28 1300 656 1313
<< psubdiffcont >>
rect 69 41 615 87
<< nsubdiffcont >>
rect 69 1313 615 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 484 1191 540 1235
rect 120 716 176 1015
rect 280 716 336 1015
rect 484 716 540 776
rect 32 703 176 716
rect 32 657 45 703
rect 91 657 176 703
rect 32 644 176 657
rect 224 703 336 716
rect 224 657 237 703
rect 283 657 336 703
rect 224 644 336 657
rect 384 703 540 716
rect 384 657 397 703
rect 443 657 540 703
rect 384 644 540 657
rect 120 385 176 644
rect 280 385 336 644
rect 484 584 540 644
rect 120 165 176 209
rect 280 165 336 209
rect 484 165 540 209
<< polycontact >>
rect 45 657 91 703
rect 237 657 283 703
rect 397 657 443 703
<< metal1 >>
rect 0 1359 684 1400
rect 0 1313 69 1359
rect 615 1313 684 1359
rect 0 1178 684 1313
rect 0 1132 409 1178
rect 455 1132 684 1178
rect 45 1075 446 1086
rect 91 1029 446 1075
rect 45 1018 446 1029
rect 42 703 94 972
rect 42 657 45 703
rect 91 657 94 703
rect 42 314 94 657
rect 234 703 286 972
rect 234 657 237 703
rect 283 657 286 703
rect 234 428 286 657
rect 394 703 446 1018
rect 394 657 397 703
rect 443 657 446 703
rect 394 382 446 657
rect 205 371 446 382
rect 251 325 446 371
rect 205 314 446 325
rect 566 1055 618 1086
rect 566 809 569 1055
rect 615 809 618 1055
rect 566 571 618 809
rect 566 325 569 571
rect 615 325 618 571
rect 566 314 618 325
rect 0 222 45 268
rect 91 222 409 268
rect 455 222 684 268
rect 0 87 684 222
rect 0 41 69 87
rect 615 41 684 87
rect 0 0 684 41
<< labels >>
rlabel metal1 s 0 0 684 268 4 vss
port 3 nsew
rlabel metal1 s 0 1132 684 1400 4 vdd
port 5 nsew
rlabel metal1 s 42 314 94 972 4 i0
port 7 nsew
rlabel metal1 s 234 428 286 972 4 i1
port 9 nsew
rlabel metal1 s 566 314 618 1086 4 q
port 11 nsew
<< end >>
