VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO buf_x2
  CLASS BLOCK ;
  FOREIGN buf_x2 ;
  ORIGIN 0.430 0.000 ;
  SIZE 4.280 BY 7.430 ;
  PIN vdd
    ANTENNADIFFAREA 2.639600 ;
    PORT
      LAYER Nwell ;
        RECT -0.430 3.400 3.850 7.430 ;
      LAYER Metal1 ;
        RECT 0.000 5.660 3.420 7.000 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 2.463600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 3.420 1.340 ;
    END
  END vss
  PIN i
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 1.570 0.960 5.430 ;
    END
  END i
  PIN q
    ANTENNADIFFAREA 1.367600 ;
    PORT
      LAYER Metal1 ;
        RECT 2.030 1.570 2.290 5.430 ;
    END
  END q
  OBS
      LAYER Metal1 ;
        RECT 0.210 1.570 0.470 5.430 ;
  END
END buf_x2
END LIBRARY

