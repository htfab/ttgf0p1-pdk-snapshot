magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 460 3782 1094
rect -86 453 86 460
rect 2662 453 3782 460
<< pwell >>
rect 86 453 2662 460
rect -86 -86 3782 453
<< mvnmos >>
rect 388 268 508 340
rect 126 124 246 196
rect 388 124 508 196
rect 820 268 940 340
rect 1188 268 1308 340
rect 820 124 940 196
rect 1188 124 1308 196
rect 1620 267 1740 339
rect 1988 267 2108 339
rect 1620 123 1740 195
rect 1988 123 2108 195
rect 2420 213 2540 285
rect 2420 69 2540 141
rect 2780 69 2900 333
rect 3004 69 3124 333
rect 3228 69 3348 333
rect 3452 69 3572 333
<< mvpmos >>
rect 126 784 226 856
rect 388 784 488 856
rect 388 640 488 712
rect 820 784 920 856
rect 1188 784 1288 856
rect 820 640 920 712
rect 1188 640 1288 712
rect 1620 784 1720 856
rect 1988 784 2088 856
rect 1620 640 1720 712
rect 1988 640 2088 712
rect 2420 784 2520 856
rect 2420 640 2520 712
rect 2780 574 2880 940
rect 3014 574 3114 940
rect 3218 574 3318 940
rect 3452 574 3552 940
<< mvndiff >>
rect 300 327 388 340
rect 300 281 313 327
rect 359 281 388 327
rect 300 268 388 281
rect 508 268 628 340
rect 568 196 628 268
rect 38 183 126 196
rect 38 137 51 183
rect 97 137 126 183
rect 38 124 126 137
rect 246 183 388 196
rect 246 137 275 183
rect 321 137 388 183
rect 246 124 388 137
rect 508 124 628 196
rect 700 268 820 340
rect 940 327 1028 340
rect 940 281 969 327
rect 1015 281 1028 327
rect 940 268 1028 281
rect 1100 327 1188 340
rect 1100 281 1113 327
rect 1159 281 1188 327
rect 1100 268 1188 281
rect 1308 268 1428 340
rect 700 196 760 268
rect 1368 196 1428 268
rect 700 124 820 196
rect 940 183 1188 196
rect 940 137 969 183
rect 1015 137 1188 183
rect 940 124 1188 137
rect 1308 124 1428 196
rect 1500 267 1620 339
rect 1740 326 1828 339
rect 1740 280 1769 326
rect 1815 280 1828 326
rect 1740 267 1828 280
rect 1900 326 1988 339
rect 1900 280 1913 326
rect 1959 280 1988 326
rect 1900 267 1988 280
rect 2108 267 2228 339
rect 1500 195 1560 267
rect 2168 195 2228 267
rect 1500 123 1620 195
rect 1740 182 1988 195
rect 1740 136 1769 182
rect 1815 136 1988 182
rect 1740 123 1988 136
rect 2108 123 2228 195
rect 2300 213 2420 285
rect 2540 272 2628 285
rect 2540 226 2569 272
rect 2615 226 2628 272
rect 2540 213 2628 226
rect 2300 141 2360 213
rect 2700 141 2780 333
rect 2300 69 2420 141
rect 2540 128 2780 141
rect 2540 82 2569 128
rect 2615 82 2780 128
rect 2540 69 2780 82
rect 2900 287 3004 333
rect 2900 147 2929 287
rect 2975 147 3004 287
rect 2900 69 3004 147
rect 3124 277 3228 333
rect 3124 137 3153 277
rect 3199 137 3228 277
rect 3124 69 3228 137
rect 3348 287 3452 333
rect 3348 147 3377 287
rect 3423 147 3452 287
rect 3348 69 3452 147
rect 3572 277 3660 333
rect 3572 137 3601 277
rect 3647 137 3660 277
rect 3572 69 3660 137
<< mvpdiff >>
rect 2700 856 2780 940
rect 38 843 126 856
rect 38 797 51 843
rect 97 797 126 843
rect 38 784 126 797
rect 226 843 388 856
rect 226 797 255 843
rect 301 797 388 843
rect 226 784 388 797
rect 488 784 608 856
rect 548 712 608 784
rect 300 699 388 712
rect 300 653 313 699
rect 359 653 388 699
rect 300 640 388 653
rect 488 640 608 712
rect 700 784 820 856
rect 920 843 1188 856
rect 920 797 949 843
rect 995 797 1188 843
rect 920 784 1188 797
rect 1288 784 1408 856
rect 700 712 760 784
rect 1348 712 1408 784
rect 700 640 820 712
rect 920 699 1008 712
rect 920 653 949 699
rect 995 653 1008 699
rect 920 640 1008 653
rect 1100 699 1188 712
rect 1100 653 1113 699
rect 1159 653 1188 699
rect 1100 640 1188 653
rect 1288 640 1408 712
rect 1500 784 1620 856
rect 1720 843 1988 856
rect 1720 797 1749 843
rect 1795 797 1988 843
rect 1720 784 1988 797
rect 2088 784 2208 856
rect 1500 712 1560 784
rect 2148 712 2208 784
rect 1500 640 1620 712
rect 1720 699 1808 712
rect 1720 653 1749 699
rect 1795 653 1808 699
rect 1720 640 1808 653
rect 1900 699 1988 712
rect 1900 653 1913 699
rect 1959 653 1988 699
rect 1900 640 1988 653
rect 2088 640 2208 712
rect 2300 784 2420 856
rect 2520 843 2780 856
rect 2520 797 2549 843
rect 2595 797 2780 843
rect 2520 784 2780 797
rect 2300 712 2360 784
rect 2300 640 2420 712
rect 2520 699 2608 712
rect 2520 653 2549 699
rect 2595 653 2608 699
rect 2520 640 2608 653
rect 2700 574 2780 784
rect 2880 861 3014 940
rect 2880 721 2939 861
rect 2985 721 3014 861
rect 2880 574 3014 721
rect 3114 927 3218 940
rect 3114 787 3143 927
rect 3189 787 3218 927
rect 3114 574 3218 787
rect 3318 861 3452 940
rect 3318 721 3347 861
rect 3393 721 3452 861
rect 3318 574 3452 721
rect 3552 927 3640 940
rect 3552 787 3581 927
rect 3627 787 3640 927
rect 3552 574 3640 787
<< mvndiffc >>
rect 313 281 359 327
rect 51 137 97 183
rect 275 137 321 183
rect 969 281 1015 327
rect 1113 281 1159 327
rect 969 137 1015 183
rect 1769 280 1815 326
rect 1913 280 1959 326
rect 1769 136 1815 182
rect 2569 226 2615 272
rect 2569 82 2615 128
rect 2929 147 2975 287
rect 3153 137 3199 277
rect 3377 147 3423 287
rect 3601 137 3647 277
<< mvpdiffc >>
rect 51 797 97 843
rect 255 797 301 843
rect 313 653 359 699
rect 949 797 995 843
rect 949 653 995 699
rect 1113 653 1159 699
rect 1749 797 1795 843
rect 1749 653 1795 699
rect 1913 653 1959 699
rect 2549 797 2595 843
rect 2549 653 2595 699
rect 2939 721 2985 861
rect 3143 787 3189 927
rect 3347 721 3393 861
rect 3581 787 3627 927
<< polysilicon >>
rect 2780 940 2880 984
rect 3014 940 3114 984
rect 3218 940 3318 984
rect 3452 940 3552 984
rect 126 856 226 900
rect 388 856 488 900
rect 820 856 920 900
rect 1188 856 1288 900
rect 1620 856 1720 900
rect 1988 856 2088 900
rect 2420 856 2520 900
rect 126 519 226 784
rect 388 712 488 784
rect 820 712 920 784
rect 1188 712 1288 784
rect 1620 712 1720 784
rect 1988 712 2088 784
rect 2420 712 2520 784
rect 126 379 143 519
rect 189 379 226 519
rect 126 240 226 379
rect 388 519 488 640
rect 388 379 401 519
rect 447 384 488 519
rect 820 519 920 640
rect 447 379 508 384
rect 388 340 508 379
rect 820 379 833 519
rect 879 384 920 519
rect 1188 519 1288 640
rect 879 379 940 384
rect 820 340 940 379
rect 1188 379 1201 519
rect 1247 384 1288 519
rect 1620 519 1720 640
rect 1247 379 1308 384
rect 1188 340 1308 379
rect 1620 379 1633 519
rect 1679 383 1720 519
rect 1988 519 2088 640
rect 1679 379 1740 383
rect 126 196 246 240
rect 388 196 508 268
rect 1620 339 1740 379
rect 1988 379 2001 519
rect 2047 383 2088 519
rect 2420 519 2520 640
rect 2047 379 2108 383
rect 1988 339 2108 379
rect 2420 379 2433 519
rect 2479 379 2520 519
rect 820 196 940 268
rect 1188 196 1308 268
rect 2420 329 2520 379
rect 2780 485 2880 574
rect 3014 485 3114 574
rect 3218 485 3318 574
rect 3452 485 3552 574
rect 2780 472 3552 485
rect 2780 426 2793 472
rect 3215 426 3552 472
rect 2780 413 3552 426
rect 2780 333 2900 413
rect 3004 333 3124 413
rect 3228 333 3348 413
rect 3452 377 3552 413
rect 3452 333 3572 377
rect 2420 285 2540 329
rect 1620 195 1740 267
rect 1988 195 2108 267
rect 126 80 246 124
rect 388 80 508 124
rect 820 80 940 124
rect 1188 80 1308 124
rect 2420 141 2540 213
rect 1620 79 1740 123
rect 1988 79 2108 123
rect 2420 25 2540 69
rect 2780 25 2900 69
rect 3004 25 3124 69
rect 3228 25 3348 69
rect 3452 25 3572 69
<< polycontact >>
rect 143 379 189 519
rect 401 379 447 519
rect 833 379 879 519
rect 1201 379 1247 519
rect 1633 379 1679 519
rect 2001 379 2047 519
rect 2433 379 2479 519
rect 2793 426 3215 472
<< metal1 >>
rect 0 927 3696 1098
rect 0 918 3143 927
rect 40 843 97 854
rect 40 797 51 843
rect 40 611 97 797
rect 255 843 301 918
rect 255 786 301 797
rect 949 843 995 918
rect 949 786 995 797
rect 1749 843 1795 918
rect 1749 786 1795 797
rect 2549 843 2595 918
rect 2549 786 2595 797
rect 2939 861 2994 872
rect 2985 721 2994 861
rect 3189 918 3581 927
rect 3143 776 3189 787
rect 3347 861 3393 872
rect 949 699 995 710
rect 302 653 313 699
rect 359 653 550 699
rect 40 607 283 611
rect 40 565 458 607
rect 40 183 86 565
rect 264 561 458 565
rect 390 519 458 561
rect 132 379 143 519
rect 189 379 200 519
rect 390 379 401 519
rect 447 379 458 519
rect 132 354 200 379
rect 504 327 550 653
rect 833 519 879 530
rect 833 327 879 379
rect 302 281 313 327
rect 359 281 879 327
rect 949 425 995 653
rect 1113 699 1159 710
rect 1113 611 1159 653
rect 1749 699 1795 710
rect 1113 565 1350 611
rect 1190 425 1201 519
rect 949 379 1201 425
rect 1247 379 1258 519
rect 949 327 1015 379
rect 1304 327 1350 565
rect 1633 519 1679 530
rect 1633 327 1679 379
rect 949 281 969 327
rect 1102 281 1113 327
rect 1159 281 1679 327
rect 1749 425 1795 653
rect 1913 699 1959 710
rect 1913 611 1959 653
rect 2549 699 2595 710
rect 1913 565 2150 611
rect 1990 425 2001 519
rect 1749 379 2001 425
rect 2047 379 2058 519
rect 2104 414 2150 565
rect 2433 519 2479 530
rect 2104 379 2433 414
rect 1749 326 1815 379
rect 2104 368 2479 379
rect 2549 472 2595 653
rect 2939 624 2994 721
rect 3627 918 3696 927
rect 3581 776 3627 787
rect 3347 624 3393 721
rect 2939 578 3393 624
rect 2549 426 2793 472
rect 3215 426 3226 472
rect 2104 326 2150 368
rect 949 270 1015 281
rect 1749 280 1769 326
rect 1902 280 1913 326
rect 1959 280 2150 326
rect 1749 269 1815 280
rect 2549 272 2615 426
rect 3272 380 3318 578
rect 2549 226 2569 272
rect 2549 215 2615 226
rect 2929 334 3423 380
rect 2929 287 2975 334
rect 275 183 321 194
rect 40 137 51 183
rect 97 137 108 183
rect 275 90 321 137
rect 969 183 1015 194
rect 969 90 1015 137
rect 1769 182 1815 193
rect 1769 90 1815 136
rect 2569 128 2615 139
rect 2929 136 2975 147
rect 3153 277 3199 288
rect 0 82 2569 90
rect 3153 90 3199 137
rect 3377 287 3423 334
rect 3377 136 3423 147
rect 3601 277 3647 288
rect 3601 90 3647 137
rect 2615 82 3696 90
rect 0 -90 3696 82
<< labels >>
flabel metal1 s 132 354 200 519 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 3696 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 3601 194 3647 288 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 3347 624 3393 872 0 FreeSans 200 0 0 0 Z
port 2 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 2939 624 2994 872 1 Z
port 2 nsew default output
rlabel metal1 s 2939 578 3393 624 1 Z
port 2 nsew default output
rlabel metal1 s 3272 380 3318 578 1 Z
port 2 nsew default output
rlabel metal1 s 2929 334 3423 380 1 Z
port 2 nsew default output
rlabel metal1 s 3377 136 3423 334 1 Z
port 2 nsew default output
rlabel metal1 s 2929 136 2975 334 1 Z
port 2 nsew default output
rlabel metal1 s 3581 786 3627 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3143 786 3189 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2549 786 2595 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1749 786 1795 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 949 786 995 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 255 786 301 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3581 776 3627 786 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3143 776 3189 786 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3153 194 3199 288 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3601 193 3647 194 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3153 193 3199 194 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 969 193 1015 194 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 275 193 321 194 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3601 139 3647 193 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3153 139 3199 193 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1769 139 1815 193 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 969 139 1015 193 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 275 139 321 193 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3601 90 3647 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3153 90 3199 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2569 90 2615 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1769 90 1815 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 969 90 1015 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 275 90 321 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3696 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3696 1008
string GDS_END 763338
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 755012
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
