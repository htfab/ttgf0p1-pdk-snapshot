magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 5910 1094
<< pwell >>
rect -86 -86 5910 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 1053 68 1173 332
rect 1277 68 1397 332
rect 1501 68 1621 332
rect 1725 68 1845 332
rect 1949 68 2069 332
rect 2173 68 2293 332
rect 2397 68 2517 332
rect 2621 68 2741 332
rect 2845 68 2965 332
rect 3069 68 3189 332
rect 3293 68 3413 332
rect 3517 68 3637 332
rect 3741 68 3861 332
rect 3965 68 4085 332
rect 4189 68 4309 332
rect 4413 68 4533 332
rect 4637 68 4757 332
rect 4861 68 4981 332
rect 5085 68 5205 332
rect 5309 68 5429 332
rect 5533 68 5653 332
<< mvpmos >>
rect 237 575 337 935
rect 441 575 541 935
rect 645 575 745 935
rect 1033 580 1133 940
rect 1325 580 1425 940
rect 1529 580 1629 940
rect 1821 580 1921 940
rect 2025 580 2125 940
rect 2229 580 2329 940
rect 2433 580 2533 940
rect 2637 580 2737 940
rect 2855 580 2955 940
rect 3079 580 3179 940
rect 3303 580 3403 940
rect 3527 580 3627 940
rect 3751 580 3851 940
rect 3975 580 4075 940
rect 4199 580 4299 940
rect 4403 580 4503 940
rect 4607 580 4707 940
rect 4811 580 4911 940
rect 5015 580 5115 940
rect 5219 580 5319 940
rect 5423 580 5523 940
<< mvndiff >>
rect 36 297 124 333
rect 36 157 49 297
rect 95 157 124 297
rect 36 69 124 157
rect 244 203 348 333
rect 244 157 273 203
rect 319 157 348 203
rect 244 69 348 157
rect 468 297 572 333
rect 468 157 497 297
rect 543 157 572 297
rect 468 69 572 157
rect 692 319 780 333
rect 692 273 721 319
rect 767 273 780 319
rect 692 69 780 273
rect 965 311 1053 332
rect 965 265 978 311
rect 1024 265 1053 311
rect 965 68 1053 265
rect 1173 127 1277 332
rect 1173 81 1202 127
rect 1248 81 1277 127
rect 1173 68 1277 81
rect 1397 311 1501 332
rect 1397 265 1426 311
rect 1472 265 1501 311
rect 1397 68 1501 265
rect 1621 127 1725 332
rect 1621 81 1650 127
rect 1696 81 1725 127
rect 1621 68 1725 81
rect 1845 209 1949 332
rect 1845 163 1874 209
rect 1920 163 1949 209
rect 1845 68 1949 163
rect 2069 297 2173 332
rect 2069 157 2098 297
rect 2144 157 2173 297
rect 2069 68 2173 157
rect 2293 319 2397 332
rect 2293 179 2322 319
rect 2368 179 2397 319
rect 2293 68 2397 179
rect 2517 297 2621 332
rect 2517 157 2546 297
rect 2592 157 2621 297
rect 2517 68 2621 157
rect 2741 319 2845 332
rect 2741 179 2770 319
rect 2816 179 2845 319
rect 2741 68 2845 179
rect 2965 297 3069 332
rect 2965 157 2994 297
rect 3040 157 3069 297
rect 2965 68 3069 157
rect 3189 274 3293 332
rect 3189 228 3218 274
rect 3264 228 3293 274
rect 3189 68 3293 228
rect 3413 127 3517 332
rect 3413 81 3442 127
rect 3488 81 3517 127
rect 3413 68 3517 81
rect 3637 319 3741 332
rect 3637 179 3666 319
rect 3712 179 3741 319
rect 3637 68 3741 179
rect 3861 127 3965 332
rect 3861 81 3890 127
rect 3936 81 3965 127
rect 3861 68 3965 81
rect 4085 319 4189 332
rect 4085 179 4114 319
rect 4160 179 4189 319
rect 4085 68 4189 179
rect 4309 127 4413 332
rect 4309 81 4338 127
rect 4384 81 4413 127
rect 4309 68 4413 81
rect 4533 319 4637 332
rect 4533 179 4562 319
rect 4608 179 4637 319
rect 4533 68 4637 179
rect 4757 127 4861 332
rect 4757 81 4786 127
rect 4832 81 4861 127
rect 4757 68 4861 81
rect 4981 319 5085 332
rect 4981 179 5010 319
rect 5056 179 5085 319
rect 4981 68 5085 179
rect 5205 127 5309 332
rect 5205 81 5234 127
rect 5280 81 5309 127
rect 5205 68 5309 81
rect 5429 280 5533 332
rect 5429 234 5458 280
rect 5504 234 5533 280
rect 5429 68 5533 234
rect 5653 297 5741 332
rect 5653 157 5682 297
rect 5728 157 5741 297
rect 5653 68 5741 157
<< mvpdiff >>
rect 1193 959 1265 972
rect 1193 940 1206 959
rect 149 845 237 935
rect 149 705 162 845
rect 208 705 237 845
rect 149 575 237 705
rect 337 845 441 935
rect 337 705 366 845
rect 412 705 441 845
rect 337 575 441 705
rect 541 845 645 935
rect 541 705 570 845
rect 616 705 645 845
rect 541 575 645 705
rect 745 753 833 935
rect 745 613 774 753
rect 820 613 833 753
rect 745 575 833 613
rect 945 753 1033 940
rect 945 613 958 753
rect 1004 613 1033 753
rect 945 580 1033 613
rect 1133 913 1206 940
rect 1252 940 1265 959
rect 1689 959 1761 972
rect 1689 940 1702 959
rect 1252 913 1325 940
rect 1133 580 1325 913
rect 1425 753 1529 940
rect 1425 613 1454 753
rect 1500 613 1529 753
rect 1425 580 1529 613
rect 1629 913 1702 940
rect 1748 940 1761 959
rect 1748 913 1821 940
rect 1629 580 1821 913
rect 1921 752 2025 940
rect 1921 612 1950 752
rect 1996 612 2025 752
rect 1921 580 2025 612
rect 2125 847 2229 940
rect 2125 801 2154 847
rect 2200 801 2229 847
rect 2125 580 2229 801
rect 2329 845 2433 940
rect 2329 705 2358 845
rect 2404 705 2433 845
rect 2329 580 2433 705
rect 2533 845 2637 940
rect 2533 705 2562 845
rect 2608 705 2637 845
rect 2533 580 2637 705
rect 2737 845 2855 940
rect 2737 705 2766 845
rect 2812 705 2855 845
rect 2737 580 2855 705
rect 2955 927 3079 940
rect 2955 787 2984 927
rect 3030 787 3079 927
rect 2955 580 3079 787
rect 3179 845 3303 940
rect 3179 705 3228 845
rect 3274 705 3303 845
rect 3179 580 3303 705
rect 3403 849 3527 940
rect 3403 803 3432 849
rect 3478 803 3527 849
rect 3403 580 3527 803
rect 3627 845 3751 940
rect 3627 705 3656 845
rect 3702 705 3751 845
rect 3627 580 3751 705
rect 3851 845 3975 940
rect 3851 799 3880 845
rect 3926 799 3975 845
rect 3851 580 3975 799
rect 4075 845 4199 940
rect 4075 705 4104 845
rect 4150 705 4199 845
rect 4075 580 4199 705
rect 4299 845 4403 940
rect 4299 799 4328 845
rect 4374 799 4403 845
rect 4299 580 4403 799
rect 4503 845 4607 940
rect 4503 705 4532 845
rect 4578 705 4607 845
rect 4503 580 4607 705
rect 4707 845 4811 940
rect 4707 799 4736 845
rect 4782 799 4811 845
rect 4707 580 4811 799
rect 4911 845 5015 940
rect 4911 705 4940 845
rect 4986 705 5015 845
rect 4911 580 5015 705
rect 5115 845 5219 940
rect 5115 799 5144 845
rect 5190 799 5219 845
rect 5115 580 5219 799
rect 5319 845 5423 940
rect 5319 705 5348 845
rect 5394 705 5423 845
rect 5319 580 5423 705
rect 5523 845 5611 940
rect 5523 799 5552 845
rect 5598 799 5611 845
rect 5523 580 5611 799
<< mvndiffc >>
rect 49 157 95 297
rect 273 157 319 203
rect 497 157 543 297
rect 721 273 767 319
rect 978 265 1024 311
rect 1202 81 1248 127
rect 1426 265 1472 311
rect 1650 81 1696 127
rect 1874 163 1920 209
rect 2098 157 2144 297
rect 2322 179 2368 319
rect 2546 157 2592 297
rect 2770 179 2816 319
rect 2994 157 3040 297
rect 3218 228 3264 274
rect 3442 81 3488 127
rect 3666 179 3712 319
rect 3890 81 3936 127
rect 4114 179 4160 319
rect 4338 81 4384 127
rect 4562 179 4608 319
rect 4786 81 4832 127
rect 5010 179 5056 319
rect 5234 81 5280 127
rect 5458 234 5504 280
rect 5682 157 5728 297
<< mvpdiffc >>
rect 162 705 208 845
rect 366 705 412 845
rect 570 705 616 845
rect 774 613 820 753
rect 958 613 1004 753
rect 1206 913 1252 959
rect 1454 613 1500 753
rect 1702 913 1748 959
rect 1950 612 1996 752
rect 2154 801 2200 847
rect 2358 705 2404 845
rect 2562 705 2608 845
rect 2766 705 2812 845
rect 2984 787 3030 927
rect 3228 705 3274 845
rect 3432 803 3478 849
rect 3656 705 3702 845
rect 3880 799 3926 845
rect 4104 705 4150 845
rect 4328 799 4374 845
rect 4532 705 4578 845
rect 4736 799 4782 845
rect 4940 705 4986 845
rect 5144 799 5190 845
rect 5348 705 5394 845
rect 5552 799 5598 845
<< polysilicon >>
rect 237 935 337 979
rect 441 935 541 979
rect 645 935 745 979
rect 1033 940 1133 984
rect 1325 940 1425 984
rect 1529 940 1629 984
rect 1821 940 1921 984
rect 2025 940 2125 984
rect 2229 940 2329 984
rect 2433 940 2533 984
rect 2637 940 2737 984
rect 2855 940 2955 984
rect 3079 940 3179 984
rect 3303 940 3403 984
rect 3527 940 3627 984
rect 3751 940 3851 984
rect 3975 940 4075 984
rect 4199 940 4299 984
rect 4403 940 4503 984
rect 4607 940 4707 984
rect 4811 940 4911 984
rect 5015 940 5115 984
rect 5219 940 5319 984
rect 5423 940 5523 984
rect 237 515 337 575
rect 441 515 541 575
rect 124 504 541 515
rect 645 542 745 575
rect 124 475 553 504
rect 645 496 658 542
rect 704 496 745 542
rect 1033 536 1133 580
rect 645 483 745 496
rect 124 414 244 475
rect 513 448 553 475
rect 1053 464 1133 536
rect 1325 464 1425 580
rect 1529 536 1629 580
rect 1529 464 1621 536
rect 1821 518 1921 580
rect 124 368 148 414
rect 194 368 244 414
rect 124 333 244 368
rect 348 414 420 427
rect 348 368 361 414
rect 407 377 420 414
rect 513 408 612 448
rect 572 377 612 408
rect 1053 414 1621 464
rect 407 368 468 377
rect 348 333 468 368
rect 572 333 692 377
rect 1053 368 1114 414
rect 1160 392 1621 414
rect 1160 368 1173 392
rect 1053 332 1173 368
rect 1277 332 1397 392
rect 1501 332 1621 392
rect 1725 505 1921 518
rect 1725 365 1738 505
rect 1784 464 1921 505
rect 2025 464 2125 580
rect 2229 464 2329 580
rect 2433 464 2533 580
rect 2637 464 2737 580
rect 2855 464 2955 580
rect 3079 547 3179 580
rect 3079 501 3105 547
rect 3151 520 3179 547
rect 3303 547 3403 580
rect 3303 520 3330 547
rect 3151 501 3330 520
rect 3376 520 3403 547
rect 3527 547 3627 580
rect 3527 520 3556 547
rect 3376 501 3556 520
rect 3602 520 3627 547
rect 3751 547 3851 580
rect 3751 520 3778 547
rect 3602 501 3778 520
rect 3824 520 3851 547
rect 3975 547 4075 580
rect 3975 520 4002 547
rect 3824 501 4002 520
rect 4048 520 4075 547
rect 4199 547 4299 580
rect 4199 520 4228 547
rect 4048 501 4228 520
rect 4274 520 4299 547
rect 4403 547 4503 580
rect 4403 520 4431 547
rect 4274 501 4431 520
rect 4477 520 4503 547
rect 4607 547 4707 580
rect 4607 520 4631 547
rect 4477 501 4631 520
rect 4677 520 4707 547
rect 4811 547 4911 580
rect 4811 520 4838 547
rect 4677 501 4838 520
rect 4884 520 4911 547
rect 5015 547 5115 580
rect 5015 520 5044 547
rect 4884 501 5044 520
rect 5090 520 5115 547
rect 5219 520 5319 580
rect 5423 520 5523 580
rect 5090 501 5523 520
rect 3079 480 5523 501
rect 1784 392 2955 464
rect 1784 365 1845 392
rect 1725 332 1845 365
rect 1949 332 2069 392
rect 2173 332 2293 392
rect 2397 332 2517 392
rect 2621 332 2741 392
rect 2845 376 2955 392
rect 3069 411 5653 432
rect 2845 332 2965 376
rect 3069 365 3101 411
rect 3147 392 3330 411
rect 3147 365 3189 392
rect 3069 332 3189 365
rect 3293 365 3330 392
rect 3376 392 3558 411
rect 3376 365 3413 392
rect 3293 332 3413 365
rect 3517 365 3558 392
rect 3604 392 3777 411
rect 3604 365 3637 392
rect 3517 332 3637 365
rect 3741 365 3777 392
rect 3823 392 4000 411
rect 3823 365 3861 392
rect 3741 332 3861 365
rect 3965 365 4000 392
rect 4046 392 4225 411
rect 4046 365 4085 392
rect 3965 332 4085 365
rect 4189 365 4225 392
rect 4271 392 4447 411
rect 4271 365 4309 392
rect 4189 332 4309 365
rect 4413 365 4447 392
rect 4493 392 4674 411
rect 4493 365 4533 392
rect 4413 332 4533 365
rect 4637 365 4674 392
rect 4720 392 4899 411
rect 4720 365 4757 392
rect 4637 332 4757 365
rect 4861 365 4899 392
rect 4945 392 5122 411
rect 4945 365 4981 392
rect 4861 332 4981 365
rect 5085 365 5122 392
rect 5168 392 5653 411
rect 5168 365 5205 392
rect 5085 332 5205 365
rect 5309 332 5429 392
rect 5533 332 5653 392
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 1053 24 1173 68
rect 1277 24 1397 68
rect 1501 24 1621 68
rect 1725 24 1845 68
rect 1949 24 2069 68
rect 2173 24 2293 68
rect 2397 24 2517 68
rect 2621 24 2741 68
rect 2845 24 2965 68
rect 3069 24 3189 68
rect 3293 24 3413 68
rect 3517 24 3637 68
rect 3741 24 3861 68
rect 3965 24 4085 68
rect 4189 24 4309 68
rect 4413 24 4533 68
rect 4637 24 4757 68
rect 4861 24 4981 68
rect 5085 24 5205 68
rect 5309 24 5429 68
rect 5533 24 5653 68
<< polycontact >>
rect 658 496 704 542
rect 148 368 194 414
rect 361 368 407 414
rect 1114 368 1160 414
rect 1738 365 1784 505
rect 3105 501 3151 547
rect 3330 501 3376 547
rect 3556 501 3602 547
rect 3778 501 3824 547
rect 4002 501 4048 547
rect 4228 501 4274 547
rect 4431 501 4477 547
rect 4631 501 4677 547
rect 4838 501 4884 547
rect 5044 501 5090 547
rect 3101 365 3147 411
rect 3330 365 3376 411
rect 3558 365 3604 411
rect 3777 365 3823 411
rect 4000 365 4046 411
rect 4225 365 4271 411
rect 4447 365 4493 411
rect 4674 365 4720 411
rect 4899 365 4945 411
rect 5122 365 5168 411
<< metal1 >>
rect 0 959 5824 1098
rect 0 918 1206 959
rect 162 845 208 856
rect 162 634 208 705
rect 366 845 412 918
rect 1252 918 1702 959
rect 1206 902 1252 913
rect 1748 927 5824 959
rect 1748 918 2984 927
rect 1702 902 1748 913
rect 366 694 412 705
rect 570 845 1996 856
rect 616 810 1996 845
rect 570 694 616 705
rect 774 753 820 764
rect 162 588 715 634
rect 361 542 715 588
rect 142 414 194 542
rect 142 368 148 414
rect 142 354 194 368
rect 361 496 658 542
rect 704 496 715 542
rect 361 414 407 496
rect 774 411 820 613
rect 361 308 407 368
rect 618 365 820 411
rect 49 297 407 308
rect 95 262 407 297
rect 497 297 543 308
rect 49 146 95 157
rect 273 203 319 214
rect 273 90 319 157
rect 618 219 664 365
rect 866 319 912 810
rect 958 753 1500 764
rect 1004 718 1454 753
rect 958 602 1004 613
rect 1114 414 1202 654
rect 1454 505 1500 613
rect 1950 752 1996 810
rect 2154 847 2200 918
rect 2154 790 2200 801
rect 2358 845 2404 856
rect 1950 547 1996 612
rect 2358 547 2404 705
rect 2562 845 2608 918
rect 2562 694 2608 705
rect 2766 845 2812 856
rect 3030 918 5824 927
rect 2984 776 3030 787
rect 3228 845 3274 856
rect 2766 547 2812 705
rect 3432 849 3478 918
rect 3432 792 3478 803
rect 3656 845 3702 856
rect 3228 698 3274 705
rect 3880 845 3926 918
rect 3880 788 3926 799
rect 4104 845 4150 856
rect 3656 698 3702 705
rect 4328 845 4374 918
rect 4328 788 4374 799
rect 4532 845 4578 856
rect 4104 698 4150 705
rect 4736 845 4782 918
rect 4736 788 4782 799
rect 4940 845 4986 856
rect 4532 698 4578 705
rect 5144 845 5190 918
rect 5144 788 5190 799
rect 5347 845 5394 856
rect 4940 698 4986 705
rect 5347 705 5348 845
rect 5347 698 5394 705
rect 3228 602 5394 698
rect 5552 845 5598 918
rect 5552 694 5598 799
rect 1454 446 1738 505
rect 1160 368 1202 414
rect 1114 357 1202 368
rect 1784 365 1795 505
rect 1950 501 3105 547
rect 3151 501 3330 547
rect 3376 501 3556 547
rect 3602 501 3778 547
rect 3824 501 4002 547
rect 4048 501 4228 547
rect 4274 501 4431 547
rect 4477 501 4631 547
rect 4677 501 4838 547
rect 4884 501 5044 547
rect 5090 501 5114 547
rect 710 273 721 319
rect 767 273 912 319
rect 1738 311 1795 365
rect 967 265 978 311
rect 1024 265 1426 311
rect 1472 265 1795 311
rect 1886 365 3101 411
rect 3147 365 3330 411
rect 3376 365 3558 411
rect 3604 365 3777 411
rect 3823 365 4000 411
rect 4046 365 4225 411
rect 4271 365 4447 411
rect 4493 365 4674 411
rect 4720 365 4899 411
rect 4945 365 5122 411
rect 5168 365 5188 411
rect 1886 219 1932 365
rect 2322 319 2368 365
rect 543 209 1932 219
rect 543 173 1874 209
rect 1863 163 1874 173
rect 1920 163 1932 209
rect 2098 297 2144 308
rect 497 146 543 157
rect 2770 319 2816 365
rect 5290 319 5396 602
rect 2322 168 2368 179
rect 2546 297 2592 308
rect 1191 90 1202 127
rect 0 81 1202 90
rect 1248 90 1259 127
rect 1639 90 1650 127
rect 1248 81 1650 90
rect 1696 90 1707 127
rect 2098 90 2144 157
rect 2770 168 2816 179
rect 2994 297 3040 308
rect 2546 90 2592 157
rect 3218 274 3666 319
rect 3264 228 3666 274
rect 3218 179 3666 228
rect 3712 179 4114 319
rect 4160 179 4562 319
rect 4608 179 5010 319
rect 5056 280 5504 319
rect 5056 234 5458 280
rect 5056 179 5504 234
rect 5682 297 5728 308
rect 2994 90 3040 157
rect 3431 90 3442 127
rect 1696 81 3442 90
rect 3488 90 3499 127
rect 3879 90 3890 127
rect 3488 81 3890 90
rect 3936 90 3947 127
rect 4327 90 4338 127
rect 3936 81 4338 90
rect 4384 90 4395 127
rect 4775 90 4786 127
rect 4384 81 4786 90
rect 4832 90 4843 127
rect 5223 90 5234 127
rect 4832 81 5234 90
rect 5280 90 5291 127
rect 5682 90 5728 157
rect 5280 81 5824 90
rect 0 -90 5824 81
<< labels >>
flabel metal1 s 142 354 194 542 0 FreeSans 200 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1114 357 1202 654 0 FreeSans 200 0 0 0 I
port 2 nsew default input
flabel metal1 s 0 918 5824 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 5682 214 5728 308 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 5347 698 5394 856 0 FreeSans 200 0 0 0 ZN
port 3 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 4940 698 4986 856 1 ZN
port 3 nsew default output
rlabel metal1 s 4532 698 4578 856 1 ZN
port 3 nsew default output
rlabel metal1 s 4104 698 4150 856 1 ZN
port 3 nsew default output
rlabel metal1 s 3656 698 3702 856 1 ZN
port 3 nsew default output
rlabel metal1 s 3228 698 3274 856 1 ZN
port 3 nsew default output
rlabel metal1 s 3228 602 5394 698 1 ZN
port 3 nsew default output
rlabel metal1 s 5290 319 5396 602 1 ZN
port 3 nsew default output
rlabel metal1 s 3218 179 5504 319 1 ZN
port 3 nsew default output
rlabel metal1 s 5552 902 5598 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5144 902 5190 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4736 902 4782 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4328 902 4374 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3880 902 3926 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3432 902 3478 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2984 902 3030 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2562 902 2608 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2154 902 2200 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1702 902 1748 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1206 902 1252 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 366 902 412 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5552 792 5598 902 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5144 792 5190 902 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4736 792 4782 902 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4328 792 4374 902 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3880 792 3926 902 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3432 792 3478 902 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2984 792 3030 902 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2562 792 2608 902 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2154 792 2200 902 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 366 792 412 902 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5552 790 5598 792 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5144 790 5190 792 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4736 790 4782 792 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4328 790 4374 792 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3880 790 3926 792 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2984 790 3030 792 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2562 790 2608 792 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2154 790 2200 792 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 366 790 412 792 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5552 788 5598 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5144 788 5190 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4736 788 4782 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4328 788 4374 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3880 788 3926 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2984 788 3030 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2562 788 2608 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 366 788 412 790 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5552 776 5598 788 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2984 776 3030 788 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2562 776 2608 788 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 366 776 412 788 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5552 694 5598 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2562 694 2608 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 366 694 412 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2994 214 3040 308 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2546 214 2592 308 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2098 214 2144 308 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5682 127 5728 214 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2994 127 3040 214 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2546 127 2592 214 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2098 127 2144 214 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 127 319 214 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5682 90 5728 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5223 90 5291 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4775 90 4843 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4327 90 4395 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3879 90 3947 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3431 90 3499 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2994 90 3040 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2546 90 2592 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2098 90 2144 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1639 90 1707 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1191 90 1259 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 5824 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5824 1008
string GDS_END 965970
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 953662
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
