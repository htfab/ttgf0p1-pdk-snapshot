magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 998 1486
<< nmos >>
rect 120 209 176 385
rect 280 209 336 385
rect 440 209 496 385
rect 600 209 656 385
<< pmos >>
rect 120 1015 176 1191
rect 280 1015 336 1191
rect 440 1015 496 1191
rect 600 1015 656 1191
<< ndiff >>
rect 32 371 120 385
rect 32 325 45 371
rect 91 325 120 371
rect 32 209 120 325
rect 176 209 280 385
rect 336 268 440 385
rect 336 222 365 268
rect 411 222 440 268
rect 336 209 440 222
rect 496 209 600 385
rect 656 371 744 385
rect 656 325 685 371
rect 731 325 744 371
rect 656 209 744 325
<< pdiff >>
rect 32 1178 120 1191
rect 32 1132 45 1178
rect 91 1132 120 1178
rect 32 1015 120 1132
rect 176 1075 280 1191
rect 176 1029 205 1075
rect 251 1029 280 1075
rect 176 1015 280 1029
rect 336 1178 440 1191
rect 336 1132 365 1178
rect 411 1132 440 1178
rect 336 1015 440 1132
rect 496 1075 600 1191
rect 496 1029 525 1075
rect 571 1029 600 1075
rect 496 1015 600 1029
rect 656 1178 744 1191
rect 656 1132 685 1178
rect 731 1132 744 1178
rect 656 1015 744 1132
<< ndiffc >>
rect 45 325 91 371
rect 365 222 411 268
rect 685 325 731 371
<< pdiffc >>
rect 45 1132 91 1178
rect 205 1029 251 1075
rect 365 1132 411 1178
rect 525 1029 571 1075
rect 685 1132 731 1178
<< psubdiff >>
rect 28 87 884 100
rect 28 41 83 87
rect 829 41 884 87
rect 28 28 884 41
<< nsubdiff >>
rect 28 1359 884 1372
rect 28 1313 83 1359
rect 829 1313 884 1359
rect 28 1300 884 1313
<< psubdiffcont >>
rect 83 41 829 87
<< nsubdiffcont >>
rect 83 1313 829 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 600 1191 656 1235
rect 120 782 176 1015
rect 32 769 176 782
rect 32 723 45 769
rect 91 723 176 769
rect 32 710 176 723
rect 120 385 176 710
rect 280 650 336 1015
rect 440 782 496 1015
rect 384 769 496 782
rect 384 723 397 769
rect 443 723 496 769
rect 384 710 496 723
rect 228 637 336 650
rect 228 591 241 637
rect 287 591 336 637
rect 228 578 336 591
rect 280 385 336 578
rect 440 385 496 710
rect 600 650 656 1015
rect 600 637 682 650
rect 600 591 623 637
rect 669 591 682 637
rect 600 578 682 591
rect 600 385 656 578
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
rect 600 165 656 209
<< polycontact >>
rect 45 723 91 769
rect 397 723 443 769
rect 241 591 287 637
rect 623 591 669 637
<< metal1 >>
rect 0 1359 912 1400
rect 0 1313 83 1359
rect 829 1313 912 1359
rect 0 1178 912 1313
rect 0 1132 45 1178
rect 91 1132 365 1178
rect 411 1132 685 1178
rect 731 1132 912 1178
rect 42 769 94 1086
rect 42 723 45 769
rect 91 723 94 769
rect 42 428 94 723
rect 140 1075 251 1086
rect 140 1029 205 1075
rect 140 1018 251 1029
rect 522 1075 574 1086
rect 522 1029 525 1075
rect 571 1029 574 1075
rect 140 780 192 1018
rect 140 769 443 780
rect 140 723 397 769
rect 140 712 443 723
rect 140 382 192 712
rect 522 648 574 1029
rect 241 637 574 648
rect 287 591 574 637
rect 241 580 574 591
rect 45 371 192 382
rect 91 325 192 371
rect 45 314 192 325
rect 522 382 574 580
rect 620 637 672 1086
rect 620 591 623 637
rect 669 591 672 637
rect 620 428 672 591
rect 522 371 731 382
rect 522 325 685 371
rect 522 314 731 325
rect 0 222 365 268
rect 411 222 912 268
rect 0 87 912 222
rect 0 41 83 87
rect 829 41 912 87
rect 0 0 912 41
<< labels >>
rlabel metal1 s 140 314 192 1086 4 q
port 3 nsew
rlabel metal1 s 0 1132 912 1400 4 vdd
port 5 nsew
rlabel metal1 s 0 0 912 268 4 vss
port 7 nsew
rlabel metal1 s 42 428 94 1086 4 nset
port 9 nsew
rlabel metal1 s 522 314 574 1086 4 nq
port 11 nsew
rlabel metal1 s 620 428 672 1086 4 nrst
port 13 nsew
<< end >>
