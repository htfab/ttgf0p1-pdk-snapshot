magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 758 1094
<< pwell >>
rect -86 -86 758 453
<< metal1 >>
rect 0 918 672 1098
rect 49 710 95 918
rect 273 766 319 872
rect 273 710 420 766
rect 477 710 523 918
rect 366 578 420 710
rect 72 454 328 542
rect 374 408 420 578
rect 273 362 420 408
rect 49 90 95 257
rect 273 189 319 362
rect 497 90 543 257
rect 0 -90 672 90
<< labels >>
rlabel metal1 s 72 454 328 542 6 I
port 1 nsew default input
rlabel metal1 s 273 189 319 362 6 ZN
port 2 nsew default output
rlabel metal1 s 273 362 420 408 6 ZN
port 2 nsew default output
rlabel metal1 s 374 408 420 578 6 ZN
port 2 nsew default output
rlabel metal1 s 366 578 420 710 6 ZN
port 2 nsew default output
rlabel metal1 s 273 710 420 766 6 ZN
port 2 nsew default output
rlabel metal1 s 273 766 319 872 6 ZN
port 2 nsew default output
rlabel metal1 s 477 710 523 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 918 672 1098 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 453 758 1094 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 758 453 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -90 672 90 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 257 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 257 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 672 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1446214
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1443520
<< end >>
