VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO and3_x1
  CLASS BLOCK ;
  FOREIGN and3_x1 ;
  ORIGIN 0.430 0.000 ;
  SIZE 5.420 BY 7.430 ;
  PIN vdd
    ANTENNADIFFAREA 3.175400 ;
    PORT
      LAYER Nwell ;
        RECT -0.430 3.400 4.990 7.430 ;
      LAYER Metal1 ;
        RECT 0.000 5.660 4.560 7.000 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 2.629800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 4.560 1.340 ;
    END
  END vss
  PIN i0
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.210 2.140 0.470 4.860 ;
    END
  END i0
  PIN i1
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.170 2.140 1.430 4.860 ;
    END
  END i1
  PIN i2
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.970 2.140 2.230 4.860 ;
    END
  END i2
  PIN q
    ANTENNADIFFAREA 1.738000 ;
    PORT
      LAYER Metal1 ;
        RECT 3.630 1.570 3.890 5.430 ;
    END
  END q
  OBS
      LAYER Metal1 ;
        RECT 0.225 5.090 3.030 5.430 ;
        RECT 2.770 1.910 3.030 5.090 ;
        RECT 0.225 1.570 3.030 1.910 ;
  END
END and3_x1
END LIBRARY

