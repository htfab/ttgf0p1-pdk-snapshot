magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 1990 1094
<< pwell >>
rect -86 -86 1990 453
<< mvnmos >>
rect 135 69 255 333
rect 359 69 479 333
rect 583 69 703 333
rect 951 68 1071 332
rect 1175 68 1295 332
rect 1399 68 1519 332
rect 1623 68 1743 332
<< mvpmos >>
rect 145 573 245 933
rect 349 573 449 933
rect 655 573 755 933
rect 1021 580 1121 940
rect 1225 580 1325 940
rect 1429 580 1529 940
rect 1633 580 1733 940
<< mvndiff >>
rect 47 287 135 333
rect 47 147 60 287
rect 106 147 135 287
rect 47 69 135 147
rect 255 193 359 333
rect 255 147 284 193
rect 330 147 359 193
rect 255 69 359 147
rect 479 287 583 333
rect 479 147 508 287
rect 554 147 583 287
rect 479 69 583 147
rect 703 320 791 333
rect 703 274 732 320
rect 778 274 791 320
rect 703 69 791 274
rect 863 217 951 332
rect 863 171 876 217
rect 922 171 951 217
rect 863 68 951 171
rect 1071 193 1175 332
rect 1071 147 1100 193
rect 1146 147 1175 193
rect 1071 68 1175 147
rect 1295 287 1399 332
rect 1295 147 1324 287
rect 1370 147 1399 287
rect 1295 68 1399 147
rect 1519 287 1623 332
rect 1519 147 1548 287
rect 1594 147 1623 287
rect 1519 68 1623 147
rect 1743 287 1831 332
rect 1743 147 1772 287
rect 1818 147 1831 287
rect 1743 68 1831 147
<< mvpdiff >>
rect 57 831 145 933
rect 57 691 70 831
rect 116 691 145 831
rect 57 573 145 691
rect 245 831 349 933
rect 245 691 274 831
rect 320 691 349 831
rect 245 573 349 691
rect 449 831 655 933
rect 449 691 580 831
rect 626 691 655 831
rect 449 573 655 691
rect 755 769 843 933
rect 755 629 784 769
rect 830 629 843 769
rect 755 573 843 629
rect 933 831 1021 940
rect 933 691 946 831
rect 992 691 1021 831
rect 933 580 1021 691
rect 1121 927 1225 940
rect 1121 881 1150 927
rect 1196 881 1225 927
rect 1121 580 1225 881
rect 1325 739 1429 940
rect 1325 599 1354 739
rect 1400 599 1429 739
rect 1325 580 1429 599
rect 1529 831 1633 940
rect 1529 691 1558 831
rect 1604 691 1633 831
rect 1529 580 1633 691
rect 1733 831 1821 940
rect 1733 691 1762 831
rect 1808 691 1821 831
rect 1733 580 1821 691
<< mvndiffc >>
rect 60 147 106 287
rect 284 147 330 193
rect 508 147 554 287
rect 732 274 778 320
rect 876 171 922 217
rect 1100 147 1146 193
rect 1324 147 1370 287
rect 1548 147 1594 287
rect 1772 147 1818 287
<< mvpdiffc >>
rect 70 691 116 831
rect 274 691 320 831
rect 580 691 626 831
rect 784 629 830 769
rect 946 691 992 831
rect 1150 881 1196 927
rect 1354 599 1400 739
rect 1558 691 1604 831
rect 1762 691 1808 831
<< polysilicon >>
rect 145 933 245 977
rect 349 933 449 977
rect 655 933 755 977
rect 1021 940 1121 984
rect 1225 940 1325 984
rect 1429 940 1529 984
rect 1633 940 1733 984
rect 145 513 245 573
rect 349 513 449 573
rect 655 540 755 573
rect 145 473 607 513
rect 655 494 668 540
rect 714 494 755 540
rect 655 481 755 494
rect 1021 547 1121 580
rect 1021 501 1048 547
rect 1094 501 1121 547
rect 1021 488 1121 501
rect 1225 539 1325 580
rect 1225 493 1238 539
rect 1284 520 1325 539
rect 1429 520 1529 580
rect 1284 493 1529 520
rect 145 425 255 473
rect 567 431 607 473
rect 135 412 255 425
rect 135 366 148 412
rect 194 366 255 412
rect 135 333 255 366
rect 359 412 479 425
rect 359 366 372 412
rect 418 366 479 412
rect 567 394 703 431
rect 359 333 479 366
rect 583 333 703 394
rect 1021 376 1071 488
rect 1225 480 1529 493
rect 951 332 1071 376
rect 1175 411 1519 432
rect 1175 365 1232 411
rect 1278 392 1519 411
rect 1278 365 1295 392
rect 1175 332 1295 365
rect 1399 332 1519 392
rect 1633 411 1733 580
rect 1633 376 1646 411
rect 1623 365 1646 376
rect 1692 376 1733 411
rect 1692 365 1743 376
rect 1623 332 1743 365
rect 135 25 255 69
rect 359 25 479 69
rect 583 25 703 69
rect 951 24 1071 68
rect 1175 24 1295 68
rect 1399 24 1519 68
rect 1623 24 1743 68
<< polycontact >>
rect 668 494 714 540
rect 1048 501 1094 547
rect 1238 493 1284 539
rect 148 366 194 412
rect 372 366 418 412
rect 1232 365 1278 411
rect 1646 365 1692 411
<< metal1 >>
rect 0 927 1904 1098
rect 0 918 1150 927
rect 70 831 116 842
rect 70 634 116 691
rect 274 831 320 918
rect 1196 918 1904 927
rect 274 680 320 691
rect 580 831 992 872
rect 1150 870 1196 881
rect 626 826 946 831
rect 580 680 626 691
rect 784 769 830 780
rect 70 588 725 634
rect 142 412 194 542
rect 142 366 148 412
rect 142 354 194 366
rect 372 540 725 588
rect 372 494 668 540
rect 714 494 725 540
rect 372 412 418 494
rect 784 448 830 629
rect 372 298 418 366
rect 640 402 830 448
rect 917 691 946 826
rect 917 444 992 691
rect 1233 796 1512 842
rect 1233 631 1279 796
rect 1048 585 1279 631
rect 1354 739 1400 750
rect 1048 547 1094 585
rect 1354 542 1400 599
rect 1466 634 1512 796
rect 1558 831 1604 918
rect 1558 680 1604 691
rect 1762 831 1818 842
rect 1808 691 1818 831
rect 1762 634 1818 691
rect 1466 588 1818 634
rect 1048 490 1094 501
rect 1140 493 1238 539
rect 1284 493 1295 539
rect 1140 444 1186 493
rect 640 298 686 402
rect 917 398 1186 444
rect 1232 411 1278 422
rect 917 356 963 398
rect 60 287 418 298
rect 106 252 418 287
rect 508 287 686 298
rect 60 136 106 147
rect 284 193 330 204
rect 284 90 330 147
rect 554 217 686 287
rect 732 320 963 356
rect 778 310 963 320
rect 1232 296 1278 365
rect 1354 298 1426 542
rect 1598 411 1692 542
rect 1598 365 1646 411
rect 1598 354 1692 365
rect 732 263 778 274
rect 1007 250 1278 296
rect 1324 287 1426 298
rect 1007 217 1053 250
rect 554 171 876 217
rect 922 171 1053 217
rect 554 147 1053 171
rect 508 136 1053 147
rect 1100 193 1146 204
rect 1100 90 1146 147
rect 1370 242 1426 287
rect 1548 287 1594 298
rect 1324 136 1370 147
rect 1548 90 1594 147
rect 1772 287 1818 588
rect 1772 136 1818 147
rect 0 -90 1904 90
<< labels >>
flabel metal1 s 142 354 194 542 0 FreeSans 200 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1598 354 1692 542 0 FreeSans 200 0 0 0 I
port 2 nsew default input
flabel metal1 s 0 918 1904 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 1548 204 1594 298 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 1354 542 1400 750 0 FreeSans 200 0 0 0 ZN
port 3 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 1354 298 1426 542 1 ZN
port 3 nsew default output
rlabel metal1 s 1324 242 1426 298 1 ZN
port 3 nsew default output
rlabel metal1 s 1324 136 1370 242 1 ZN
port 3 nsew default output
rlabel metal1 s 1558 870 1604 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1150 870 1196 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 274 870 320 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1558 680 1604 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 274 680 320 870 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1548 90 1594 204 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1100 90 1146 204 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 284 90 330 204 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1904 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1904 1008
string GDS_END 929554
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 923694
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
