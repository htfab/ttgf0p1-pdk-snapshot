magic
tech gf180mcuD
magscale 1 10
timestamp 1753371985
<< nwell >>
rect -86 354 1206 870
<< pwell >>
rect -86 -86 1206 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 756 68 812 268
rect 916 68 972 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
<< ndiff >>
rect 28 127 116 268
rect 28 81 41 127
rect 87 81 116 127
rect 28 68 116 81
rect 172 68 276 268
rect 332 251 436 268
rect 332 205 361 251
rect 407 205 436 251
rect 332 68 436 205
rect 492 68 596 268
rect 652 127 756 268
rect 652 81 681 127
rect 727 81 756 127
rect 652 68 756 81
rect 812 251 916 268
rect 812 205 841 251
rect 887 205 916 251
rect 812 68 916 205
rect 972 127 1062 268
rect 972 81 1001 127
rect 1047 81 1062 127
rect 972 68 1062 81
<< pdiff >>
rect 28 600 116 716
rect 28 554 41 600
rect 87 554 116 600
rect 28 440 116 554
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 600 436 716
rect 332 554 361 600
rect 407 554 436 600
rect 332 440 436 554
rect 492 703 596 716
rect 492 657 521 703
rect 567 657 596 703
rect 492 440 596 657
rect 652 639 756 716
rect 652 593 681 639
rect 727 593 756 639
rect 652 440 756 593
rect 812 499 916 716
rect 812 453 841 499
rect 887 453 916 499
rect 812 440 916 453
rect 972 652 1062 716
rect 972 606 1001 652
rect 1047 606 1062 652
rect 972 440 1062 606
<< ndiffc >>
rect 41 81 87 127
rect 361 205 407 251
rect 681 81 727 127
rect 841 205 887 251
rect 1001 81 1047 127
<< pdiffc >>
rect 41 554 87 600
rect 201 657 247 703
rect 361 554 407 600
rect 521 657 567 703
rect 681 593 727 639
rect 841 453 887 499
rect 1001 606 1047 652
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 116 390 172 440
rect 91 377 172 390
rect 91 331 107 377
rect 153 331 172 377
rect 91 318 172 331
rect 116 268 172 318
rect 276 390 332 440
rect 436 390 492 440
rect 276 377 492 390
rect 596 386 652 440
rect 276 331 289 377
rect 479 331 492 377
rect 276 318 492 331
rect 276 268 332 318
rect 436 268 492 318
rect 572 373 653 386
rect 572 327 590 373
rect 636 327 653 373
rect 572 314 653 327
rect 756 373 812 440
rect 916 392 972 440
rect 916 375 1025 392
rect 916 373 964 375
rect 756 329 964 373
rect 1010 329 1025 375
rect 756 327 1025 329
rect 596 268 652 314
rect 756 268 812 327
rect 916 313 1025 327
rect 916 268 972 313
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
<< polycontact >>
rect 107 331 153 377
rect 289 331 479 377
rect 590 327 636 373
rect 964 329 1010 375
<< metal1 >>
rect 0 724 1120 844
rect 201 703 247 724
rect 201 646 247 657
rect 521 703 567 724
rect 521 646 567 657
rect 681 652 1047 678
rect 681 639 1001 652
rect 41 600 87 616
rect 87 554 361 600
rect 407 593 681 600
rect 727 632 1001 639
rect 1001 594 1047 606
rect 407 554 727 593
rect 41 539 87 554
rect 129 462 618 508
rect 129 391 175 462
rect 91 377 175 391
rect 91 331 107 377
rect 153 331 175 377
rect 91 318 175 331
rect 276 377 492 390
rect 276 331 289 377
rect 479 331 492 377
rect 276 318 492 331
rect 572 386 618 462
rect 829 499 887 524
rect 829 453 841 499
rect 572 373 653 386
rect 572 327 590 373
rect 636 327 653 373
rect 572 314 653 327
rect 829 251 887 453
rect 947 375 1025 462
rect 947 329 964 375
rect 1010 329 1025 375
rect 947 313 1025 329
rect 336 205 361 251
rect 407 205 841 251
rect 887 205 898 251
rect 41 127 87 138
rect 41 60 87 81
rect 681 127 727 138
rect 681 60 727 81
rect 1001 127 1047 138
rect 1001 60 1047 81
rect 0 -60 1120 60
<< labels >>
flabel metal1 s 0 724 1120 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1120 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 829 205 887 524 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 947 313 1025 462 0 FreeSans 200 0 0 0 C
port 6 nsew signal input
flabel metal1 276 318 492 390 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel metal1 91 318 175 391 0 FreeSans 200 0 0 0 A
port 8 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1120 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
