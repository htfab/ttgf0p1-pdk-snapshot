VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO nsnrlatch_x0
  CLASS BLOCK ;
  FOREIGN nsnrlatch_x0 ;
  ORIGIN 0.430 0.000 ;
  SIZE 5.420 BY 7.430 ;
  PIN q
    ANTENNAGATEAREA 0.492800 ;
    ANTENNADIFFAREA 0.844800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.700 5.090 1.255 5.430 ;
        RECT 0.700 3.900 0.960 5.090 ;
        RECT 0.700 3.560 2.215 3.900 ;
        RECT 0.700 1.910 0.960 3.560 ;
        RECT 0.225 1.570 0.960 1.910 ;
    END
  END q
  PIN vdd
    ANTENNADIFFAREA 2.772800 ;
    PORT
      LAYER Nwell ;
        RECT -0.430 3.400 4.990 7.430 ;
      LAYER Metal1 ;
        RECT 0.000 5.660 4.560 7.000 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 1.998400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 4.560 1.340 ;
    END
  END vss
  PIN nset
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.210 2.140 0.470 5.430 ;
    END
  END nset
  PIN nq
    ANTENNAGATEAREA 0.492800 ;
    ANTENNADIFFAREA 0.844800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.610 3.240 2.870 5.430 ;
        RECT 1.205 2.900 2.870 3.240 ;
        RECT 2.610 1.910 2.870 2.900 ;
        RECT 2.610 1.570 3.655 1.910 ;
    END
  END nq
  PIN nrst
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 3.100 2.140 3.360 5.430 ;
    END
  END nrst
END nsnrlatch_x0
END LIBRARY

