magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
use M1_NWELL4310590548733_128x8m81  M1_NWELL4310590548733_128x8m81_0
timestamp 1755005639
transform 1 0 887 0 1 2626
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_0
timestamp 1755005639
transform 1 0 296 0 1 2790
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_1
timestamp 1755005639
transform 1 0 296 0 1 2268
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_0
timestamp 1755005639
transform 1 0 1170 0 1 2821
box 0 0 1 1
use M1_POLY24310590548734_128x8m81  M1_POLY24310590548734_128x8m81_1
timestamp 1755005639
transform 1 0 1170 0 1 2310
box 0 0 1 1
use M2_M14310590548751_128x8m81  M2_M14310590548751_128x8m81_0
timestamp 1755005639
transform 1 0 874 0 1 6580
box 0 0 1 1
use M2_M14310590548751_128x8m81  M2_M14310590548751_128x8m81_1
timestamp 1755005639
transform 1 0 1322 0 1 6580
box 0 0 1 1
use M2_M14310590548751_128x8m81  M2_M14310590548751_128x8m81_2
timestamp 1755005639
transform 1 0 202 0 1 6580
box 0 0 1 1
use M2_M14310590548753_128x8m81  M2_M14310590548753_128x8m81_0
timestamp 1755005639
transform 1 0 1098 0 1 1994
box 0 0 1 1
use M2_M14310590548753_128x8m81  M2_M14310590548753_128x8m81_1
timestamp 1755005639
transform 1 0 650 0 1 1994
box 0 0 1 1
use M2_M14310590548754_128x8m81  M2_M14310590548754_128x8m81_0
timestamp 1755005639
transform 1 0 218 0 1 2271
box 0 0 1 1
use M2_M14310590548755_128x8m81  M2_M14310590548755_128x8m81_0
timestamp 1755005639
transform 1 0 1098 0 1 4302
box 0 0 1 1
use M2_M14310590548755_128x8m81  M2_M14310590548755_128x8m81_1
timestamp 1755005639
transform 1 0 650 0 1 4302
box 0 0 1 1
use M3_M24310590548752_128x8m81  M3_M24310590548752_128x8m81_0
timestamp 1755005639
transform 1 0 202 0 1 6580
box 0 0 1 1
use M3_M24310590548752_128x8m81  M3_M24310590548752_128x8m81_1
timestamp 1755005639
transform 1 0 1322 0 1 6580
box 0 0 1 1
use M3_M24310590548752_128x8m81  M3_M24310590548752_128x8m81_2
timestamp 1755005639
transform 1 0 874 0 1 6580
box 0 0 1 1
use nmos_5p04310590548758_128x8m81  nmos_5p04310590548758_128x8m81_0
timestamp 1755005639
transform 1 0 926 0 1 340
box 0 0 1 1
use nmos_5p04310590548758_128x8m81  nmos_5p04310590548758_128x8m81_1
timestamp 1755005639
transform 1 0 702 0 1 340
box 0 0 1 1
use nmos_5p04310590548758_128x8m81  nmos_5p04310590548758_128x8m81_2
timestamp 1755005639
transform 1 0 254 0 1 340
box 0 0 1 1
use nmos_5p04310590548758_128x8m81  nmos_5p04310590548758_128x8m81_3
timestamp 1755005639
transform 1 0 1150 0 1 340
box 0 0 1 1
use pmos_5p04310590548759_128x8m81  pmos_5p04310590548759_128x8m81_0
timestamp 1755005639
transform 1 0 254 0 1 2971
box 0 0 1 1
use pmos_5p04310590548759_128x8m81  pmos_5p04310590548759_128x8m81_1
timestamp 1755005639
transform 1 0 702 0 1 2971
box 0 0 1 1
use pmos_5p04310590548759_128x8m81  pmos_5p04310590548759_128x8m81_2
timestamp 1755005639
transform 1 0 926 0 1 2971
box 0 0 1 1
use pmos_5p04310590548759_128x8m81  pmos_5p04310590548759_128x8m81_3
timestamp 1755005639
transform 1 0 1150 0 1 2971
box 0 0 1 1
<< properties >>
string GDS_END 846104
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 842830
string path 4.370 15.035 4.370 13.055 
<< end >>
