magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 534 1094
<< pwell >>
rect -86 -86 534 453
<< metal1 >>
rect 0 918 448 1098
rect 49 710 95 918
rect 126 366 194 506
rect 49 90 95 257
rect 142 242 194 366
rect 253 189 319 872
rect 0 -90 448 90
<< labels >>
rlabel metal1 s 142 242 194 366 6 I
port 1 nsew default input
rlabel metal1 s 126 366 194 506 6 I
port 1 nsew default input
rlabel metal1 s 253 189 319 872 6 ZN
port 2 nsew default output
rlabel metal1 s 49 710 95 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 918 448 1098 6 VDD
port 3 nsew power bidirectional abutment
rlabel nwell s -86 453 534 1094 6 VNW
port 4 nsew power bidirectional
rlabel pwell s -86 -86 534 453 6 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 0 -90 448 90 8 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 257 6 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 448 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1443454
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1441240
<< end >>
