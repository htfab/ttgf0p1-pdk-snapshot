* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__aoi31_2.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__aoi31_2 VDD VNW VPW VSS A B C Y D
X0 a_28_440# A VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X1 VSS D Y VPW nfet_03v3 ad=0.2625p pd=1.525u as=0.26p ps=1.52u w=1u l=0.28u
X2 VSS A a_28_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X3 a_28_440# C VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X4 Y C a_492_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X5 VDD B a_28_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X6 a_28_68# B a_492_68# VPW nfet_03v3 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.28u
X7 Y D a_28_440# VNW pfet_03v3 ad=0.36225p pd=1.905u as=0.3588p ps=1.9u w=1.38u l=0.28u
X8 a_28_440# B VDD VNW pfet_03v3 ad=0.8004p pd=2.54u as=0.3588p ps=1.9u w=1.38u l=0.28u
X9 VDD C a_28_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.8004p ps=2.54u w=1.38u l=0.28u
X10 a_492_68# C Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.28u
X11 a_492_68# B a_28_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X12 Y D VSS VPW nfet_03v3 ad=0.44p pd=2.88u as=0.2625p ps=1.525u w=1u l=0.28u
X13 VDD A a_28_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X14 a_28_440# D Y VNW pfet_03v3 ad=0.6072p pd=3.64u as=0.36225p ps=1.905u w=1.38u l=0.28u
X15 a_28_68# A VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
.ends

