magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 1226 1486
<< nmos >>
rect 120 209 176 385
rect 280 209 336 385
rect 440 209 496 385
rect 600 209 656 385
rect 804 209 860 584
<< pmos >>
rect 120 1015 176 1191
rect 280 1015 336 1191
rect 440 1015 496 1191
rect 600 1015 656 1191
rect 804 776 860 1191
<< ndiff >>
rect 716 385 804 584
rect 32 268 120 385
rect 32 222 45 268
rect 91 222 120 268
rect 32 209 120 222
rect 176 371 280 385
rect 176 325 205 371
rect 251 325 280 371
rect 176 209 280 325
rect 336 268 440 385
rect 336 222 365 268
rect 411 222 440 268
rect 336 209 440 222
rect 496 371 600 385
rect 496 325 525 371
rect 571 325 600 371
rect 496 209 600 325
rect 656 268 804 385
rect 656 222 729 268
rect 775 222 804 268
rect 656 209 804 222
rect 860 571 948 584
rect 860 325 889 571
rect 935 325 948 571
rect 860 209 948 325
<< pdiff >>
rect 32 1075 120 1191
rect 32 1029 45 1075
rect 91 1029 120 1075
rect 32 1015 120 1029
rect 176 1015 280 1191
rect 336 1015 440 1191
rect 496 1015 600 1191
rect 656 1178 804 1191
rect 656 1132 729 1178
rect 775 1132 804 1178
rect 656 1015 804 1132
rect 716 776 804 1015
rect 860 1055 948 1191
rect 860 809 889 1055
rect 935 809 948 1055
rect 860 776 948 809
<< ndiffc >>
rect 45 222 91 268
rect 205 325 251 371
rect 365 222 411 268
rect 525 325 571 371
rect 729 222 775 268
rect 889 325 935 571
<< pdiffc >>
rect 45 1029 91 1075
rect 729 1132 775 1178
rect 889 809 935 1055
<< psubdiff >>
rect 28 87 1112 100
rect 28 41 47 87
rect 1093 41 1112 87
rect 28 28 1112 41
<< nsubdiff >>
rect 28 1359 1112 1372
rect 28 1313 47 1359
rect 1093 1313 1112 1359
rect 28 1300 1112 1313
<< psubdiffcont >>
rect 47 41 1093 87
<< nsubdiffcont >>
rect 47 1313 1093 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 600 1191 656 1235
rect 804 1191 860 1235
rect 120 716 176 1015
rect 280 716 336 1015
rect 440 716 496 1015
rect 600 716 656 1015
rect 804 716 860 776
rect 32 703 176 716
rect 32 657 45 703
rect 91 657 176 703
rect 32 644 176 657
rect 224 703 336 716
rect 224 657 237 703
rect 283 657 336 703
rect 224 644 336 657
rect 384 703 496 716
rect 384 657 397 703
rect 443 657 496 703
rect 384 644 496 657
rect 544 703 656 716
rect 544 657 557 703
rect 603 657 656 703
rect 544 644 656 657
rect 704 703 860 716
rect 704 657 717 703
rect 763 657 860 703
rect 704 644 860 657
rect 120 385 176 644
rect 280 385 336 644
rect 440 385 496 644
rect 600 385 656 644
rect 804 584 860 644
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
rect 600 165 656 209
rect 804 165 860 209
<< polycontact >>
rect 45 657 91 703
rect 237 657 283 703
rect 397 657 443 703
rect 557 657 603 703
rect 717 657 763 703
<< metal1 >>
rect 0 1359 1140 1400
rect 0 1313 47 1359
rect 1093 1313 1140 1359
rect 0 1178 1140 1313
rect 0 1132 729 1178
rect 775 1132 1140 1178
rect 45 1075 766 1086
rect 91 1029 766 1075
rect 45 1018 766 1029
rect 42 703 94 972
rect 42 657 45 703
rect 91 657 94 703
rect 42 314 94 657
rect 234 703 286 972
rect 234 657 237 703
rect 283 657 286 703
rect 234 428 286 657
rect 394 703 446 972
rect 394 657 397 703
rect 443 657 446 703
rect 394 428 446 657
rect 554 703 606 972
rect 554 657 557 703
rect 603 657 606 703
rect 554 428 606 657
rect 714 703 766 1018
rect 714 657 717 703
rect 763 657 766 703
rect 714 382 766 657
rect 205 371 766 382
rect 251 325 525 371
rect 571 325 766 371
rect 205 314 766 325
rect 886 1055 938 1086
rect 886 809 889 1055
rect 935 809 938 1055
rect 886 571 938 809
rect 886 325 889 571
rect 935 325 938 571
rect 886 314 938 325
rect 0 222 45 268
rect 91 222 365 268
rect 411 222 729 268
rect 775 222 1140 268
rect 0 87 1140 222
rect 0 41 47 87
rect 1093 41 1140 87
rect 0 0 1140 41
<< labels >>
rlabel metal1 s 0 0 1140 268 4 vss
port 3 nsew
rlabel metal1 s 0 1132 1140 1400 4 vdd
port 5 nsew
rlabel metal1 s 42 314 94 972 4 i0
port 7 nsew
rlabel metal1 s 234 428 286 972 4 i1
port 9 nsew
rlabel metal1 s 394 428 446 972 4 i2
port 11 nsew
rlabel metal1 s 554 428 606 972 4 i3
port 13 nsew
rlabel metal1 s 886 314 938 1086 4 q
port 15 nsew
<< end >>
