magic
tech gf180mcuD
timestamp 1755005639
<< properties >>
string GDS_END 253850
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 252826
<< end >>
