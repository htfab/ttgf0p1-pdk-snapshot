magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 1430 1094
<< pwell >>
rect -86 -86 1430 453
<< metal1 >>
rect 0 918 1344 1098
rect 69 710 115 918
rect 731 603 777 872
rect 1149 710 1195 918
rect 731 557 991 603
rect 142 443 203 542
rect 360 454 428 542
rect 584 454 652 542
rect 49 90 95 316
rect 497 90 543 316
rect 814 354 866 511
rect 926 228 991 557
rect 1038 354 1090 511
rect 0 -90 1344 90
<< obsm1 >>
rect 273 362 767 408
rect 273 154 319 362
rect 721 182 767 362
rect 1169 182 1215 316
rect 721 136 1215 182
<< labels >>
rlabel metal1 s 584 454 652 542 6 A1
port 1 nsew default input
rlabel metal1 s 360 454 428 542 6 A2
port 2 nsew default input
rlabel metal1 s 142 443 203 542 6 A3
port 3 nsew default input
rlabel metal1 s 814 354 866 511 6 B1
port 4 nsew default input
rlabel metal1 s 1038 354 1090 511 6 B2
port 5 nsew default input
rlabel metal1 s 926 228 991 557 6 ZN
port 6 nsew default output
rlabel metal1 s 731 557 991 603 6 ZN
port 6 nsew default output
rlabel metal1 s 731 603 777 872 6 ZN
port 6 nsew default output
rlabel metal1 s 1149 710 1195 918 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 69 710 115 918 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 918 1344 1098 6 VDD
port 7 nsew power bidirectional abutment
rlabel nwell s -86 453 1430 1094 6 VNW
port 8 nsew power bidirectional
rlabel pwell s -86 -86 1430 453 6 VPW
port 9 nsew ground bidirectional
rlabel metal1 s 0 -90 1344 90 8 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 316 6 VSS
port 10 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 316 6 VSS
port 10 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1344 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 166272
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 162082
<< end >>
