* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__xnor2_4.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__xnor2_4 VDD VNW VPW VSS B A Y
X0 VSS a_556_68# Y VPW nfet_03v3 ad=0.26p pd=1.52u as=0.285p ps=1.57u w=1u l=0.28u
X1 VDD a_556_68# Y VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3933p ps=1.95u w=1.38u l=0.28u
X2 Y a_556_68# VSS VPW nfet_03v3 ad=0.285p pd=1.57u as=0.26p ps=1.52u w=1u l=0.28u
X3 a_332_440# A VDD VNW pfet_03v3 ad=0.5796p pd=2.22u as=0.3588p ps=1.9u w=1.38u l=0.28u
X4 VSS A a_28_68# VPW nfet_03v3 ad=0.54p pd=2.08u as=0.44p ps=2.88u w=1u l=0.28u
X5 a_556_68# a_500_24# a_444_68# VPW nfet_03v3 ad=0.62p pd=2.24u as=0.14p ps=1.28u w=1u l=0.28u
X6 Y a_556_68# VDD VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.3588p ps=1.9u w=1.38u l=0.28u
X7 a_500_24# A a_556_68# VPW nfet_03v3 ad=0.31p pd=1.62u as=0.62p ps=2.24u w=1u l=0.28u
X8 a_500_24# a_28_68# a_556_68# VNW pfet_03v3 ad=0.7866p pd=2.52u as=0.4968p ps=2.1u w=1.38u l=0.28u
X9 VDD B a_500_24# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.7866p ps=2.52u w=1.38u l=0.28u
X10 VSS B a_500_24# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.31p ps=1.62u w=1u l=0.28u
X11 VSS a_556_68# Y VPW nfet_03v3 ad=0.56p pd=3.12u as=0.26p ps=1.52u w=1u l=0.28u
X12 VDD a_556_68# Y VNW pfet_03v3 ad=0.7314p pd=3.82u as=0.3588p ps=1.9u w=1.38u l=0.28u
X13 a_444_68# a_28_68# VSS VPW nfet_03v3 ad=0.14p pd=1.28u as=0.54p ps=2.08u w=1u l=0.28u
X14 Y a_556_68# VSS VPW nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.28u
X15 Y a_556_68# VDD VNW pfet_03v3 ad=0.3933p pd=1.95u as=0.3588p ps=1.9u w=1.38u l=0.28u
X16 VDD A a_28_68# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.6072p ps=3.64u w=1.38u l=0.28u
X17 a_556_68# a_500_24# a_332_440# VNW pfet_03v3 ad=0.4968p pd=2.1u as=0.5796p ps=2.22u w=1.38u l=0.28u
.ends

