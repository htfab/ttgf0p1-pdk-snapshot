* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__diode_2.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__diode_2 VDD VNW VPW VSS DIODE
D0 DIODE VNW diode_pd2nw_03v3 pj=1.93u area=0.2295p
D1 VPW DIODE diode_nd2ps_03v3 pj=1.83u area=0.209p
.ends

