magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< psubdiff >>
rect 13097 70975 69968 71000
rect 13097 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69968 70975
rect 13097 70871 69968 70929
rect 13097 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69968 70871
rect 13097 70803 69968 70825
rect 13097 70767 13291 70803
rect 13097 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13291 70767
rect 13097 70663 13291 70721
rect 13097 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13291 70663
rect 13097 70559 13291 70617
rect 13097 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13291 70559
rect 13097 70455 13291 70513
rect 13097 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13291 70455
rect 13097 70351 13291 70409
rect 13097 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13291 70351
rect 13097 70247 13291 70305
rect 13097 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13291 70247
rect 13097 70143 13291 70201
rect 13097 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13291 70143
rect 13097 70039 13291 70097
rect 13097 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13291 70039
rect 13097 69935 13291 69993
rect 13097 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13291 69935
rect 13097 69831 13291 69889
rect 13097 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13291 69831
rect 13097 69727 13291 69785
rect 69774 70720 69968 70803
rect 69774 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69968 70720
rect 69774 70616 69968 70674
rect 69774 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69968 70616
rect 69774 70512 69968 70570
rect 69774 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69968 70512
rect 69774 70408 69968 70466
rect 69774 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69968 70408
rect 69774 70304 69968 70362
rect 69774 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69968 70304
rect 69774 70200 69968 70258
rect 69774 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69968 70200
rect 69774 70096 69968 70154
rect 69774 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69968 70096
rect 69774 69968 69968 70050
rect 69774 69946 71000 69968
rect 69774 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69774 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69774 69842 71000 69862
rect 69774 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69774 69774 70824 69796
rect 13097 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13291 69727
rect 13097 69623 13291 69681
rect 13097 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13291 69623
rect 13097 69519 13291 69577
rect 13097 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13291 69519
rect 13097 69415 13291 69473
rect 13097 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13291 69415
rect 13097 69311 13291 69369
rect 13097 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13291 69311
rect 13097 69207 13291 69265
rect 13097 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13291 69207
rect 13097 69103 13291 69161
rect 13097 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13291 69103
rect 13097 68999 13291 69057
rect 13097 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13291 68999
rect 13097 68895 13291 68953
rect 13097 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13291 68895
rect 13097 68791 13291 68849
rect 13097 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13291 68791
rect 13097 68687 13291 68745
rect 13097 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13291 68687
rect 13097 68583 13291 68641
rect 13097 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13291 68583
rect 13097 68479 13291 68537
rect 13097 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13291 68479
rect 13097 68375 13291 68433
rect 13097 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13291 68375
rect 13097 68271 13291 68329
rect 13097 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13291 68271
rect 13097 68167 13291 68225
rect 13097 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13291 68167
rect 13097 68063 13291 68121
rect 13097 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13291 68063
rect 13097 67959 13291 68017
rect 13097 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13291 67959
rect 13097 67855 13291 67913
rect 13097 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13291 67855
rect 13097 67751 13291 67809
rect 13097 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13291 67751
rect 13097 67647 13291 67705
rect 13097 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13291 67647
rect 13097 67543 13291 67601
rect 13097 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13291 67543
rect 13097 67439 13291 67497
rect 13097 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13291 67439
rect 13097 67335 13291 67393
rect 13097 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13291 67335
rect 13097 67231 13291 67289
rect 13097 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13291 67231
rect 13097 67127 13291 67185
rect 13097 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13291 67127
rect 13097 67023 13291 67081
rect 13097 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13291 67023
rect 13097 66919 13291 66977
rect 13097 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13291 66919
rect 13097 66815 13291 66873
rect 13097 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13291 66815
rect 13097 66711 13291 66769
rect 13097 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13291 66711
rect 13097 66607 13291 66665
rect 13097 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13291 66607
rect 13097 66503 13291 66561
rect 13097 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13291 66503
rect 13097 66399 13291 66457
rect 13097 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13291 66399
rect 13097 66295 13291 66353
rect 13097 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13291 66295
rect 13097 66191 13291 66249
rect 13097 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13291 66191
rect 13097 66087 13291 66145
rect 13097 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13291 66087
rect 13097 65983 13291 66041
rect 13097 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13291 65983
rect 13097 65879 13291 65937
rect 13097 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13291 65879
rect 13097 65775 13291 65833
rect 13097 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13291 65775
rect 13097 65671 13291 65729
rect 13097 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13291 65671
rect 13097 65567 13291 65625
rect 13097 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13291 65567
rect 13097 65463 13291 65521
rect 13097 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13291 65463
rect 13097 65359 13291 65417
rect 13097 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13291 65359
rect 13097 65255 13291 65313
rect 13097 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13291 65255
rect 13097 65151 13291 65209
rect 13097 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13291 65151
rect 13097 65047 13291 65105
rect 13097 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13291 65047
rect 13097 64943 13291 65001
rect 13097 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13291 64943
rect 13097 64839 13291 64897
rect 13097 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13291 64839
rect 13097 64735 13291 64793
rect 13097 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13291 64735
rect 13097 64631 13291 64689
rect 13097 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13291 64631
rect 13097 64527 13291 64585
rect 13097 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13291 64527
rect 13097 64423 13291 64481
rect 13097 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13291 64423
rect 13097 64319 13291 64377
rect 13097 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13291 64319
rect 13097 64215 13291 64273
rect 13097 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13291 64215
rect 13097 64111 13291 64169
rect 13097 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13291 64111
rect 13097 64007 13291 64065
rect 13097 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13291 64007
rect 13097 63903 13291 63961
rect 13097 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13291 63903
rect 13097 63799 13291 63857
rect 13097 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13291 63799
rect 13097 63695 13291 63753
rect 13097 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13291 63695
rect 13097 63591 13291 63649
rect 13097 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13291 63591
rect 13097 63487 13291 63545
rect 13097 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13291 63487
rect 13097 63383 13291 63441
rect 13097 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13291 63383
rect 13097 63279 13291 63337
rect 13097 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13291 63279
rect 13097 63175 13291 63233
rect 13097 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13291 63175
rect 13097 63071 13291 63129
rect 13097 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13291 63071
rect 13097 62967 13291 63025
rect 13097 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13291 62967
rect 13097 62863 13291 62921
rect 13097 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13291 62863
rect 13097 62759 13291 62817
rect 13097 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13291 62759
rect 13097 62655 13291 62713
rect 13097 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13291 62655
rect 13097 62551 13291 62609
rect 13097 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13291 62551
rect 13097 62447 13291 62505
rect 13097 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13291 62447
rect 13097 62343 13291 62401
rect 13097 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13291 62343
rect 13097 62239 13291 62297
rect 13097 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13291 62239
rect 13097 62135 13291 62193
rect 13097 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13291 62135
rect 13097 62031 13291 62089
rect 13097 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13291 62031
rect 13097 61927 13291 61985
rect 13097 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13291 61927
rect 13097 61823 13291 61881
rect 13097 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13291 61823
rect 13097 61719 13291 61777
rect 13097 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13291 61719
rect 13097 61615 13291 61673
rect 13097 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13291 61615
rect 13097 61511 13291 61569
rect 13097 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13291 61511
rect 13097 61407 13291 61465
rect 13097 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13291 61407
rect 13097 61303 13291 61361
rect 13097 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13291 61303
rect 13097 61199 13291 61257
rect 13097 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13291 61199
rect 13097 61095 13291 61153
rect 13097 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13291 61095
rect 13097 60991 13291 61049
rect 13097 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13291 60991
rect 13097 60887 13291 60945
rect 13097 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13291 60887
rect 13097 60783 13291 60841
rect 13097 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13291 60783
rect 13097 60679 13291 60737
rect 13097 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13291 60679
rect 13097 60575 13291 60633
rect 13097 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13291 60575
rect 13097 60471 13291 60529
rect 13097 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13291 60471
rect 13097 60367 13291 60425
rect 13097 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13291 60367
rect 13097 60263 13291 60321
rect 13097 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13291 60263
rect 13097 60159 13291 60217
rect 13097 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13291 60159
rect 13097 60055 13291 60113
rect 13097 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13291 60055
rect 13097 59951 13291 60009
rect 13097 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13291 59951
rect 13097 59847 13291 59905
rect 13097 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13291 59847
rect 13097 59743 13291 59801
rect 13097 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13291 59743
rect 13097 59639 13291 59697
rect 13097 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13291 59639
rect 13097 59535 13291 59593
rect 13097 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13291 59535
rect 13097 59431 13291 59489
rect 13097 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13291 59431
rect 13097 59327 13291 59385
rect 13097 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13291 59327
rect 13097 59223 13291 59281
rect 13097 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13291 59223
rect 13097 59119 13291 59177
rect 13097 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13291 59119
rect 13097 59015 13291 59073
rect 13097 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13291 59015
rect 13097 58911 13291 58969
rect 13097 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13291 58911
rect 13097 58807 13291 58865
rect 13097 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13291 58807
rect 13097 58703 13291 58761
rect 13097 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13291 58703
rect 13097 58599 13291 58657
rect 13097 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13291 58599
rect 13097 58495 13291 58553
rect 13097 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13291 58495
rect 13097 58391 13291 58449
rect 13097 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13291 58391
rect 13097 58287 13291 58345
rect 13097 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13291 58287
rect 13097 58183 13291 58241
rect 13097 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13291 58183
rect 13097 58079 13291 58137
rect 13097 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13291 58079
rect 13097 57975 13291 58033
rect 13097 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13291 57975
rect 13097 57871 13291 57929
rect 13097 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13291 57871
rect 13097 57767 13291 57825
rect 13097 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13291 57767
rect 13097 57663 13291 57721
rect 13097 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13291 57663
rect 13097 57559 13291 57617
rect 13097 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13291 57559
rect 13097 57455 13291 57513
rect 13097 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13291 57455
rect 13097 57351 13291 57409
rect 13097 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13291 57351
rect 13097 57247 13291 57305
rect 13097 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13291 57247
rect 13097 57143 13291 57201
rect 13097 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13291 57143
rect 13097 57039 13291 57097
rect 13097 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13291 57039
rect 13097 56935 13291 56993
rect 13097 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13291 56935
rect 13097 56831 13291 56889
rect 13097 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13291 56831
rect 13097 56727 13291 56785
rect 13097 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13291 56727
rect 13097 56623 13291 56681
rect 13097 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13291 56623
rect 13097 56519 13291 56577
rect 13097 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13291 56519
rect 13097 56415 13291 56473
rect 13097 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13291 56415
rect 13097 56311 13291 56369
rect 13097 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13291 56311
rect 13097 56207 13291 56265
rect 13097 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13291 56207
rect 13097 56103 13291 56161
rect 13097 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13291 56103
rect 13097 55999 13291 56057
rect 13097 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13291 55999
rect 13097 55895 13291 55953
rect 13097 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13291 55895
rect 13097 55791 13291 55849
rect 13097 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13291 55791
rect 13097 55687 13291 55745
rect 13097 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13291 55687
rect 13097 55583 13291 55641
rect 13097 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13291 55583
rect 13097 55479 13291 55537
rect 13097 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13291 55479
rect 13097 55375 13291 55433
rect 13097 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13291 55375
rect 13097 55271 13291 55329
rect 13097 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13291 55271
rect 13097 55167 13291 55225
rect 13097 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13291 55167
rect 13097 55063 13291 55121
rect 13097 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13291 55063
rect 13097 54959 13291 55017
rect 13097 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13291 54959
rect 13097 54855 13291 54913
rect 13097 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13291 54855
rect 13097 54751 13291 54809
rect 13097 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13291 54751
rect 13097 54647 13291 54705
rect 13097 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13291 54647
rect 13097 54543 13291 54601
rect 13097 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13291 54543
rect 13097 54439 13291 54497
rect 13097 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13291 54439
rect 13097 54335 13291 54393
rect 13097 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13291 54335
rect 13097 54231 13291 54289
rect 13097 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13291 54231
rect 13097 54127 13291 54185
rect 13097 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13291 54127
rect 13097 54023 13291 54081
rect 13097 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13291 54023
rect 13097 53919 13291 53977
rect 13097 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13291 53919
rect 13097 53815 13291 53873
rect 13097 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13291 53815
rect 13097 53711 13291 53769
rect 13097 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13291 53711
rect 13097 53607 13291 53665
rect 13097 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13291 53607
rect 13097 53503 13291 53561
rect 13097 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13291 53503
rect 13097 53399 13291 53457
rect 13097 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13291 53399
rect 13097 53295 13291 53353
rect 13097 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13291 53295
rect 13097 53191 13291 53249
rect 13097 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13291 53191
rect 13097 53087 13291 53145
rect 13097 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13291 53087
rect 13097 52983 13291 53041
rect 13097 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13291 52983
rect 13097 52879 13291 52937
rect 13097 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13291 52879
rect 13097 52775 13291 52833
rect 13097 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13291 52775
rect 13097 52671 13291 52729
rect 13097 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13291 52671
rect 13097 52567 13291 52625
rect 13097 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13291 52567
rect 13097 52463 13291 52521
rect 13097 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13291 52463
rect 13097 52359 13291 52417
rect 13097 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13291 52359
rect 13097 52255 13291 52313
rect 13097 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13291 52255
rect 13097 52151 13291 52209
rect 13097 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13291 52151
rect 13097 52047 13291 52105
rect 13097 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13291 52047
rect 13097 51943 13291 52001
rect 13097 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13291 51943
rect 13097 51839 13291 51897
rect 13097 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13291 51839
rect 13097 51735 13291 51793
rect 13097 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13291 51735
rect 13097 51631 13291 51689
rect 13097 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13291 51631
rect 13097 51527 13291 51585
rect 13097 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13291 51527
rect 13097 51423 13291 51481
rect 13097 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13291 51423
rect 13097 51319 13291 51377
rect 13097 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13291 51319
rect 13097 51215 13291 51273
rect 13097 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13291 51215
rect 13097 51111 13291 51169
rect 13097 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13291 51111
rect 13097 51007 13291 51065
rect 13097 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13291 51007
rect 13097 50903 13291 50961
rect 13097 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13291 50903
rect 13097 50799 13291 50857
rect 13097 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13291 50799
rect 13097 50695 13291 50753
rect 13097 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13291 50695
rect 13097 50591 13291 50649
rect 13097 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13291 50591
rect 13097 50487 13291 50545
rect 13097 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13291 50487
rect 13097 50383 13291 50441
rect 13097 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13291 50383
rect 13097 50279 13291 50337
rect 13097 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13291 50279
rect 13097 50175 13291 50233
rect 13097 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13291 50175
rect 13097 50071 13291 50129
rect 13097 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13291 50071
rect 13097 49967 13291 50025
rect 13097 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13291 49967
rect 13097 49863 13291 49921
rect 13097 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13291 49863
rect 13097 49759 13291 49817
rect 13097 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13291 49759
rect 13097 49655 13291 49713
rect 13097 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13291 49655
rect 13097 49551 13291 49609
rect 13097 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13291 49551
rect 13097 49447 13291 49505
rect 13097 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13291 49447
rect 13097 49343 13291 49401
rect 13097 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13291 49343
rect 13097 49239 13291 49297
rect 13097 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13291 49239
rect 13097 49135 13291 49193
rect 13097 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13291 49135
rect 13097 49031 13291 49089
rect 13097 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13291 49031
rect 13097 48927 13291 48985
rect 13097 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13291 48927
rect 13097 48823 13291 48881
rect 13097 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13291 48823
rect 13097 48719 13291 48777
rect 13097 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13291 48719
rect 13097 48615 13291 48673
rect 13097 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13291 48615
rect 13097 48511 13291 48569
rect 13097 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13291 48511
rect 13097 48407 13291 48465
rect 13097 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13291 48407
rect 13097 48303 13291 48361
rect 13097 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13291 48303
rect 13097 48199 13291 48257
rect 13097 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13291 48199
rect 13097 48095 13291 48153
rect 13097 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13291 48095
rect 13097 47991 13291 48049
rect 13097 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13291 47991
rect 13097 47887 13291 47945
rect 13097 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13291 47887
rect 13097 47783 13291 47841
rect 13097 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13291 47783
rect 13097 47679 13291 47737
rect 13097 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13291 47679
rect 13097 47575 13291 47633
rect 13097 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13291 47575
rect 13097 47471 13291 47529
rect 13097 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13291 47471
rect 13097 47367 13291 47425
rect 13097 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13291 47367
rect 13097 47263 13291 47321
rect 13097 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13291 47263
rect 13097 47159 13291 47217
rect 13097 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13291 47159
rect 13097 47055 13291 47113
rect 13097 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13291 47055
rect 13097 46951 13291 47009
rect 13097 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13291 46951
rect 13097 46847 13291 46905
rect 13097 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13291 46847
rect 13097 46743 13291 46801
rect 13097 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13291 46743
rect 13097 46639 13291 46697
rect 13097 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13291 46639
rect 13097 46535 13291 46593
rect 13097 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13291 46535
rect 13097 46431 13291 46489
rect 13097 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13291 46431
rect 13097 46327 13291 46385
rect 13097 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13291 46327
rect 13097 46223 13291 46281
rect 13097 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13291 46223
rect 13097 46119 13291 46177
rect 13097 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13291 46119
rect 13097 46015 13291 46073
rect 13097 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13291 46015
rect 13097 45911 13291 45969
rect 13097 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13291 45911
rect 13097 45807 13291 45865
rect 13097 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13291 45807
rect 13097 45703 13291 45761
rect 13097 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13291 45703
rect 13097 45599 13291 45657
rect 13097 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13291 45599
rect 13097 45495 13291 45553
rect 13097 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13291 45495
rect 13097 45391 13291 45449
rect 13097 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13291 45391
rect 13097 45287 13291 45345
rect 13097 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13291 45287
rect 13097 45183 13291 45241
rect 13097 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13291 45183
rect 13097 45079 13291 45137
rect 13097 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13291 45079
rect 13097 44892 13291 45033
rect 70802 69758 70824 69774
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70802 69700 71000 69758
rect 70802 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70802 69596 71000 69654
rect 70802 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70802 69492 71000 69550
rect 70802 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70802 69388 71000 69446
rect 70802 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70802 69284 71000 69342
rect 70802 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70802 69180 71000 69238
rect 70802 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70802 69076 71000 69134
rect 70802 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70802 68972 71000 69030
rect 70802 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70802 68868 71000 68926
rect 70802 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70802 68764 71000 68822
rect 70802 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70802 68660 71000 68718
rect 70802 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70802 68556 71000 68614
rect 70802 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70802 68452 71000 68510
rect 70802 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70802 68348 71000 68406
rect 70802 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70802 68244 71000 68302
rect 70802 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70802 68140 71000 68198
rect 70802 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70802 68036 71000 68094
rect 70802 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70802 67932 71000 67990
rect 70802 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70802 67828 71000 67886
rect 70802 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70802 67724 71000 67782
rect 70802 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70802 67620 71000 67678
rect 70802 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70802 67516 71000 67574
rect 70802 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70802 67412 71000 67470
rect 70802 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70802 67308 71000 67366
rect 70802 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70802 67204 71000 67262
rect 70802 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70802 67100 71000 67158
rect 70802 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70802 66996 71000 67054
rect 70802 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70802 66892 71000 66950
rect 70802 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70802 66788 71000 66846
rect 70802 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70802 66684 71000 66742
rect 70802 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70802 66580 71000 66638
rect 70802 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70802 66476 71000 66534
rect 70802 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70802 66372 71000 66430
rect 70802 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70802 66268 71000 66326
rect 70802 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70802 66164 71000 66222
rect 70802 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70802 66060 71000 66118
rect 70802 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70802 65956 71000 66014
rect 70802 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70802 65852 71000 65910
rect 70802 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70802 65748 71000 65806
rect 70802 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70802 65644 71000 65702
rect 70802 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70802 65540 71000 65598
rect 70802 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70802 65436 71000 65494
rect 70802 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70802 65332 71000 65390
rect 70802 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70802 65228 71000 65286
rect 70802 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70802 65124 71000 65182
rect 70802 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70802 65020 71000 65078
rect 70802 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70802 64916 71000 64974
rect 70802 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70802 64812 71000 64870
rect 70802 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70802 64708 71000 64766
rect 70802 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70802 64604 71000 64662
rect 70802 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70802 64500 71000 64558
rect 70802 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70802 64396 71000 64454
rect 70802 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70802 64292 71000 64350
rect 70802 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70802 64188 71000 64246
rect 70802 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70802 64084 71000 64142
rect 70802 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70802 63980 71000 64038
rect 70802 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70802 63876 71000 63934
rect 70802 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70802 63772 71000 63830
rect 70802 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70802 63668 71000 63726
rect 70802 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70802 63564 71000 63622
rect 70802 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70802 63460 71000 63518
rect 70802 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70802 63356 71000 63414
rect 70802 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70802 63252 71000 63310
rect 70802 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70802 63148 71000 63206
rect 70802 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70802 63044 71000 63102
rect 70802 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70802 62940 71000 62998
rect 70802 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70802 62836 71000 62894
rect 70802 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70802 62732 71000 62790
rect 70802 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70802 62628 71000 62686
rect 70802 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70802 62524 71000 62582
rect 70802 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70802 62420 71000 62478
rect 70802 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70802 62316 71000 62374
rect 70802 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70802 62212 71000 62270
rect 70802 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70802 62108 71000 62166
rect 70802 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70802 62004 71000 62062
rect 70802 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70802 61900 71000 61958
rect 70802 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70802 61796 71000 61854
rect 70802 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70802 61692 71000 61750
rect 70802 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70802 61588 71000 61646
rect 70802 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70802 61484 71000 61542
rect 70802 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70802 61380 71000 61438
rect 70802 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70802 61276 71000 61334
rect 70802 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70802 61172 71000 61230
rect 70802 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70802 61068 71000 61126
rect 70802 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70802 60964 71000 61022
rect 70802 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70802 60860 71000 60918
rect 70802 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70802 60756 71000 60814
rect 70802 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70802 60652 71000 60710
rect 70802 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70802 60548 71000 60606
rect 70802 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70802 60444 71000 60502
rect 70802 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70802 60340 71000 60398
rect 70802 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70802 60236 71000 60294
rect 70802 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70802 60132 71000 60190
rect 70802 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70802 60028 71000 60086
rect 70802 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70802 59924 71000 59982
rect 70802 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70802 59820 71000 59878
rect 70802 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70802 59716 71000 59774
rect 70802 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70802 59612 71000 59670
rect 70802 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70802 59508 71000 59566
rect 70802 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70802 59404 71000 59462
rect 70802 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70802 59300 71000 59358
rect 70802 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70802 59196 71000 59254
rect 70802 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70802 59092 71000 59150
rect 70802 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70802 58988 71000 59046
rect 70802 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70802 58884 71000 58942
rect 70802 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70802 58780 71000 58838
rect 70802 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70802 58676 71000 58734
rect 70802 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70802 58572 71000 58630
rect 70802 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70802 58468 71000 58526
rect 70802 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70802 58364 71000 58422
rect 70802 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70802 58260 71000 58318
rect 70802 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70802 58156 71000 58214
rect 70802 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70802 58052 71000 58110
rect 70802 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70802 57948 71000 58006
rect 70802 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70802 57844 71000 57902
rect 70802 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70802 57740 71000 57798
rect 70802 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70802 57636 71000 57694
rect 70802 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70802 57532 71000 57590
rect 70802 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70802 57428 71000 57486
rect 70802 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70802 57324 71000 57382
rect 70802 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70802 57220 71000 57278
rect 70802 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70802 57116 71000 57174
rect 70802 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70802 57012 71000 57070
rect 70802 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70802 56908 71000 56966
rect 70802 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70802 56804 71000 56862
rect 70802 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70802 56700 71000 56758
rect 70802 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70802 56596 71000 56654
rect 70802 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70802 56492 71000 56550
rect 70802 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70802 56388 71000 56446
rect 70802 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70802 56284 71000 56342
rect 70802 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70802 56180 71000 56238
rect 70802 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70802 56076 71000 56134
rect 70802 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70802 55972 71000 56030
rect 70802 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70802 55868 71000 55926
rect 70802 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70802 55764 71000 55822
rect 70802 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70802 55660 71000 55718
rect 70802 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70802 55556 71000 55614
rect 70802 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70802 55452 71000 55510
rect 70802 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70802 55348 71000 55406
rect 70802 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70802 55244 71000 55302
rect 70802 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70802 55140 71000 55198
rect 70802 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70802 55036 71000 55094
rect 70802 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70802 54932 71000 54990
rect 70802 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70802 54828 71000 54886
rect 70802 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70802 54724 71000 54782
rect 70802 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70802 54620 71000 54678
rect 70802 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70802 54516 71000 54574
rect 70802 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70802 54412 71000 54470
rect 70802 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70802 54308 71000 54366
rect 70802 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70802 54204 71000 54262
rect 70802 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70802 54100 71000 54158
rect 70802 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70802 53996 71000 54054
rect 70802 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70802 53892 71000 53950
rect 70802 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70802 53788 71000 53846
rect 70802 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70802 53684 71000 53742
rect 70802 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70802 53580 71000 53638
rect 70802 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70802 53476 71000 53534
rect 70802 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70802 53372 71000 53430
rect 70802 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70802 53268 71000 53326
rect 70802 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70802 53164 71000 53222
rect 70802 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70802 53060 71000 53118
rect 70802 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70802 52956 71000 53014
rect 70802 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70802 52852 71000 52910
rect 70802 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70802 52748 71000 52806
rect 70802 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70802 52644 71000 52702
rect 70802 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70802 52540 71000 52598
rect 70802 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70802 52436 71000 52494
rect 70802 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70802 52332 71000 52390
rect 70802 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70802 52228 71000 52286
rect 70802 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70802 52124 71000 52182
rect 70802 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70802 52020 71000 52078
rect 70802 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70802 51916 71000 51974
rect 70802 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70802 51812 71000 51870
rect 70802 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70802 51708 71000 51766
rect 70802 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70802 51604 71000 51662
rect 70802 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70802 51500 71000 51558
rect 70802 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70802 51396 71000 51454
rect 70802 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70802 51292 71000 51350
rect 70802 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70802 51188 71000 51246
rect 70802 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70802 51084 71000 51142
rect 70802 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70802 50980 71000 51038
rect 70802 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70802 50876 71000 50934
rect 70802 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70802 50772 71000 50830
rect 70802 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70802 50668 71000 50726
rect 70802 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70802 50564 71000 50622
rect 70802 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70802 50460 71000 50518
rect 70802 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70802 50356 71000 50414
rect 70802 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70802 50252 71000 50310
rect 70802 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70802 50148 71000 50206
rect 70802 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70802 50044 71000 50102
rect 70802 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70802 49940 71000 49998
rect 70802 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70802 49836 71000 49894
rect 70802 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70802 49732 71000 49790
rect 70802 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70802 49628 71000 49686
rect 70802 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70802 49524 71000 49582
rect 70802 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70802 49420 71000 49478
rect 70802 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70802 49316 71000 49374
rect 70802 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70802 49212 71000 49270
rect 70802 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70802 49108 71000 49166
rect 70802 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70802 49004 71000 49062
rect 70802 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70802 48900 71000 48958
rect 70802 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70802 48796 71000 48854
rect 70802 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70802 48692 71000 48750
rect 70802 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70802 48588 71000 48646
rect 70802 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70802 48484 71000 48542
rect 70802 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70802 48380 71000 48438
rect 70802 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70802 48276 71000 48334
rect 70802 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70802 48172 71000 48230
rect 70802 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70802 48068 71000 48126
rect 70802 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70802 47964 71000 48022
rect 70802 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70802 47860 71000 47918
rect 70802 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70802 47756 71000 47814
rect 70802 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70802 47652 71000 47710
rect 70802 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70802 47548 71000 47606
rect 70802 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70802 47444 71000 47502
rect 70802 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70802 47340 71000 47398
rect 70802 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70802 47236 71000 47294
rect 70802 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70802 47132 71000 47190
rect 70802 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70802 47028 71000 47086
rect 70802 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70802 46924 71000 46982
rect 70802 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70802 46820 71000 46878
rect 70802 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70802 46716 71000 46774
rect 70802 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70802 46612 71000 46670
rect 70802 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70802 46508 71000 46566
rect 70802 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70802 46404 71000 46462
rect 70802 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70802 46300 71000 46358
rect 70802 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70802 46196 71000 46254
rect 70802 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70802 46092 71000 46150
rect 70802 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70802 45988 71000 46046
rect 70802 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70802 45884 71000 45942
rect 70802 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70802 45780 71000 45838
rect 70802 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70802 45676 71000 45734
rect 70802 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70802 45572 71000 45630
rect 70802 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70802 45468 71000 45526
rect 70802 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70802 45364 71000 45422
rect 70802 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70802 45260 71000 45318
rect 70802 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70802 45156 71000 45214
rect 70802 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70802 45052 71000 45110
rect 70802 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70802 44948 71000 45006
tri 13291 44892 13323 44924 sw
rect 70802 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 13097 44847 13323 44892
tri 13323 44847 13368 44892 sw
rect 13097 44844 13368 44847
tri 13097 44831 13110 44844 ne
rect 13110 44831 13368 44844
tri 13110 44785 13155 44831 ne
rect 13155 44824 13368 44831
rect 13155 44785 13254 44824
tri 13155 44740 13201 44785 ne
rect 13201 44778 13254 44785
rect 13300 44802 13368 44824
tri 13368 44802 13413 44847 sw
rect 70802 44844 71000 44902
rect 13300 44786 13413 44802
tri 13413 44786 13429 44802 sw
rect 70802 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
rect 13300 44778 13429 44786
rect 13201 44741 13429 44778
tri 13429 44741 13474 44786 sw
rect 13201 44740 13474 44741
tri 13201 44708 13233 44740 ne
rect 13233 44708 13474 44740
tri 13233 44663 13278 44708 ne
rect 13278 44696 13474 44708
tri 13474 44696 13519 44741 sw
rect 70802 44740 71000 44798
rect 13278 44692 13519 44696
rect 13278 44663 13386 44692
tri 13278 44618 13323 44663 ne
rect 13323 44646 13386 44663
rect 13432 44651 13519 44692
tri 13519 44651 13565 44696 sw
rect 70802 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
rect 13432 44646 13565 44651
rect 13323 44618 13565 44646
tri 13565 44618 13597 44651 sw
rect 70802 44636 71000 44694
tri 13323 44573 13368 44618 ne
rect 13368 44573 13597 44618
tri 13597 44573 13643 44618 sw
rect 70802 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
tri 13368 44527 13413 44573 ne
rect 13413 44560 13643 44573
rect 13413 44527 13518 44560
tri 13413 44482 13459 44527 ne
rect 13459 44514 13518 44527
rect 13564 44527 13643 44560
tri 13643 44527 13688 44573 sw
rect 70802 44532 71000 44590
rect 13564 44514 13688 44527
rect 13459 44482 13688 44514
tri 13688 44482 13733 44527 sw
rect 70802 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
tri 13459 44467 13474 44482 ne
rect 13474 44467 13733 44482
tri 13733 44467 13749 44482 sw
tri 13474 44421 13519 44467 ne
rect 13519 44428 13749 44467
rect 13519 44421 13650 44428
tri 13519 44376 13565 44421 ne
rect 13565 44382 13650 44421
rect 13696 44421 13749 44428
tri 13749 44421 13794 44467 sw
rect 70802 44428 71000 44486
rect 13696 44382 13794 44421
rect 13565 44376 13794 44382
tri 13794 44376 13839 44421 sw
rect 70802 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
tri 13565 44331 13610 44376 ne
rect 13610 44331 13839 44376
tri 13839 44331 13884 44376 sw
tri 13610 44298 13643 44331 ne
rect 13643 44298 13884 44331
tri 13884 44298 13917 44331 sw
rect 70802 44324 71000 44382
tri 13643 44253 13688 44298 ne
rect 13688 44296 13917 44298
rect 13688 44253 13782 44296
tri 13688 44208 13733 44253 ne
rect 13733 44250 13782 44253
rect 13828 44286 13917 44296
tri 13917 44286 13929 44298 sw
rect 13828 44250 13929 44286
rect 13733 44241 13929 44250
tri 13929 44241 13975 44286 sw
rect 70802 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
rect 13733 44208 13975 44241
tri 13733 44163 13778 44208 ne
rect 13778 44195 13975 44208
tri 13975 44195 14020 44241 sw
rect 70802 44220 71000 44278
rect 13778 44164 14020 44195
rect 13778 44163 13914 44164
tri 13778 44159 13781 44163 ne
rect 13781 44159 13914 44163
tri 13781 44114 13827 44159 ne
rect 13827 44118 13914 44159
rect 13960 44159 14020 44164
tri 14020 44159 14056 44195 sw
rect 70802 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
rect 13960 44118 14056 44159
rect 13827 44114 14056 44118
tri 14056 44114 14101 44159 sw
rect 70802 44116 71000 44174
tri 13827 44069 13872 44114 ne
rect 13872 44069 14101 44114
tri 14101 44069 14146 44114 sw
rect 70802 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
tri 13872 44024 13917 44069 ne
rect 13917 44032 14146 44069
rect 13917 44024 14046 44032
tri 13917 44011 13929 44024 ne
rect 13929 44011 14046 44024
tri 13929 43966 13975 44011 ne
rect 13975 43986 14046 44011
rect 14092 44024 14146 44032
tri 14146 44024 14191 44069 sw
rect 14092 44011 14191 44024
tri 14191 44011 14204 44024 sw
rect 70802 44012 71000 44070
rect 14092 43986 14204 44011
rect 13975 43966 14204 43986
tri 14204 43966 14249 44011 sw
rect 70802 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
tri 13975 43921 14020 43966 ne
rect 14020 43921 14249 43966
tri 14249 43921 14294 43966 sw
tri 14020 43876 14065 43921 ne
rect 14065 43900 14294 43921
rect 14065 43876 14178 43900
tri 14065 43840 14101 43876 ne
rect 14101 43854 14178 43876
rect 14224 43876 14294 43900
tri 14294 43876 14339 43921 sw
rect 70802 43908 71000 43966
rect 14224 43854 14339 43876
rect 14101 43840 14339 43854
tri 14339 43840 14375 43876 sw
rect 70802 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
tri 14101 43795 14146 43840 ne
rect 14146 43795 14375 43840
tri 14375 43795 14421 43840 sw
rect 70802 43804 71000 43862
tri 14146 43749 14191 43795 ne
rect 14191 43768 14421 43795
rect 14191 43749 14310 43768
tri 14191 43704 14237 43749 ne
rect 14237 43722 14310 43749
rect 14356 43749 14421 43768
tri 14421 43749 14466 43795 sw
rect 70802 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 14356 43722 14466 43749
rect 14237 43704 14466 43722
tri 14466 43704 14511 43749 sw
tri 14237 43692 14249 43704 ne
rect 14249 43692 14511 43704
tri 14511 43692 14523 43704 sw
rect 70802 43700 71000 43758
tri 14249 43647 14294 43692 ne
rect 14294 43647 14523 43692
tri 14523 43647 14569 43692 sw
rect 70802 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
tri 14294 43601 14339 43647 ne
rect 14339 43636 14569 43647
rect 14339 43601 14442 43636
tri 14339 43556 14385 43601 ne
rect 14385 43590 14442 43601
rect 14488 43601 14569 43636
tri 14569 43601 14614 43647 sw
rect 14488 43590 14614 43601
rect 14385 43556 14614 43590
tri 14614 43556 14659 43601 sw
rect 70802 43596 71000 43654
tri 14385 43520 14421 43556 ne
rect 14421 43520 14659 43556
tri 14659 43520 14695 43556 sw
rect 70802 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
tri 14421 43475 14466 43520 ne
rect 14466 43504 14695 43520
rect 14466 43475 14574 43504
tri 14466 43430 14511 43475 ne
rect 14511 43458 14574 43475
rect 14620 43475 14695 43504
tri 14695 43475 14740 43520 sw
rect 70802 43492 71000 43550
rect 14620 43458 14740 43475
rect 14511 43430 14740 43458
tri 14740 43430 14785 43475 sw
rect 70802 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
tri 14511 43385 14556 43430 ne
rect 14556 43385 14785 43430
tri 14785 43385 14831 43430 sw
rect 70802 43388 71000 43446
tri 14556 43372 14569 43385 ne
rect 14569 43372 14831 43385
tri 14831 43372 14843 43385 sw
tri 14569 43327 14614 43372 ne
rect 14614 43327 14706 43372
tri 14614 43282 14659 43327 ne
rect 14659 43326 14706 43327
rect 14752 43327 14843 43372
tri 14843 43327 14888 43372 sw
rect 70802 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
rect 14752 43326 14888 43327
rect 14659 43282 14888 43326
tri 14888 43282 14933 43327 sw
rect 70802 43284 71000 43342
tri 14659 43237 14704 43282 ne
rect 14704 43240 14933 43282
rect 14704 43237 14838 43240
tri 14704 43201 14740 43237 ne
rect 14740 43201 14838 43237
tri 14740 43155 14785 43201 ne
rect 14785 43194 14838 43201
rect 14884 43237 14933 43240
tri 14933 43237 14979 43282 sw
rect 70802 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 14884 43201 14979 43237
tri 14979 43201 15015 43237 sw
rect 14884 43194 15015 43201
rect 14785 43191 15015 43194
tri 15015 43191 15024 43201 sw
rect 14785 43155 15024 43191
tri 14785 43110 14831 43155 ne
rect 14831 43146 15024 43155
tri 15024 43146 15069 43191 sw
rect 70802 43180 71000 43238
rect 14831 43110 15069 43146
tri 14831 43065 14876 43110 ne
rect 14876 43108 15069 43110
rect 14876 43065 14970 43108
tri 14876 43062 14879 43065 ne
rect 14879 43062 14970 43065
rect 15016 43101 15069 43108
tri 15069 43101 15114 43146 sw
rect 70802 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
rect 15016 43062 15114 43101
tri 15114 43062 15153 43101 sw
rect 70802 43076 71000 43134
tri 14879 43017 14924 43062 ne
rect 14924 43017 15153 43062
tri 15153 43017 15199 43062 sw
rect 70802 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
tri 14924 42971 14969 43017 ne
rect 14969 42976 15199 43017
rect 14969 42971 15102 42976
tri 14969 42926 15015 42971 ne
rect 15015 42930 15102 42971
rect 15148 42971 15199 42976
tri 15199 42971 15244 43017 sw
rect 70802 42972 71000 43030
rect 15148 42930 15244 42971
rect 15015 42926 15244 42930
tri 15244 42926 15289 42971 sw
rect 70802 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
tri 15015 42917 15024 42926 ne
rect 15024 42917 15289 42926
tri 15289 42917 15298 42926 sw
tri 15024 42872 15069 42917 ne
rect 15069 42872 15298 42917
tri 15298 42872 15343 42917 sw
tri 15069 42827 15114 42872 ne
rect 15114 42844 15343 42872
rect 15114 42827 15234 42844
tri 15114 42781 15159 42827 ne
rect 15159 42798 15234 42827
rect 15280 42827 15343 42844
tri 15343 42827 15389 42872 sw
rect 70802 42868 71000 42926
rect 15280 42798 15389 42827
rect 15159 42781 15389 42798
tri 15389 42781 15434 42827 sw
rect 70802 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
tri 15159 42742 15199 42781 ne
rect 15199 42742 15434 42781
tri 15434 42742 15473 42781 sw
rect 70802 42764 71000 42822
tri 15199 42697 15244 42742 ne
rect 15244 42712 15473 42742
rect 15244 42697 15366 42712
tri 15244 42652 15289 42697 ne
rect 15289 42666 15366 42697
rect 15412 42697 15473 42712
tri 15473 42697 15518 42742 sw
rect 70802 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
rect 15412 42666 15518 42697
rect 15289 42652 15518 42666
tri 15518 42652 15563 42697 sw
rect 70802 42660 71000 42718
tri 15289 42607 15334 42652 ne
rect 15334 42607 15563 42652
tri 15563 42607 15609 42652 sw
rect 70802 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
tri 15334 42597 15343 42607 ne
rect 15343 42597 15609 42607
tri 15609 42597 15618 42607 sw
tri 15343 42552 15389 42597 ne
rect 15389 42580 15618 42597
rect 15389 42552 15498 42580
tri 15389 42507 15434 42552 ne
rect 15434 42534 15498 42552
rect 15544 42552 15618 42580
tri 15618 42552 15663 42597 sw
rect 70802 42556 71000 42614
rect 15544 42534 15663 42552
rect 15434 42507 15663 42534
tri 15663 42507 15708 42552 sw
rect 70802 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
tri 15434 42462 15479 42507 ne
rect 15479 42462 15708 42507
tri 15708 42462 15753 42507 sw
tri 15479 42423 15518 42462 ne
rect 15518 42448 15753 42462
rect 15518 42423 15630 42448
tri 15518 42377 15563 42423 ne
rect 15563 42402 15630 42423
rect 15676 42423 15753 42448
tri 15753 42423 15793 42462 sw
rect 70802 42452 71000 42510
rect 15676 42402 15793 42423
rect 15563 42377 15793 42402
tri 15793 42377 15838 42423 sw
rect 70802 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
tri 15563 42332 15609 42377 ne
rect 15609 42332 15838 42377
tri 15838 42332 15883 42377 sw
rect 70802 42348 71000 42406
tri 15609 42287 15654 42332 ne
rect 15654 42316 15883 42332
rect 15654 42287 15762 42316
tri 15654 42278 15663 42287 ne
rect 15663 42278 15762 42287
tri 15663 42233 15708 42278 ne
rect 15708 42270 15762 42278
rect 15808 42287 15883 42316
tri 15883 42287 15928 42332 sw
rect 70802 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 15808 42278 15928 42287
tri 15928 42278 15937 42287 sw
rect 15808 42270 15937 42278
rect 15708 42233 15937 42270
tri 15937 42233 15983 42278 sw
rect 70802 42244 71000 42302
tri 15708 42187 15753 42233 ne
rect 15753 42187 15983 42233
tri 15983 42187 16028 42233 sw
rect 70802 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
tri 15753 42142 15799 42187 ne
rect 15799 42184 16028 42187
rect 15799 42142 15894 42184
tri 15799 42103 15838 42142 ne
rect 15838 42138 15894 42142
rect 15940 42142 16028 42184
tri 16028 42142 16073 42187 sw
rect 15940 42138 16073 42142
rect 15838 42103 16073 42138
tri 16073 42103 16112 42142 sw
rect 70802 42140 71000 42198
tri 15838 42058 15883 42103 ne
rect 15883 42097 16112 42103
tri 16112 42097 16118 42103 sw
rect 15883 42058 16118 42097
tri 15883 42013 15928 42058 ne
rect 15928 42052 16118 42058
tri 16118 42052 16163 42097 sw
rect 70802 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
rect 15928 42013 16026 42052
tri 15928 41967 15973 42013 ne
rect 15973 42006 16026 42013
rect 16072 42007 16163 42052
tri 16163 42007 16209 42052 sw
rect 70802 42036 71000 42094
rect 16072 42006 16209 42007
rect 15973 41967 16209 42006
tri 15973 41964 15977 41967 ne
rect 15977 41964 16209 41967
tri 16209 41964 16251 42007 sw
rect 70802 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
tri 15977 41919 16022 41964 ne
rect 16022 41920 16251 41964
rect 16022 41919 16158 41920
tri 16022 41874 16067 41919 ne
rect 16067 41874 16158 41919
rect 16204 41919 16251 41920
tri 16251 41919 16296 41964 sw
rect 70802 41932 71000 41990
rect 16204 41874 16296 41919
tri 16296 41874 16341 41919 sw
rect 70802 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
tri 16067 41829 16112 41874 ne
rect 16112 41829 16341 41874
tri 16341 41829 16387 41874 sw
tri 16112 41823 16118 41829 ne
rect 16118 41823 16387 41829
tri 16387 41823 16393 41829 sw
rect 70802 41828 71000 41886
tri 16118 41777 16163 41823 ne
rect 16163 41788 16393 41823
rect 16163 41777 16290 41788
tri 16163 41732 16209 41777 ne
rect 16209 41742 16290 41777
rect 16336 41777 16393 41788
tri 16393 41777 16438 41823 sw
rect 70802 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 16336 41742 16438 41777
rect 16209 41732 16438 41742
tri 16438 41732 16483 41777 sw
tri 16209 41687 16254 41732 ne
rect 16254 41687 16483 41732
tri 16483 41687 16528 41732 sw
rect 70802 41724 71000 41782
tri 16254 41645 16296 41687 ne
rect 16296 41656 16528 41687
rect 16296 41645 16422 41656
tri 16296 41599 16341 41645 ne
rect 16341 41610 16422 41645
rect 16468 41645 16528 41656
tri 16528 41645 16571 41687 sw
rect 70802 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
rect 16468 41610 16571 41645
rect 16341 41599 16571 41610
tri 16571 41599 16616 41645 sw
rect 70802 41620 71000 41678
tri 16341 41554 16387 41599 ne
rect 16387 41554 16616 41599
tri 16616 41554 16661 41599 sw
rect 70802 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
tri 16387 41509 16432 41554 ne
rect 16432 41524 16661 41554
rect 16432 41509 16554 41524
tri 16432 41503 16438 41509 ne
rect 16438 41503 16554 41509
tri 16438 41458 16483 41503 ne
rect 16483 41478 16554 41503
rect 16600 41509 16661 41524
tri 16661 41509 16706 41554 sw
rect 70802 41516 71000 41574
rect 16600 41503 16706 41509
tri 16706 41503 16712 41509 sw
rect 16600 41478 16712 41503
rect 16483 41458 16712 41478
tri 16712 41458 16757 41503 sw
rect 70802 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
tri 16483 41413 16528 41458 ne
rect 16528 41413 16757 41458
tri 16757 41413 16803 41458 sw
tri 16528 41367 16573 41413 ne
rect 16573 41392 16803 41413
rect 16573 41367 16686 41392
tri 16573 41325 16616 41367 ne
rect 16616 41346 16686 41367
rect 16732 41367 16803 41392
tri 16803 41367 16848 41413 sw
rect 70802 41412 71000 41470
rect 16732 41346 16848 41367
rect 16616 41325 16848 41346
tri 16848 41325 16890 41367 sw
rect 70802 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
tri 16616 41280 16661 41325 ne
rect 16661 41280 16890 41325
tri 16890 41280 16935 41325 sw
rect 70802 41308 71000 41366
tri 16661 41235 16706 41280 ne
rect 16706 41260 16935 41280
rect 16706 41235 16818 41260
tri 16706 41189 16751 41235 ne
rect 16751 41214 16818 41235
rect 16864 41235 16935 41260
tri 16935 41235 16981 41280 sw
rect 70802 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
rect 16864 41214 16981 41235
rect 16751 41189 16981 41214
tri 16981 41189 17026 41235 sw
rect 70802 41204 71000 41262
tri 16751 41183 16757 41189 ne
rect 16757 41183 17026 41189
tri 17026 41183 17032 41189 sw
tri 16757 41138 16803 41183 ne
rect 16803 41138 17032 41183
tri 17032 41138 17077 41183 sw
rect 70802 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
tri 16803 41093 16848 41138 ne
rect 16848 41128 17077 41138
rect 16848 41093 16950 41128
tri 16848 41048 16893 41093 ne
rect 16893 41082 16950 41093
rect 16996 41093 17077 41128
tri 17077 41093 17122 41138 sw
rect 70802 41100 71000 41158
rect 16996 41082 17122 41093
rect 16893 41048 17122 41082
tri 17122 41048 17167 41093 sw
rect 70802 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
tri 16893 41005 16935 41048 ne
rect 16935 41005 17167 41048
tri 17167 41005 17210 41048 sw
tri 16935 40960 16981 41005 ne
rect 16981 41003 17210 41005
tri 17210 41003 17213 41005 sw
rect 16981 40996 17213 41003
rect 16981 40960 17082 40996
tri 16981 40915 17026 40960 ne
rect 17026 40950 17082 40960
rect 17128 40957 17213 40996
tri 17213 40957 17258 41003 sw
rect 70802 40996 71000 41054
rect 17128 40950 17258 40957
rect 17026 40915 17258 40950
tri 17026 40870 17071 40915 ne
rect 17071 40912 17258 40915
tri 17258 40912 17303 40957 sw
rect 70802 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
rect 17071 40870 17303 40912
tri 17071 40867 17074 40870 ne
rect 17074 40867 17303 40870
tri 17303 40867 17348 40912 sw
rect 70802 40892 71000 40950
tri 17074 40821 17119 40867 ne
rect 17119 40864 17349 40867
rect 17119 40821 17214 40864
tri 17119 40776 17165 40821 ne
rect 17165 40818 17214 40821
rect 17260 40821 17349 40864
tri 17349 40821 17394 40867 sw
rect 70802 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 17260 40818 17394 40821
rect 17165 40776 17394 40818
tri 17394 40776 17439 40821 sw
rect 70802 40788 71000 40846
tri 17165 40731 17210 40776 ne
rect 17210 40732 17439 40776
rect 17210 40731 17346 40732
tri 17210 40728 17213 40731 ne
rect 17213 40728 17346 40731
tri 17213 40683 17258 40728 ne
rect 17258 40686 17346 40728
rect 17392 40731 17439 40732
tri 17439 40731 17484 40776 sw
rect 70802 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
rect 17392 40728 17484 40731
tri 17484 40728 17487 40731 sw
rect 17392 40686 17487 40728
rect 17258 40683 17487 40686
tri 17487 40683 17532 40728 sw
rect 70802 40684 71000 40742
tri 17258 40638 17303 40683 ne
rect 17303 40638 17532 40683
tri 17532 40638 17577 40683 sw
rect 70802 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
tri 17303 40593 17348 40638 ne
rect 17348 40600 17577 40638
rect 17348 40593 17478 40600
tri 17348 40547 17393 40593 ne
rect 17393 40554 17478 40593
rect 17524 40593 17577 40600
tri 17577 40593 17623 40638 sw
rect 17524 40554 17623 40593
rect 17393 40547 17623 40554
tri 17623 40547 17668 40593 sw
rect 70802 40580 71000 40638
tri 17394 40502 17439 40547 ne
rect 17439 40502 17668 40547
tri 17668 40502 17713 40547 sw
rect 70802 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
tri 17439 40457 17484 40502 ne
rect 17484 40468 17713 40502
rect 17484 40457 17610 40468
tri 17484 40411 17529 40457 ne
rect 17529 40422 17610 40457
rect 17656 40457 17713 40468
tri 17713 40457 17759 40502 sw
rect 70802 40476 71000 40534
rect 17656 40422 17759 40457
rect 17529 40411 17759 40422
tri 17759 40411 17804 40457 sw
rect 70802 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
tri 17529 40409 17532 40411 ne
rect 17532 40409 17804 40411
tri 17804 40409 17807 40411 sw
tri 17532 40363 17577 40409 ne
rect 17577 40363 17807 40409
tri 17807 40363 17852 40409 sw
rect 70802 40372 71000 40430
tri 17577 40318 17623 40363 ne
rect 17623 40336 17852 40363
rect 17623 40318 17742 40336
tri 17623 40273 17668 40318 ne
rect 17668 40290 17742 40318
rect 17788 40318 17852 40336
tri 17852 40318 17897 40363 sw
rect 70802 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 17788 40290 17897 40318
rect 17668 40273 17897 40290
tri 17897 40273 17942 40318 sw
tri 17668 40228 17713 40273 ne
rect 17713 40228 17942 40273
tri 17942 40228 17987 40273 sw
rect 70802 40268 71000 40326
rect 17713 40227 17987 40228
tri 17987 40227 17988 40228 sw
tri 17713 40182 17759 40227 ne
rect 17759 40204 17988 40227
rect 17759 40182 17874 40204
tri 17759 40137 17804 40182 ne
rect 17804 40158 17874 40182
rect 17920 40182 17988 40204
tri 17988 40182 18033 40227 sw
rect 70802 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
rect 17920 40158 18033 40182
rect 17804 40137 18033 40158
tri 18033 40137 18078 40182 sw
rect 70802 40164 71000 40222
tri 17804 40092 17849 40137 ne
rect 17849 40092 18078 40137
tri 18078 40092 18123 40137 sw
rect 70802 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
tri 17849 40089 17852 40092 ne
rect 17852 40089 18123 40092
tri 18123 40089 18126 40092 sw
tri 17852 40044 17897 40089 ne
rect 17897 40072 18126 40089
rect 17897 40044 18006 40072
tri 17897 39999 17942 40044 ne
rect 17942 40026 18006 40044
rect 18052 40044 18126 40072
tri 18126 40044 18171 40089 sw
rect 70802 40060 71000 40118
rect 18052 40026 18171 40044
rect 17942 39999 18171 40026
tri 18171 39999 18217 40044 sw
rect 70802 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
tri 17942 39953 17987 39999 ne
rect 17987 39953 18217 39999
tri 18217 39953 18262 39999 sw
rect 70802 39956 71000 40014
tri 17987 39908 18033 39953 ne
rect 18033 39940 18262 39953
rect 18033 39908 18138 39940
tri 18033 39863 18078 39908 ne
rect 18078 39894 18138 39908
rect 18184 39908 18262 39940
tri 18262 39908 18307 39953 sw
rect 70802 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
rect 18184 39894 18307 39908
rect 18078 39863 18307 39894
tri 18307 39863 18353 39908 sw
tri 18078 39817 18123 39863 ne
rect 18123 39817 18353 39863
tri 18353 39817 18398 39863 sw
rect 70802 39852 71000 39910
tri 18123 39772 18169 39817 ne
rect 18169 39808 18398 39817
rect 18169 39772 18270 39808
tri 18169 39769 18171 39772 ne
rect 18171 39769 18270 39772
tri 18171 39724 18217 39769 ne
rect 18217 39762 18270 39769
rect 18316 39772 18398 39808
tri 18398 39772 18443 39817 sw
rect 70802 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 18316 39769 18443 39772
tri 18443 39769 18446 39772 sw
rect 18316 39762 18446 39769
rect 18217 39724 18446 39762
tri 18446 39724 18491 39769 sw
rect 70802 39748 71000 39806
tri 18217 39679 18262 39724 ne
rect 18262 39679 18491 39724
tri 18491 39679 18537 39724 sw
rect 70802 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
tri 18262 39634 18307 39679 ne
rect 18307 39676 18537 39679
rect 18307 39633 18402 39676
tri 18307 39589 18352 39633 ne
rect 18352 39630 18402 39633
rect 18448 39633 18537 39676
tri 18537 39633 18582 39679 sw
rect 70802 39644 71000 39702
rect 18448 39630 18582 39633
rect 18352 39589 18582 39630
tri 18582 39589 18627 39633 sw
rect 70802 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
tri 18352 39543 18397 39589 ne
rect 18397 39544 18627 39589
rect 18397 39543 18534 39544
tri 18397 39498 18443 39543 ne
rect 18443 39498 18534 39543
rect 18580 39543 18627 39544
tri 18627 39543 18672 39589 sw
rect 18580 39498 18672 39543
tri 18672 39498 18717 39543 sw
rect 70802 39540 71000 39598
tri 18443 39453 18488 39498 ne
rect 18488 39453 18717 39498
tri 18717 39453 18762 39498 sw
rect 70802 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
tri 18488 39449 18491 39453 ne
rect 18491 39449 18762 39453
tri 18762 39449 18766 39453 sw
tri 18491 39404 18537 39449 ne
rect 18537 39412 18766 39449
rect 18537 39404 18666 39412
tri 18537 39359 18582 39404 ne
rect 18582 39366 18666 39404
rect 18712 39404 18766 39412
tri 18766 39404 18811 39449 sw
rect 70802 39436 71000 39494
rect 18712 39366 18811 39404
rect 18582 39359 18811 39366
tri 18811 39359 18856 39404 sw
rect 70802 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
tri 18582 39314 18627 39359 ne
rect 18627 39314 18856 39359
tri 18856 39314 18901 39359 sw
rect 70802 39332 71000 39390
tri 18627 39269 18672 39314 ne
rect 18672 39280 18901 39314
rect 18672 39269 18798 39280
tri 18672 39224 18717 39269 ne
rect 18717 39234 18798 39269
rect 18844 39269 18901 39280
tri 18901 39269 18946 39314 sw
rect 70802 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
rect 18844 39234 18946 39269
rect 18717 39224 18946 39234
tri 18946 39224 18991 39269 sw
rect 70802 39228 71000 39286
tri 18717 39179 18762 39224 ne
rect 18762 39179 18991 39224
tri 18991 39179 19037 39224 sw
rect 70802 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
tri 18762 39133 18807 39179 ne
rect 18807 39148 19037 39179
rect 18807 39133 18930 39148
tri 18807 39130 18811 39133 ne
rect 18811 39130 18930 39133
tri 18811 39085 18856 39130 ne
rect 18856 39102 18930 39130
rect 18976 39133 19037 39148
tri 19037 39133 19082 39179 sw
rect 18976 39130 19082 39133
tri 19082 39130 19085 39133 sw
rect 18976 39102 19085 39130
rect 18856 39085 19085 39102
tri 19085 39085 19131 39130 sw
rect 70802 39124 71000 39182
tri 18856 39039 18901 39085 ne
rect 18901 39039 19131 39085
tri 19131 39039 19176 39085 sw
rect 70802 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
tri 18901 38994 18947 39039 ne
rect 18947 39016 19176 39039
rect 18947 38994 19062 39016
tri 18947 38949 18991 38994 ne
rect 18991 38970 19062 38994
rect 19108 38994 19176 39016
tri 19176 38994 19221 39039 sw
rect 70802 39020 71000 39078
rect 19108 38970 19221 38994
rect 18991 38949 19221 38970
tri 19221 38949 19266 38994 sw
rect 70802 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
tri 18991 38904 19037 38949 ne
rect 19037 38904 19266 38949
tri 19266 38904 19311 38949 sw
rect 70802 38916 71000 38974
tri 19037 38859 19082 38904 ne
rect 19082 38884 19311 38904
rect 19082 38859 19194 38884
tri 19082 38814 19127 38859 ne
rect 19127 38838 19194 38859
rect 19240 38859 19311 38884
tri 19311 38859 19356 38904 sw
rect 70802 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 19240 38838 19356 38859
rect 19127 38814 19356 38838
tri 19356 38814 19401 38859 sw
tri 19127 38810 19131 38814 ne
rect 19131 38810 19401 38814
tri 19401 38810 19405 38814 sw
rect 70802 38812 71000 38870
tri 19131 38765 19176 38810 ne
rect 19176 38765 19405 38810
tri 19405 38765 19450 38810 sw
rect 70802 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
tri 19176 38720 19221 38765 ne
rect 19221 38752 19450 38765
rect 19221 38720 19326 38752
tri 19221 38675 19266 38720 ne
rect 19266 38706 19326 38720
rect 19372 38720 19450 38752
tri 19450 38720 19495 38765 sw
rect 19372 38706 19495 38720
rect 19266 38675 19495 38706
tri 19495 38675 19541 38720 sw
rect 70802 38708 71000 38766
tri 19266 38630 19311 38675 ne
rect 19311 38671 19541 38675
tri 19541 38671 19544 38675 sw
rect 19311 38630 19544 38671
tri 19311 38585 19356 38630 ne
rect 19356 38626 19544 38630
tri 19544 38626 19589 38671 sw
rect 70802 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
rect 19356 38620 19589 38626
rect 19356 38585 19458 38620
tri 19356 38539 19401 38585 ne
rect 19401 38574 19458 38585
rect 19504 38581 19589 38620
tri 19589 38581 19634 38626 sw
rect 70802 38604 71000 38662
rect 19504 38574 19634 38581
rect 19401 38539 19634 38574
tri 19401 38536 19405 38539 ne
rect 19405 38536 19634 38539
tri 19634 38536 19679 38581 sw
rect 70802 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
tri 19405 38494 19447 38536 ne
rect 19447 38494 19679 38536
tri 19679 38494 19721 38536 sw
rect 70802 38500 71000 38558
tri 19447 38449 19492 38494 ne
rect 19492 38488 19721 38494
rect 19492 38449 19590 38488
tri 19492 38404 19537 38449 ne
rect 19537 38442 19590 38449
rect 19636 38449 19721 38488
tri 19721 38449 19766 38494 sw
rect 70802 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 19636 38442 19766 38449
rect 19537 38404 19766 38442
tri 19766 38404 19811 38449 sw
tri 19537 38359 19582 38404 ne
rect 19582 38359 19811 38404
tri 19811 38359 19857 38404 sw
rect 70802 38396 71000 38454
tri 19582 38352 19589 38359 ne
rect 19589 38356 19857 38359
rect 19589 38352 19722 38356
tri 19589 38307 19634 38352 ne
rect 19634 38310 19722 38352
rect 19768 38352 19857 38356
tri 19857 38352 19863 38359 sw
rect 19768 38310 19863 38352
rect 19634 38307 19863 38310
tri 19863 38307 19909 38352 sw
rect 70802 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
tri 19634 38261 19679 38307 ne
rect 19679 38261 19909 38307
tri 19909 38261 19954 38307 sw
rect 70802 38292 71000 38350
tri 19679 38216 19725 38261 ne
rect 19725 38224 19954 38261
rect 19725 38216 19854 38224
tri 19725 38175 19766 38216 ne
rect 19766 38178 19854 38216
rect 19900 38216 19954 38224
tri 19954 38216 19999 38261 sw
rect 70802 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
rect 19900 38178 19999 38216
rect 19766 38175 19999 38178
tri 19999 38175 20041 38216 sw
rect 70802 38188 71000 38246
tri 19766 38129 19811 38175 ne
rect 19811 38129 20041 38175
tri 20041 38129 20086 38175 sw
rect 70802 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
tri 19811 38084 19857 38129 ne
rect 19857 38092 20086 38129
rect 19857 38084 19986 38092
tri 19857 38039 19902 38084 ne
rect 19902 38046 19986 38084
rect 20032 38084 20086 38092
tri 20086 38084 20131 38129 sw
rect 70802 38084 71000 38142
rect 20032 38046 20131 38084
rect 19902 38039 20131 38046
tri 20131 38039 20176 38084 sw
tri 19902 38032 19909 38039 ne
rect 19909 38032 20176 38039
tri 20176 38032 20183 38039 sw
rect 70802 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
tri 19909 37987 19954 38032 ne
rect 19954 37987 20183 38032
tri 20183 37987 20228 38032 sw
tri 19954 37942 19999 37987 ne
rect 19999 37960 20228 37987
rect 19999 37942 20118 37960
tri 19999 37897 20044 37942 ne
rect 20044 37914 20118 37942
rect 20164 37942 20228 37960
tri 20228 37942 20273 37987 sw
rect 70802 37980 71000 38038
rect 20164 37914 20273 37942
rect 20044 37897 20273 37914
tri 20273 37897 20319 37942 sw
rect 70802 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
tri 20044 37855 20086 37897 ne
rect 20086 37855 20319 37897
tri 20319 37855 20360 37897 sw
rect 70802 37876 71000 37934
tri 20086 37810 20131 37855 ne
rect 20131 37828 20360 37855
rect 20131 37810 20250 37828
tri 20131 37765 20176 37810 ne
rect 20176 37782 20250 37810
rect 20296 37810 20360 37828
tri 20360 37810 20405 37855 sw
rect 70802 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
rect 20296 37782 20405 37810
rect 20176 37765 20405 37782
tri 20405 37765 20451 37810 sw
rect 70802 37772 71000 37830
tri 20176 37719 20221 37765 ne
rect 20221 37719 20451 37765
tri 20451 37719 20496 37765 sw
rect 70802 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
tri 20221 37713 20228 37719 ne
rect 20228 37713 20496 37719
tri 20496 37713 20503 37719 sw
tri 20228 37667 20273 37713 ne
rect 20273 37696 20503 37713
rect 20273 37667 20382 37696
tri 20273 37622 20319 37667 ne
rect 20319 37650 20382 37667
rect 20428 37667 20503 37696
tri 20503 37667 20548 37713 sw
rect 70802 37668 71000 37726
rect 20428 37650 20548 37667
rect 20319 37622 20548 37650
tri 20548 37622 20593 37667 sw
rect 70802 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
tri 20319 37577 20364 37622 ne
rect 20364 37577 20593 37622
tri 20593 37577 20638 37622 sw
tri 20364 37535 20405 37577 ne
rect 20405 37574 20638 37577
tri 20638 37574 20641 37577 sw
rect 20405 37564 20641 37574
rect 20405 37535 20514 37564
tri 20405 37490 20451 37535 ne
rect 20451 37518 20514 37535
rect 20560 37529 20641 37564
tri 20641 37529 20687 37574 sw
rect 70802 37564 71000 37622
rect 20560 37518 20687 37529
rect 20451 37490 20687 37518
tri 20451 37445 20496 37490 ne
rect 20496 37483 20687 37490
tri 20687 37483 20732 37529 sw
rect 70802 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
rect 20496 37445 20732 37483
tri 20496 37438 20503 37445 ne
rect 20503 37438 20732 37445
tri 20732 37438 20777 37483 sw
rect 70802 37460 71000 37518
tri 20503 37400 20541 37438 ne
rect 20541 37432 20777 37438
rect 20541 37400 20646 37432
tri 20541 37355 20586 37400 ne
rect 20586 37386 20646 37400
rect 20692 37400 20777 37432
tri 20777 37400 20815 37438 sw
rect 70802 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
rect 20692 37386 20815 37400
rect 20586 37355 20815 37386
tri 20815 37355 20861 37400 sw
rect 70802 37356 71000 37414
tri 20586 37309 20631 37355 ne
rect 20631 37309 20861 37355
tri 20861 37309 20906 37355 sw
rect 70802 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
tri 20631 37264 20677 37309 ne
rect 20677 37300 20906 37309
rect 20677 37264 20778 37300
tri 20677 37254 20687 37264 ne
rect 20687 37254 20778 37264
rect 20824 37264 20906 37300
tri 20906 37264 20951 37309 sw
rect 20824 37254 20951 37264
tri 20951 37254 20961 37264 sw
tri 20687 37209 20732 37254 ne
rect 20732 37209 20961 37254
tri 20961 37209 21006 37254 sw
rect 70802 37252 71000 37310
tri 20732 37164 20777 37209 ne
rect 20777 37168 21006 37209
rect 20777 37164 20910 37168
tri 20777 37119 20822 37164 ne
rect 20822 37122 20910 37164
rect 20956 37164 21006 37168
tri 21006 37164 21051 37209 sw
rect 70802 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
rect 20956 37122 21051 37164
rect 20822 37119 21051 37122
tri 21051 37119 21097 37164 sw
rect 70802 37148 71000 37206
tri 20822 37080 20861 37119 ne
rect 20861 37080 21097 37119
tri 21097 37080 21135 37119 sw
rect 70802 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
tri 20861 37035 20906 37080 ne
rect 20906 37036 21135 37080
rect 20906 37035 21042 37036
tri 20906 36990 20951 37035 ne
rect 20951 36990 21042 37035
rect 21088 37035 21135 37036
tri 21135 37035 21180 37080 sw
rect 70802 37044 71000 37102
rect 21088 36990 21180 37035
tri 21180 36990 21225 37035 sw
rect 70802 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
tri 20951 36945 20996 36990 ne
rect 20996 36945 21225 36990
tri 21225 36945 21271 36990 sw
tri 20996 36935 21006 36945 ne
rect 21006 36935 21271 36945
tri 21271 36935 21281 36945 sw
rect 70802 36940 71000 36998
tri 21006 36889 21051 36935 ne
rect 21051 36904 21281 36935
rect 21051 36889 21174 36904
tri 21051 36844 21097 36889 ne
rect 21097 36858 21174 36889
rect 21220 36889 21281 36904
tri 21281 36889 21326 36935 sw
rect 70802 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
rect 21220 36858 21326 36889
rect 21097 36844 21326 36858
tri 21326 36844 21371 36889 sw
tri 21097 36799 21142 36844 ne
rect 21142 36799 21371 36844
tri 21371 36799 21416 36844 sw
rect 70802 36836 71000 36894
tri 21142 36761 21180 36799 ne
rect 21180 36772 21416 36799
rect 21180 36761 21306 36772
tri 21180 36715 21225 36761 ne
rect 21225 36726 21306 36761
rect 21352 36761 21416 36772
tri 21416 36761 21455 36799 sw
rect 70802 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
rect 21352 36726 21455 36761
rect 21225 36715 21455 36726
tri 21455 36715 21500 36761 sw
rect 70802 36732 71000 36790
tri 21225 36670 21271 36715 ne
rect 21271 36670 21500 36715
tri 21500 36670 21545 36715 sw
rect 70802 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
tri 21271 36625 21316 36670 ne
rect 21316 36640 21545 36670
rect 21316 36625 21438 36640
tri 21316 36615 21326 36625 ne
rect 21326 36615 21438 36625
tri 21326 36570 21371 36615 ne
rect 21371 36594 21438 36615
rect 21484 36625 21545 36640
tri 21545 36625 21590 36670 sw
rect 70802 36628 71000 36686
rect 21484 36615 21590 36625
tri 21590 36615 21600 36625 sw
rect 21484 36594 21600 36615
rect 21371 36570 21600 36594
tri 21600 36570 21645 36615 sw
rect 70802 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
tri 21371 36525 21416 36570 ne
rect 21416 36525 21645 36570
tri 21645 36525 21691 36570 sw
tri 21416 36479 21461 36525 ne
rect 21461 36508 21691 36525
rect 21461 36479 21570 36508
tri 21461 36441 21500 36479 ne
rect 21500 36462 21570 36479
rect 21616 36479 21691 36508
tri 21691 36479 21736 36525 sw
rect 70802 36524 71000 36582
rect 21616 36476 21736 36479
tri 21736 36476 21739 36479 sw
rect 70802 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
rect 21616 36462 21739 36476
rect 21500 36441 21739 36462
tri 21500 36396 21545 36441 ne
rect 21545 36431 21739 36441
tri 21739 36431 21784 36476 sw
rect 21545 36396 21784 36431
tri 21545 36351 21590 36396 ne
rect 21590 36386 21784 36396
tri 21784 36386 21829 36431 sw
rect 70802 36420 71000 36478
rect 21590 36376 21829 36386
rect 21590 36351 21702 36376
tri 21590 36341 21600 36351 ne
rect 21600 36341 21702 36351
tri 21600 36305 21635 36341 ne
rect 21635 36330 21702 36341
rect 21748 36341 21829 36376
tri 21829 36341 21875 36386 sw
rect 70802 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 21748 36330 21875 36341
rect 21635 36305 21875 36330
tri 21875 36305 21910 36341 sw
rect 70802 36316 71000 36374
tri 21635 36260 21681 36305 ne
rect 21681 36260 21910 36305
tri 21910 36260 21955 36305 sw
rect 70802 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
tri 21681 36215 21726 36260 ne
rect 21726 36244 21955 36260
rect 21726 36215 21834 36244
tri 21726 36170 21771 36215 ne
rect 21771 36198 21834 36215
rect 21880 36215 21955 36244
tri 21955 36215 22000 36260 sw
rect 21880 36198 22000 36215
rect 21771 36170 22000 36198
tri 22000 36170 22045 36215 sw
rect 70802 36212 71000 36270
tri 21771 36157 21784 36170 ne
rect 21784 36157 22045 36170
tri 22045 36157 22059 36170 sw
rect 70802 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
tri 21784 36111 21829 36157 ne
rect 21829 36112 22059 36157
rect 21829 36111 21966 36112
tri 21829 36066 21875 36111 ne
rect 21875 36066 21966 36111
rect 22012 36111 22059 36112
tri 22059 36111 22104 36157 sw
rect 22012 36066 22104 36111
tri 22104 36066 22149 36111 sw
rect 70802 36108 71000 36166
tri 21875 36021 21920 36066 ne
rect 21920 36021 22149 36066
tri 22149 36021 22194 36066 sw
rect 70802 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
tri 21920 35986 21955 36021 ne
rect 21955 35986 22194 36021
tri 22194 35986 22229 36021 sw
rect 70802 36004 71000 36062
tri 21955 35941 22000 35986 ne
rect 22000 35980 22229 35986
rect 22000 35941 22098 35980
tri 22000 35895 22045 35941 ne
rect 22045 35934 22098 35941
rect 22144 35941 22229 35980
tri 22229 35941 22275 35986 sw
rect 70802 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 22144 35934 22275 35941
rect 22045 35895 22275 35934
tri 22275 35895 22320 35941 sw
rect 70802 35900 71000 35958
tri 22045 35850 22091 35895 ne
rect 22091 35850 22320 35895
tri 22320 35850 22365 35895 sw
rect 70802 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
tri 22091 35837 22104 35850 ne
rect 22104 35848 22365 35850
rect 22104 35837 22230 35848
tri 22104 35792 22149 35837 ne
rect 22149 35802 22230 35837
rect 22276 35837 22365 35848
tri 22365 35837 22378 35850 sw
rect 22276 35802 22378 35837
rect 22149 35792 22378 35802
tri 22378 35792 22423 35837 sw
rect 70802 35796 71000 35854
tri 22149 35747 22194 35792 ne
rect 22194 35747 22423 35792
tri 22423 35747 22469 35792 sw
rect 70802 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
tri 22194 35701 22239 35747 ne
rect 22239 35716 22469 35747
rect 22239 35701 22362 35716
tri 22239 35666 22275 35701 ne
rect 22275 35670 22362 35701
rect 22408 35701 22469 35716
tri 22469 35701 22514 35747 sw
rect 22408 35670 22514 35701
rect 22275 35666 22514 35670
tri 22514 35666 22549 35701 sw
rect 70802 35692 71000 35750
tri 22275 35621 22320 35666 ne
rect 22320 35621 22549 35666
tri 22549 35621 22594 35666 sw
rect 70802 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
tri 22320 35576 22365 35621 ne
rect 22365 35584 22594 35621
rect 22365 35576 22494 35584
tri 22365 35531 22410 35576 ne
rect 22410 35538 22494 35576
rect 22540 35576 22594 35584
tri 22594 35576 22639 35621 sw
rect 70802 35588 71000 35646
rect 22540 35538 22639 35576
rect 22410 35531 22639 35538
tri 22639 35531 22685 35576 sw
rect 70802 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
tri 22410 35517 22423 35531 ne
rect 22423 35517 22685 35531
tri 22685 35517 22698 35531 sw
tri 22423 35472 22469 35517 ne
rect 22469 35472 22698 35517
tri 22698 35472 22743 35517 sw
rect 70802 35484 71000 35542
tri 22469 35427 22514 35472 ne
rect 22514 35452 22743 35472
rect 22514 35427 22626 35452
tri 22514 35382 22559 35427 ne
rect 22559 35406 22626 35427
rect 22672 35427 22743 35452
tri 22743 35427 22788 35472 sw
rect 70802 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 22672 35406 22788 35427
rect 22559 35382 22788 35406
tri 22788 35382 22833 35427 sw
tri 22559 35347 22594 35382 ne
rect 22594 35379 22833 35382
tri 22833 35379 22837 35382 sw
rect 70802 35380 71000 35438
rect 22594 35347 22837 35379
tri 22594 35301 22639 35347 ne
rect 22639 35333 22837 35347
tri 22837 35333 22882 35379 sw
rect 70802 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
rect 22639 35320 22882 35333
rect 22639 35301 22758 35320
tri 22639 35256 22685 35301 ne
rect 22685 35274 22758 35301
rect 22804 35288 22882 35320
tri 22882 35288 22927 35333 sw
rect 22804 35274 22927 35288
rect 22685 35256 22927 35274
tri 22685 35243 22698 35256 ne
rect 22698 35243 22927 35256
tri 22927 35243 22972 35288 sw
rect 70802 35276 71000 35334
tri 22698 35211 22730 35243 ne
rect 22730 35211 22972 35243
tri 22972 35211 23004 35243 sw
rect 70802 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
tri 22730 35166 22775 35211 ne
rect 22775 35188 23004 35211
rect 22775 35166 22890 35188
tri 22775 35121 22820 35166 ne
rect 22820 35142 22890 35166
rect 22936 35166 23004 35188
tri 23004 35166 23049 35211 sw
rect 70802 35172 71000 35230
rect 22936 35142 23049 35166
rect 22820 35121 23049 35142
tri 23049 35121 23095 35166 sw
rect 70802 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
tri 22820 35075 22865 35121 ne
rect 22865 35075 23095 35121
tri 23095 35075 23140 35121 sw
tri 22865 35059 22882 35075 ne
rect 22882 35059 23140 35075
tri 23140 35059 23156 35075 sw
rect 70802 35068 71000 35126
tri 22882 35014 22927 35059 ne
rect 22927 35056 23156 35059
rect 22927 35014 23022 35056
tri 22927 34969 22972 35014 ne
rect 22972 35010 23022 35014
rect 23068 35014 23156 35056
tri 23156 35014 23201 35059 sw
rect 70802 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
rect 23068 35010 23201 35014
rect 22972 34969 23201 35010
tri 23201 34969 23247 35014 sw
tri 22972 34923 23017 34969 ne
rect 23017 34924 23247 34969
rect 23017 34923 23154 34924
tri 23017 34891 23049 34923 ne
rect 23049 34891 23154 34923
tri 23049 34846 23095 34891 ne
rect 23095 34878 23154 34891
rect 23200 34923 23247 34924
tri 23247 34923 23292 34969 sw
rect 70802 34964 71000 35022
rect 23200 34891 23292 34923
tri 23292 34891 23324 34923 sw
rect 70802 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 23200 34878 23324 34891
rect 23095 34846 23324 34878
tri 23324 34846 23369 34891 sw
rect 70802 34860 71000 34918
tri 23095 34801 23140 34846 ne
rect 23140 34801 23369 34846
tri 23369 34801 23414 34846 sw
rect 70802 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
tri 23140 34756 23185 34801 ne
rect 23185 34792 23414 34801
rect 23185 34756 23286 34792
tri 23185 34739 23201 34756 ne
rect 23201 34746 23286 34756
rect 23332 34756 23414 34792
tri 23414 34756 23459 34801 sw
rect 70802 34756 71000 34814
rect 23332 34746 23459 34756
rect 23201 34739 23459 34746
tri 23459 34739 23476 34756 sw
tri 23201 34694 23247 34739 ne
rect 23247 34694 23476 34739
tri 23476 34694 23521 34739 sw
rect 70802 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
tri 23247 34649 23292 34694 ne
rect 23292 34660 23521 34694
rect 23292 34649 23418 34660
tri 23292 34604 23337 34649 ne
rect 23337 34614 23418 34649
rect 23464 34649 23521 34660
tri 23521 34649 23566 34694 sw
rect 70802 34652 71000 34710
rect 23464 34614 23566 34649
rect 23337 34604 23566 34614
tri 23566 34604 23611 34649 sw
rect 70802 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
tri 23337 34572 23369 34604 ne
rect 23369 34572 23611 34604
tri 23611 34572 23643 34604 sw
tri 23369 34527 23414 34572 ne
rect 23414 34528 23643 34572
rect 23414 34527 23550 34528
tri 23414 34481 23459 34527 ne
rect 23459 34482 23550 34527
rect 23596 34527 23643 34528
tri 23643 34527 23689 34572 sw
rect 70802 34548 71000 34606
rect 23596 34482 23689 34527
rect 23459 34481 23689 34482
tri 23689 34481 23734 34527 sw
rect 70802 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
tri 23459 34436 23505 34481 ne
rect 23505 34436 23734 34481
tri 23734 34436 23779 34481 sw
rect 70802 34444 71000 34502
tri 23505 34420 23521 34436 ne
rect 23521 34420 23779 34436
tri 23779 34420 23795 34436 sw
tri 23521 34375 23566 34420 ne
rect 23566 34396 23795 34420
rect 23566 34375 23682 34396
tri 23566 34329 23611 34375 ne
rect 23611 34350 23682 34375
rect 23728 34375 23795 34396
tri 23795 34375 23841 34420 sw
rect 70802 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
rect 23728 34350 23841 34375
rect 23611 34329 23841 34350
tri 23841 34329 23886 34375 sw
rect 70802 34340 71000 34398
tri 23611 34284 23657 34329 ne
rect 23657 34284 23886 34329
tri 23886 34284 23931 34329 sw
rect 70802 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
tri 23657 34252 23689 34284 ne
rect 23689 34281 23931 34284
tri 23931 34281 23934 34284 sw
rect 23689 34264 23934 34281
rect 23689 34252 23814 34264
tri 23689 34207 23734 34252 ne
rect 23734 34218 23814 34252
rect 23860 34236 23934 34264
tri 23934 34236 23979 34281 sw
rect 70802 34236 71000 34294
rect 23860 34218 23979 34236
rect 23734 34207 23979 34218
tri 23734 34162 23779 34207 ne
rect 23779 34191 23979 34207
tri 23979 34191 24025 34236 sw
rect 23779 34162 24025 34191
tri 23779 34145 23795 34162 ne
rect 23795 34145 24025 34162
tri 24025 34145 24070 34191 sw
rect 70802 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
tri 23795 34117 23824 34145 ne
rect 23824 34132 24070 34145
rect 23824 34117 23946 34132
tri 23824 34071 23869 34117 ne
rect 23869 34086 23946 34117
rect 23992 34117 24070 34132
tri 24070 34117 24099 34145 sw
rect 70802 34132 71000 34190
rect 23992 34086 24099 34117
rect 23869 34071 24099 34086
tri 24099 34071 24144 34117 sw
rect 70802 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
tri 23869 34026 23915 34071 ne
rect 23915 34026 24144 34071
tri 24144 34026 24189 34071 sw
rect 70802 34028 71000 34086
tri 23915 33981 23960 34026 ne
rect 23960 34000 24189 34026
rect 23960 33981 24078 34000
tri 23960 33961 23979 33981 ne
rect 23979 33961 24078 33981
tri 23979 33916 24025 33961 ne
rect 24025 33954 24078 33961
rect 24124 33981 24189 34000
tri 24189 33981 24234 34026 sw
rect 70802 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 24124 33961 24234 33981
tri 24234 33961 24254 33981 sw
rect 24124 33954 24254 33961
rect 24025 33916 24254 33954
tri 24254 33916 24299 33961 sw
rect 70802 33924 71000 33982
tri 24025 33871 24070 33916 ne
rect 24070 33871 24299 33916
tri 24299 33871 24344 33916 sw
rect 70802 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
tri 24070 33826 24115 33871 ne
rect 24115 33868 24344 33871
rect 24115 33826 24210 33868
tri 24115 33797 24144 33826 ne
rect 24144 33822 24210 33826
rect 24256 33826 24344 33868
tri 24344 33826 24389 33871 sw
rect 24256 33822 24389 33826
rect 24144 33797 24389 33822
tri 24389 33797 24418 33826 sw
rect 70802 33820 71000 33878
tri 24144 33752 24189 33797 ne
rect 24189 33752 24418 33797
tri 24418 33752 24463 33797 sw
rect 70802 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
tri 24189 33707 24234 33752 ne
rect 24234 33736 24463 33752
rect 24234 33707 24342 33736
tri 24234 33661 24279 33707 ne
rect 24279 33690 24342 33707
rect 24388 33707 24463 33736
tri 24463 33707 24509 33752 sw
rect 70802 33716 71000 33774
rect 24388 33690 24509 33707
rect 24279 33661 24509 33690
tri 24509 33661 24554 33707 sw
rect 70802 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
tri 24279 33642 24299 33661 ne
rect 24299 33642 24554 33661
tri 24554 33642 24573 33661 sw
tri 24299 33597 24344 33642 ne
rect 24344 33604 24573 33642
rect 24344 33597 24474 33604
tri 24344 33551 24389 33597 ne
rect 24389 33558 24474 33597
rect 24520 33597 24573 33604
tri 24573 33597 24619 33642 sw
rect 70802 33612 71000 33670
rect 24520 33558 24619 33597
rect 24389 33551 24619 33558
tri 24619 33551 24664 33597 sw
rect 70802 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
tri 24389 33506 24435 33551 ne
rect 24435 33506 24664 33551
tri 24664 33506 24709 33551 sw
rect 70802 33508 71000 33566
tri 24435 33477 24463 33506 ne
rect 24463 33477 24709 33506
tri 24709 33477 24738 33506 sw
tri 24463 33432 24509 33477 ne
rect 24509 33472 24738 33477
rect 24509 33432 24606 33472
tri 24509 33387 24554 33432 ne
rect 24554 33426 24606 33432
rect 24652 33432 24738 33472
tri 24738 33432 24783 33477 sw
rect 70802 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 24652 33426 24783 33432
rect 24554 33387 24783 33426
tri 24783 33387 24828 33432 sw
rect 70802 33404 71000 33462
tri 24554 33342 24599 33387 ne
rect 24599 33342 24828 33387
tri 24828 33342 24873 33387 sw
rect 70802 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
tri 24599 33322 24619 33342 ne
rect 24619 33340 24873 33342
rect 24619 33322 24738 33340
tri 24619 33277 24664 33322 ne
rect 24664 33294 24738 33322
rect 24784 33322 24873 33340
tri 24873 33322 24893 33342 sw
rect 24784 33294 24893 33322
rect 24664 33277 24893 33294
tri 24893 33277 24938 33322 sw
rect 70802 33300 71000 33358
tri 24664 33232 24709 33277 ne
rect 24709 33232 24938 33277
tri 24938 33232 24983 33277 sw
rect 70802 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
tri 24709 33187 24754 33232 ne
rect 24754 33208 24983 33232
rect 24754 33187 24870 33208
tri 24754 33158 24783 33187 ne
rect 24783 33162 24870 33187
rect 24916 33187 24983 33208
tri 24983 33187 25029 33232 sw
rect 70802 33196 71000 33254
rect 24916 33183 25029 33187
tri 25029 33183 25032 33187 sw
rect 24916 33162 25032 33183
rect 24783 33158 25032 33162
tri 24783 33113 24828 33158 ne
rect 24828 33138 25032 33158
tri 25032 33138 25077 33183 sw
rect 70802 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
rect 24828 33113 25077 33138
tri 24828 33067 24873 33113 ne
rect 24873 33093 25077 33113
tri 25077 33093 25122 33138 sw
rect 24873 33076 25122 33093
rect 24873 33067 25002 33076
tri 24873 33048 24893 33067 ne
rect 24893 33048 25002 33067
tri 24893 33022 24919 33048 ne
rect 24919 33030 25002 33048
rect 25048 33048 25122 33076
tri 25122 33048 25167 33093 sw
rect 70802 33092 71000 33150
rect 25048 33030 25167 33048
rect 24919 33022 25167 33030
tri 25167 33022 25193 33048 sw
rect 70802 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
tri 24919 32977 24964 33022 ne
rect 24964 32977 25193 33022
tri 25193 32977 25238 33022 sw
rect 70802 32988 71000 33046
tri 24964 32932 25009 32977 ne
rect 25009 32944 25238 32977
rect 25009 32932 25134 32944
tri 25009 32887 25054 32932 ne
rect 25054 32898 25134 32932
rect 25180 32932 25238 32944
tri 25238 32932 25283 32977 sw
rect 70802 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 25180 32898 25283 32932
rect 25054 32887 25283 32898
tri 25283 32887 25329 32932 sw
tri 25054 32864 25077 32887 ne
rect 25077 32864 25329 32887
tri 25329 32864 25351 32887 sw
rect 70802 32884 71000 32942
tri 25077 32819 25122 32864 ne
rect 25122 32819 25351 32864
tri 25351 32819 25397 32864 sw
rect 70802 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
tri 25122 32773 25167 32819 ne
rect 25167 32812 25397 32819
rect 25167 32773 25266 32812
tri 25167 32728 25213 32773 ne
rect 25213 32766 25266 32773
rect 25312 32773 25397 32812
tri 25397 32773 25442 32819 sw
rect 70802 32780 71000 32838
rect 25312 32766 25442 32773
rect 25213 32728 25442 32766
tri 25442 32728 25487 32773 sw
rect 70802 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
tri 25213 32703 25238 32728 ne
rect 25238 32703 25487 32728
tri 25487 32703 25513 32728 sw
tri 25238 32657 25283 32703 ne
rect 25283 32680 25513 32703
rect 25283 32657 25398 32680
tri 25283 32612 25329 32657 ne
rect 25329 32634 25398 32657
rect 25444 32657 25513 32680
tri 25513 32657 25558 32703 sw
rect 70802 32676 71000 32734
rect 25444 32634 25558 32657
rect 25329 32612 25558 32634
tri 25558 32612 25603 32657 sw
rect 70802 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
tri 25329 32567 25374 32612 ne
rect 25374 32567 25603 32612
tri 25603 32567 25648 32612 sw
rect 70802 32572 71000 32630
tri 25374 32544 25397 32567 ne
rect 25397 32548 25648 32567
rect 25397 32544 25530 32548
tri 25397 32499 25442 32544 ne
rect 25442 32502 25530 32544
rect 25576 32544 25648 32548
tri 25648 32544 25671 32567 sw
rect 25576 32502 25671 32544
rect 25442 32499 25671 32502
tri 25671 32499 25716 32544 sw
rect 70802 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
tri 25442 32454 25487 32499 ne
rect 25487 32454 25716 32499
tri 25716 32454 25761 32499 sw
rect 70802 32468 71000 32526
tri 25487 32409 25532 32454 ne
rect 25532 32416 25761 32454
rect 25532 32409 25662 32416
tri 25532 32383 25558 32409 ne
rect 25558 32383 25662 32409
tri 25558 32338 25603 32383 ne
rect 25603 32370 25662 32383
rect 25708 32409 25761 32416
tri 25761 32409 25807 32454 sw
rect 70802 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
rect 25708 32383 25807 32409
tri 25807 32383 25832 32409 sw
rect 25708 32370 25832 32383
rect 25603 32338 25832 32370
tri 25832 32338 25877 32383 sw
rect 70802 32364 71000 32422
tri 25603 32293 25648 32338 ne
rect 25648 32293 25877 32338
tri 25877 32293 25923 32338 sw
rect 70802 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
tri 25648 32247 25693 32293 ne
rect 25693 32284 25923 32293
rect 25693 32247 25794 32284
tri 25693 32225 25716 32247 ne
rect 25716 32238 25794 32247
rect 25840 32247 25923 32284
tri 25923 32247 25968 32293 sw
rect 70802 32260 71000 32318
rect 25840 32238 25968 32247
rect 25716 32225 25968 32238
tri 25968 32225 25991 32247 sw
tri 25716 32179 25761 32225 ne
rect 25761 32179 25991 32225
tri 25991 32179 26036 32225 sw
rect 70802 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
tri 25761 32134 25807 32179 ne
rect 25807 32152 26036 32179
rect 25807 32134 25926 32152
tri 25807 32089 25852 32134 ne
rect 25852 32106 25926 32134
rect 25972 32134 26036 32152
tri 26036 32134 26081 32179 sw
rect 70802 32156 71000 32214
rect 25972 32106 26081 32134
rect 25852 32089 26081 32106
tri 26081 32089 26126 32134 sw
rect 70802 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
tri 25852 32063 25877 32089 ne
rect 25877 32086 26126 32089
tri 26126 32086 26129 32089 sw
rect 25877 32063 26129 32086
tri 25877 32018 25923 32063 ne
rect 25923 32041 26129 32063
tri 26129 32041 26175 32086 sw
rect 70802 32052 71000 32110
rect 25923 32020 26175 32041
rect 25923 32018 26058 32020
tri 25923 31973 25968 32018 ne
rect 25968 31974 26058 32018
rect 26104 31995 26175 32020
tri 26175 31995 26220 32041 sw
rect 70802 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 26104 31974 26220 31995
rect 25968 31973 26220 31974
tri 25968 31950 25991 31973 ne
rect 25991 31950 26220 31973
tri 26220 31950 26265 31995 sw
tri 25991 31928 26013 31950 ne
rect 26013 31928 26265 31950
tri 26265 31928 26287 31950 sw
rect 70802 31948 71000 32006
tri 26013 31883 26058 31928 ne
rect 26058 31888 26287 31928
rect 26058 31883 26190 31888
tri 26058 31837 26103 31883 ne
rect 26103 31842 26190 31883
rect 26236 31883 26287 31888
tri 26287 31883 26333 31928 sw
rect 70802 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
rect 26236 31842 26333 31883
rect 26103 31837 26333 31842
tri 26333 31837 26378 31883 sw
rect 70802 31844 71000 31902
tri 26103 31792 26149 31837 ne
rect 26149 31792 26378 31837
tri 26378 31792 26423 31837 sw
rect 70802 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
tri 26149 31766 26175 31792 ne
rect 26175 31766 26423 31792
tri 26423 31766 26449 31792 sw
tri 26175 31721 26220 31766 ne
rect 26220 31756 26449 31766
rect 26220 31721 26322 31756
tri 26220 31676 26265 31721 ne
rect 26265 31710 26322 31721
rect 26368 31721 26449 31756
tri 26449 31721 26494 31766 sw
rect 70802 31740 71000 31798
rect 26368 31710 26494 31721
rect 26265 31676 26494 31710
tri 26494 31676 26539 31721 sw
rect 70802 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
tri 26265 31631 26310 31676 ne
rect 26310 31631 26539 31676
tri 26539 31631 26585 31676 sw
rect 70802 31636 71000 31694
tri 26310 31608 26333 31631 ne
rect 26333 31624 26585 31631
rect 26333 31608 26454 31624
tri 26333 31563 26378 31608 ne
rect 26378 31578 26454 31608
rect 26500 31608 26585 31624
tri 26585 31608 26607 31631 sw
rect 26500 31578 26607 31608
rect 26378 31563 26607 31578
tri 26607 31563 26652 31608 sw
rect 70802 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
tri 26378 31518 26423 31563 ne
rect 26423 31518 26652 31563
tri 26652 31518 26697 31563 sw
rect 70802 31532 71000 31590
tri 26423 31473 26468 31518 ne
rect 26468 31492 26697 31518
rect 26468 31473 26586 31492
tri 26468 31447 26494 31473 ne
rect 26494 31447 26586 31473
tri 26494 31401 26539 31447 ne
rect 26539 31446 26586 31447
rect 26632 31473 26697 31492
tri 26697 31473 26743 31518 sw
rect 70802 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 26632 31447 26743 31473
tri 26743 31447 26769 31473 sw
rect 26632 31446 26769 31447
rect 26539 31401 26769 31446
tri 26769 31401 26814 31447 sw
rect 70802 31428 71000 31486
tri 26539 31356 26585 31401 ne
rect 26585 31360 26814 31401
rect 26585 31356 26718 31360
tri 26585 31311 26630 31356 ne
rect 26630 31314 26718 31356
rect 26764 31356 26814 31360
tri 26814 31356 26859 31401 sw
rect 70802 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
rect 26764 31314 26859 31356
rect 26630 31311 26859 31314
tri 26859 31311 26904 31356 sw
rect 70802 31324 71000 31382
tri 26630 31289 26652 31311 ne
rect 26652 31289 26904 31311
tri 26904 31289 26927 31311 sw
tri 26652 31243 26697 31289 ne
rect 26697 31243 26927 31289
tri 26927 31243 26972 31289 sw
rect 70802 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
tri 26697 31198 26743 31243 ne
rect 26743 31228 26972 31243
rect 26743 31198 26850 31228
tri 26743 31153 26788 31198 ne
rect 26788 31182 26850 31198
rect 26896 31198 26972 31228
tri 26972 31198 27017 31243 sw
rect 70802 31220 71000 31278
rect 26896 31182 27017 31198
rect 26788 31153 27017 31182
tri 27017 31153 27062 31198 sw
rect 70802 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
tri 26788 31127 26814 31153 ne
rect 26814 31127 27062 31153
tri 27062 31127 27088 31153 sw
tri 26814 31082 26859 31127 ne
rect 26859 31096 27088 31127
rect 26859 31082 26982 31096
tri 26859 31037 26904 31082 ne
rect 26904 31050 26982 31082
rect 27028 31082 27088 31096
tri 27088 31082 27133 31127 sw
rect 70802 31116 71000 31174
rect 27028 31050 27133 31082
rect 26904 31037 27133 31050
tri 27133 31037 27179 31082 sw
rect 70802 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
tri 26904 30991 26949 31037 ne
rect 26949 30991 27179 31037
tri 27179 30991 27224 31037 sw
rect 70802 31012 71000 31070
tri 26949 30969 26972 30991 ne
rect 26972 30988 27224 30991
tri 27224 30988 27227 30991 sw
rect 26972 30969 27227 30988
tri 26972 30924 27017 30969 ne
rect 27017 30964 27227 30969
rect 27017 30924 27114 30964
tri 27017 30879 27062 30924 ne
rect 27062 30918 27114 30924
rect 27160 30943 27227 30964
tri 27227 30943 27272 30988 sw
rect 70802 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
rect 27160 30918 27272 30943
rect 27062 30898 27272 30918
tri 27272 30898 27317 30943 sw
rect 70802 30908 71000 30966
rect 27062 30879 27317 30898
tri 27062 30853 27088 30879 ne
rect 27088 30853 27317 30879
tri 27317 30853 27363 30898 sw
rect 70802 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
tri 27088 30833 27107 30853 ne
rect 27107 30833 27363 30853
tri 27363 30833 27382 30853 sw
tri 27107 30788 27153 30833 ne
rect 27153 30832 27382 30833
rect 27153 30788 27246 30832
tri 27153 30743 27198 30788 ne
rect 27198 30786 27246 30788
rect 27292 30788 27382 30832
tri 27382 30788 27427 30833 sw
rect 70802 30804 71000 30862
rect 27292 30786 27427 30788
rect 27198 30743 27427 30786
tri 27427 30743 27472 30788 sw
rect 70802 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
tri 27198 30698 27243 30743 ne
rect 27243 30700 27472 30743
rect 27243 30698 27378 30700
tri 27243 30669 27272 30698 ne
rect 27272 30669 27378 30698
tri 27272 30623 27317 30669 ne
rect 27317 30654 27378 30669
rect 27424 30698 27472 30700
tri 27472 30698 27517 30743 sw
rect 70802 30700 71000 30758
rect 27424 30669 27517 30698
tri 27517 30669 27547 30698 sw
rect 27424 30654 27547 30669
rect 27317 30623 27547 30654
tri 27547 30623 27592 30669 sw
rect 70802 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
tri 27317 30578 27363 30623 ne
rect 27363 30578 27592 30623
tri 27592 30578 27637 30623 sw
rect 70802 30596 71000 30654
tri 27363 30533 27408 30578 ne
rect 27408 30568 27637 30578
rect 27408 30533 27510 30568
tri 27408 30514 27427 30533 ne
rect 27427 30522 27510 30533
rect 27556 30533 27637 30568
tri 27637 30533 27682 30578 sw
rect 70802 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 27556 30522 27682 30533
rect 27427 30514 27682 30522
tri 27682 30514 27701 30533 sw
tri 27427 30469 27472 30514 ne
rect 27472 30469 27701 30514
tri 27701 30469 27747 30514 sw
rect 70802 30492 71000 30550
tri 27472 30423 27517 30469 ne
rect 27517 30436 27747 30469
rect 27517 30423 27642 30436
tri 27517 30378 27563 30423 ne
rect 27563 30390 27642 30423
rect 27688 30423 27747 30436
tri 27747 30423 27792 30469 sw
rect 70802 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
rect 27688 30390 27792 30423
rect 27563 30378 27792 30390
tri 27792 30378 27837 30423 sw
rect 70802 30388 71000 30446
tri 27563 30349 27592 30378 ne
rect 27592 30349 27837 30378
tri 27837 30349 27866 30378 sw
tri 27592 30304 27637 30349 ne
rect 27637 30304 27866 30349
tri 27866 30304 27911 30349 sw
rect 70802 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
tri 27637 30259 27682 30304 ne
rect 27682 30259 27774 30304
tri 27682 30213 27727 30259 ne
rect 27727 30258 27774 30259
rect 27820 30259 27911 30304
tri 27911 30259 27957 30304 sw
rect 70802 30284 71000 30342
rect 27820 30258 27957 30259
rect 27727 30213 27957 30258
tri 27957 30213 28002 30259 sw
rect 70802 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
tri 27727 30194 27747 30213 ne
rect 27747 30194 28002 30213
tri 28002 30194 28021 30213 sw
tri 27747 30149 27792 30194 ne
rect 27792 30172 28021 30194
rect 27792 30149 27906 30172
tri 27792 30104 27837 30149 ne
rect 27837 30126 27906 30149
rect 27952 30149 28021 30172
tri 28021 30149 28066 30194 sw
rect 70802 30180 71000 30238
rect 27952 30126 28066 30149
rect 27837 30104 28066 30126
tri 28066 30104 28111 30149 sw
rect 70802 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
tri 27837 30059 27882 30104 ne
rect 27882 30059 28111 30104
tri 28111 30059 28157 30104 sw
rect 70802 30076 71000 30134
tri 27882 30029 27911 30059 ne
rect 27911 30040 28157 30059
rect 27911 30029 28038 30040
tri 27911 29984 27957 30029 ne
rect 27957 29994 28038 30029
rect 28084 30029 28157 30040
tri 28157 30029 28186 30059 sw
rect 70802 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 28084 29994 28186 30029
rect 27957 29984 28186 29994
tri 28186 29984 28231 30029 sw
tri 27957 29939 28002 29984 ne
rect 28002 29939 28231 29984
tri 28231 29939 28276 29984 sw
rect 70802 29972 71000 30030
tri 28002 29894 28047 29939 ne
rect 28047 29908 28276 29939
rect 28047 29894 28170 29908
tri 28047 29875 28066 29894 ne
rect 28066 29875 28170 29894
tri 28066 29829 28111 29875 ne
rect 28111 29862 28170 29875
rect 28216 29894 28276 29908
tri 28276 29894 28321 29939 sw
rect 70802 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
rect 28216 29891 28321 29894
tri 28321 29891 28325 29894 sw
rect 28216 29862 28325 29891
rect 28111 29845 28325 29862
tri 28325 29845 28370 29891 sw
rect 70802 29868 71000 29926
rect 28111 29829 28370 29845
tri 28111 29784 28157 29829 ne
rect 28157 29800 28370 29829
tri 28370 29800 28415 29845 sw
rect 70802 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
rect 28157 29784 28415 29800
tri 28157 29755 28186 29784 ne
rect 28186 29776 28415 29784
rect 28186 29755 28302 29776
tri 28186 29739 28202 29755 ne
rect 28202 29739 28302 29755
tri 28202 29694 28247 29739 ne
rect 28247 29730 28302 29739
rect 28348 29755 28415 29776
tri 28415 29755 28460 29800 sw
rect 70802 29764 71000 29822
rect 28348 29739 28460 29755
tri 28460 29739 28476 29755 sw
rect 28348 29730 28476 29739
rect 28247 29694 28476 29730
tri 28476 29694 28521 29739 sw
rect 70802 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
tri 28247 29649 28292 29694 ne
rect 28292 29649 28521 29694
tri 28521 29649 28567 29694 sw
rect 70802 29660 71000 29718
tri 28292 29603 28337 29649 ne
rect 28337 29644 28567 29649
rect 28337 29603 28434 29644
tri 28337 29571 28370 29603 ne
rect 28370 29598 28434 29603
rect 28480 29603 28567 29644
tri 28567 29603 28612 29649 sw
rect 70802 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
rect 28480 29598 28612 29603
rect 28370 29571 28612 29598
tri 28612 29571 28644 29603 sw
tri 28370 29526 28415 29571 ne
rect 28415 29526 28644 29571
tri 28644 29526 28689 29571 sw
rect 70802 29556 71000 29614
tri 28415 29481 28460 29526 ne
rect 28460 29512 28689 29526
rect 28460 29481 28566 29512
tri 28460 29435 28505 29481 ne
rect 28505 29466 28566 29481
rect 28612 29481 28689 29512
tri 28689 29481 28735 29526 sw
rect 70802 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 28612 29466 28735 29481
rect 28505 29435 28735 29466
tri 28735 29435 28780 29481 sw
rect 70802 29452 71000 29510
tri 28505 29419 28521 29435 ne
rect 28521 29419 28780 29435
tri 28780 29419 28796 29435 sw
tri 28521 29374 28567 29419 ne
rect 28567 29380 28796 29419
rect 28567 29374 28698 29380
tri 28567 29329 28612 29374 ne
rect 28612 29334 28698 29374
rect 28744 29374 28796 29380
tri 28796 29374 28841 29419 sw
rect 70802 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
rect 28744 29334 28841 29374
rect 28612 29329 28841 29334
tri 28841 29329 28886 29374 sw
rect 70802 29348 71000 29406
tri 28612 29284 28657 29329 ne
rect 28657 29284 28886 29329
tri 28886 29284 28931 29329 sw
rect 70802 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
tri 28657 29251 28689 29284 ne
rect 28689 29251 28931 29284
tri 28931 29251 28964 29284 sw
tri 28689 29206 28735 29251 ne
rect 28735 29248 28964 29251
rect 28735 29206 28830 29248
tri 28735 29161 28780 29206 ne
rect 28780 29202 28830 29206
rect 28876 29206 28964 29248
tri 28964 29206 29009 29251 sw
rect 70802 29244 71000 29302
rect 28876 29202 29009 29206
rect 28780 29161 29009 29202
tri 29009 29161 29054 29206 sw
rect 70802 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
tri 28780 29116 28825 29161 ne
rect 28825 29116 29054 29161
tri 29054 29116 29099 29161 sw
rect 70802 29140 71000 29198
tri 28825 29100 28841 29116 ne
rect 28841 29100 28962 29116
tri 28841 29055 28886 29100 ne
rect 28886 29070 28962 29100
rect 29008 29100 29099 29116
tri 29099 29100 29115 29116 sw
rect 29008 29070 29115 29100
rect 28886 29055 29115 29070
tri 29115 29055 29161 29100 sw
rect 70802 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
tri 28886 29009 28931 29055 ne
rect 28931 29009 29161 29055
tri 29161 29009 29206 29055 sw
rect 70802 29036 71000 29094
tri 28931 28964 28977 29009 ne
rect 28977 28984 29206 29009
rect 28977 28964 29094 28984
tri 28977 28932 29009 28964 ne
rect 29009 28938 29094 28964
rect 29140 28964 29206 28984
tri 29206 28964 29251 29009 sw
rect 70802 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
rect 29140 28938 29251 28964
rect 29009 28932 29251 28938
tri 29251 28932 29283 28964 sw
rect 70802 28932 71000 28990
tri 29009 28887 29054 28932 ne
rect 29054 28887 29283 28932
tri 29283 28887 29329 28932 sw
tri 29054 28841 29099 28887 ne
rect 29099 28852 29329 28887
rect 29099 28841 29226 28852
tri 29099 28796 29145 28841 ne
rect 29145 28806 29226 28841
rect 29272 28841 29329 28852
tri 29329 28841 29374 28887 sw
rect 70802 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
rect 29272 28806 29374 28841
rect 29145 28796 29374 28806
tri 29374 28796 29419 28841 sw
rect 70802 28828 71000 28886
tri 29145 28780 29161 28796 ne
rect 29161 28793 29419 28796
tri 29419 28793 29422 28796 sw
rect 29161 28780 29422 28793
tri 29161 28735 29206 28780 ne
rect 29206 28748 29422 28780
tri 29422 28748 29467 28793 sw
rect 70802 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
rect 29206 28735 29467 28748
tri 29206 28690 29251 28735 ne
rect 29251 28720 29467 28735
rect 29251 28690 29358 28720
tri 29251 28657 29283 28690 ne
rect 29283 28674 29358 28690
rect 29404 28703 29467 28720
tri 29467 28703 29513 28748 sw
rect 70802 28724 71000 28782
rect 29404 28674 29513 28703
rect 29283 28657 29513 28674
tri 29513 28657 29558 28703 sw
rect 70802 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
tri 29283 28645 29296 28657 ne
rect 29296 28645 29558 28657
tri 29558 28645 29571 28657 sw
tri 29296 28599 29341 28645 ne
rect 29341 28599 29571 28645
tri 29571 28599 29616 28645 sw
rect 70802 28620 71000 28678
tri 29341 28554 29387 28599 ne
rect 29387 28588 29616 28599
rect 29387 28554 29490 28588
tri 29387 28509 29432 28554 ne
rect 29432 28542 29490 28554
rect 29536 28554 29616 28588
tri 29616 28554 29661 28599 sw
rect 70802 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 29536 28542 29661 28554
rect 29432 28509 29661 28542
tri 29661 28509 29706 28554 sw
rect 70802 28516 71000 28574
tri 29432 28473 29467 28509 ne
rect 29467 28473 29706 28509
tri 29706 28473 29742 28509 sw
tri 29467 28428 29513 28473 ne
rect 29513 28456 29742 28473
rect 29513 28428 29622 28456
tri 29513 28383 29558 28428 ne
rect 29558 28410 29622 28428
rect 29668 28428 29742 28456
tri 29742 28428 29787 28473 sw
rect 70802 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
rect 29668 28410 29787 28428
rect 29558 28383 29787 28410
tri 29787 28383 29832 28428 sw
rect 70802 28412 71000 28470
tri 29558 28338 29603 28383 ne
rect 29603 28338 29832 28383
tri 29832 28338 29877 28383 sw
rect 70802 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
tri 29603 28325 29616 28338 ne
rect 29616 28325 29877 28338
tri 29877 28325 29890 28338 sw
tri 29616 28280 29661 28325 ne
rect 29661 28324 29890 28325
rect 29661 28280 29754 28324
tri 29661 28235 29706 28280 ne
rect 29706 28278 29754 28280
rect 29800 28280 29890 28324
tri 29890 28280 29935 28325 sw
rect 70802 28308 71000 28366
rect 29800 28278 29935 28280
rect 29706 28235 29935 28278
tri 29935 28235 29981 28280 sw
rect 70802 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
tri 29706 28189 29751 28235 ne
rect 29751 28192 29981 28235
rect 29751 28189 29886 28192
tri 29751 28154 29787 28189 ne
rect 29787 28154 29886 28189
tri 29787 28109 29832 28154 ne
rect 29832 28146 29886 28154
rect 29932 28189 29981 28192
tri 29981 28189 30026 28235 sw
rect 70802 28204 71000 28262
rect 29932 28154 30026 28189
tri 30026 28154 30061 28189 sw
rect 70802 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
rect 29932 28146 30061 28154
rect 29832 28109 30061 28146
tri 30061 28109 30107 28154 sw
tri 29832 28063 29877 28109 ne
rect 29877 28063 30107 28109
tri 30107 28063 30152 28109 sw
rect 70802 28100 71000 28158
tri 29877 28018 29923 28063 ne
rect 29923 28060 30152 28063
rect 29923 28018 30018 28060
tri 29923 28005 29935 28018 ne
rect 29935 28014 30018 28018
rect 30064 28018 30152 28060
tri 30152 28018 30197 28063 sw
rect 70802 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 30064 28014 30197 28018
rect 29935 28005 30197 28014
tri 30197 28005 30210 28018 sw
tri 29935 27960 29981 28005 ne
rect 29981 27960 30210 28005
tri 30210 27960 30255 28005 sw
rect 70802 27996 71000 28054
tri 29981 27915 30026 27960 ne
rect 30026 27928 30255 27960
rect 30026 27915 30150 27928
tri 30026 27870 30071 27915 ne
rect 30071 27882 30150 27915
rect 30196 27915 30255 27928
tri 30255 27915 30300 27960 sw
rect 70802 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
rect 30196 27882 30300 27915
rect 30071 27870 30300 27882
tri 30300 27870 30345 27915 sw
rect 70802 27892 71000 27950
tri 30071 27834 30107 27870 ne
rect 30107 27834 30345 27870
tri 30345 27834 30381 27870 sw
rect 70802 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
tri 30107 27789 30152 27834 ne
rect 30152 27796 30381 27834
rect 30152 27789 30282 27796
tri 30152 27744 30197 27789 ne
rect 30197 27750 30282 27789
rect 30328 27789 30381 27796
tri 30381 27789 30426 27834 sw
rect 30328 27750 30426 27789
rect 30197 27744 30426 27750
tri 30426 27744 30471 27789 sw
rect 70802 27788 71000 27846
tri 30197 27699 30242 27744 ne
rect 30242 27699 30471 27744
tri 30471 27699 30517 27744 sw
rect 70802 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
tri 30242 27686 30255 27699 ne
rect 30255 27695 30517 27699
tri 30517 27695 30520 27699 sw
rect 30255 27686 30520 27695
tri 30255 27641 30300 27686 ne
rect 30300 27664 30520 27686
rect 30300 27641 30414 27664
tri 30300 27595 30345 27641 ne
rect 30345 27618 30414 27641
rect 30460 27650 30520 27664
tri 30520 27650 30565 27695 sw
rect 70802 27684 71000 27742
rect 30460 27618 30565 27650
rect 30345 27605 30565 27618
tri 30565 27605 30610 27650 sw
rect 70802 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 30345 27595 30610 27605
tri 30345 27560 30381 27595 ne
rect 30381 27560 30610 27595
tri 30610 27560 30655 27605 sw
rect 70802 27580 71000 27638
tri 30381 27550 30391 27560 ne
rect 30391 27550 30655 27560
tri 30655 27550 30665 27560 sw
tri 30391 27505 30436 27550 ne
rect 30436 27532 30665 27550
rect 30436 27505 30546 27532
tri 30436 27460 30481 27505 ne
rect 30481 27486 30546 27505
rect 30592 27505 30665 27532
tri 30665 27505 30710 27550 sw
rect 70802 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
rect 30592 27486 30710 27505
rect 30481 27460 30710 27486
tri 30710 27460 30755 27505 sw
rect 70802 27476 71000 27534
tri 30481 27415 30526 27460 ne
rect 30526 27415 30755 27460
tri 30755 27415 30801 27460 sw
rect 70802 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
tri 30526 27376 30565 27415 ne
rect 30565 27400 30801 27415
rect 30565 27376 30678 27400
tri 30565 27331 30610 27376 ne
rect 30610 27354 30678 27376
rect 30724 27376 30801 27400
tri 30801 27376 30839 27415 sw
rect 30724 27354 30839 27376
rect 30610 27331 30839 27354
tri 30839 27331 30885 27376 sw
rect 70802 27372 71000 27430
tri 30610 27285 30655 27331 ne
rect 30655 27285 30885 27331
tri 30885 27285 30930 27331 sw
rect 70802 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
tri 30655 27240 30701 27285 ne
rect 30701 27268 30930 27285
rect 30701 27240 30810 27268
tri 30701 27231 30710 27240 ne
rect 30710 27231 30810 27240
tri 30710 27185 30755 27231 ne
rect 30755 27222 30810 27231
rect 30856 27240 30930 27268
tri 30930 27240 30975 27285 sw
rect 70802 27268 71000 27326
rect 30856 27231 30975 27240
tri 30975 27231 30985 27240 sw
rect 30856 27222 30985 27231
rect 30755 27185 30985 27222
tri 30985 27185 31030 27231 sw
rect 70802 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
tri 30755 27140 30801 27185 ne
rect 30801 27140 31030 27185
tri 31030 27140 31075 27185 sw
rect 70802 27164 71000 27222
tri 30801 27095 30846 27140 ne
rect 30846 27136 31075 27140
rect 30846 27095 30942 27136
tri 30846 27056 30885 27095 ne
rect 30885 27090 30942 27095
rect 30988 27095 31075 27136
tri 31075 27095 31120 27140 sw
rect 70802 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
rect 30988 27090 31120 27095
rect 30885 27056 31120 27090
tri 31120 27056 31159 27095 sw
rect 70802 27060 71000 27118
tri 30885 27011 30930 27056 ne
rect 30930 27011 31159 27056
tri 31159 27011 31204 27056 sw
rect 70802 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
tri 30930 26966 30975 27011 ne
rect 30975 27004 31204 27011
rect 30975 26966 31074 27004
tri 30975 26921 31020 26966 ne
rect 31020 26958 31074 26966
rect 31120 26966 31204 27004
tri 31204 26966 31249 27011 sw
rect 31120 26958 31249 26966
rect 31020 26921 31249 26958
tri 31249 26921 31295 26966 sw
rect 70802 26956 71000 27014
tri 31020 26911 31030 26921 ne
rect 31030 26911 31295 26921
tri 31295 26911 31304 26921 sw
tri 31030 26866 31075 26911 ne
rect 31075 26872 31304 26911
rect 31075 26866 31206 26872
tri 31075 26821 31120 26866 ne
rect 31120 26826 31206 26866
rect 31252 26866 31304 26872
tri 31304 26866 31349 26911 sw
rect 70802 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
rect 31252 26826 31349 26866
rect 31120 26821 31349 26826
tri 31349 26821 31395 26866 sw
rect 70802 26852 71000 26910
tri 31120 26775 31165 26821 ne
rect 31165 26775 31395 26821
tri 31395 26775 31440 26821 sw
rect 70802 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
tri 31165 26737 31204 26775 ne
rect 31204 26740 31440 26775
rect 31204 26737 31338 26740
tri 31204 26691 31249 26737 ne
rect 31249 26694 31338 26737
rect 31384 26737 31440 26740
tri 31440 26737 31479 26775 sw
rect 70802 26748 71000 26806
rect 31384 26694 31479 26737
rect 31249 26691 31479 26694
tri 31479 26691 31524 26737 sw
rect 70802 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
tri 31249 26646 31295 26691 ne
rect 31295 26646 31524 26691
tri 31524 26646 31569 26691 sw
tri 31295 26601 31340 26646 ne
rect 31340 26608 31569 26646
rect 31340 26601 31470 26608
tri 31340 26591 31349 26601 ne
rect 31349 26591 31470 26601
tri 31349 26546 31395 26591 ne
rect 31395 26562 31470 26591
rect 31516 26601 31569 26608
tri 31569 26601 31614 26646 sw
rect 70802 26644 71000 26702
rect 31516 26598 31614 26601
tri 31614 26598 31617 26601 sw
rect 70802 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
rect 31516 26562 31617 26598
rect 31395 26553 31617 26562
tri 31617 26553 31663 26598 sw
rect 31395 26546 31663 26553
tri 31395 26501 31440 26546 ne
rect 31440 26507 31663 26546
tri 31663 26507 31708 26553 sw
rect 70802 26540 71000 26598
rect 31440 26501 31708 26507
tri 31440 26462 31479 26501 ne
rect 31479 26476 31708 26501
rect 31479 26462 31602 26476
tri 31479 26456 31485 26462 ne
rect 31485 26456 31602 26462
tri 31485 26411 31530 26456 ne
rect 31530 26430 31602 26456
rect 31648 26462 31708 26476
tri 31708 26462 31753 26507 sw
rect 70802 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
rect 31648 26456 31753 26462
tri 31753 26456 31759 26462 sw
rect 31648 26430 31759 26456
rect 31530 26411 31759 26430
tri 31759 26411 31805 26456 sw
rect 70802 26436 71000 26494
tri 31530 26365 31575 26411 ne
rect 31575 26365 31805 26411
tri 31805 26365 31850 26411 sw
rect 70802 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
tri 31575 26320 31621 26365 ne
rect 31621 26344 31850 26365
rect 31621 26320 31734 26344
tri 31621 26278 31663 26320 ne
rect 31663 26298 31734 26320
rect 31780 26320 31850 26344
tri 31850 26320 31895 26365 sw
rect 70802 26332 71000 26390
rect 31780 26298 31895 26320
rect 31663 26278 31895 26298
tri 31895 26278 31937 26320 sw
rect 70802 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
tri 31663 26233 31708 26278 ne
rect 31708 26233 31937 26278
tri 31937 26233 31982 26278 sw
tri 31708 26188 31753 26233 ne
rect 31753 26212 31982 26233
rect 31753 26188 31866 26212
tri 31753 26143 31798 26188 ne
rect 31798 26166 31866 26188
rect 31912 26188 31982 26212
tri 31982 26188 32027 26233 sw
rect 70802 26228 71000 26286
rect 31912 26166 32027 26188
rect 31798 26143 32027 26166
tri 32027 26143 32073 26188 sw
rect 70802 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
tri 31798 26136 31805 26143 ne
rect 31805 26136 32073 26143
tri 32073 26136 32079 26143 sw
tri 31805 26091 31850 26136 ne
rect 31850 26091 32079 26136
tri 32079 26091 32124 26136 sw
rect 70802 26124 71000 26182
tri 31850 26046 31895 26091 ne
rect 31895 26080 32124 26091
rect 31895 26046 31998 26080
tri 31895 26001 31940 26046 ne
rect 31940 26034 31998 26046
rect 32044 26046 32124 26080
tri 32124 26046 32169 26091 sw
rect 70802 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 32044 26034 32169 26046
rect 31940 26001 32169 26034
tri 32169 26001 32215 26046 sw
rect 70802 26020 71000 26078
tri 31940 25959 31982 26001 ne
rect 31982 25959 32215 26001
tri 32215 25959 32257 26001 sw
rect 70802 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
tri 31982 25913 32027 25959 ne
rect 32027 25948 32257 25959
rect 32027 25913 32130 25948
tri 32027 25868 32073 25913 ne
rect 32073 25902 32130 25913
rect 32176 25913 32257 25948
tri 32257 25913 32302 25959 sw
rect 70802 25916 71000 25974
rect 32176 25902 32302 25913
rect 32073 25868 32302 25902
tri 32302 25868 32347 25913 sw
rect 70802 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
tri 32073 25823 32118 25868 ne
rect 32118 25823 32347 25868
tri 32347 25823 32392 25868 sw
tri 32118 25817 32124 25823 ne
rect 32124 25817 32392 25823
tri 32392 25817 32399 25823 sw
tri 32124 25771 32169 25817 ne
rect 32169 25816 32399 25817
rect 32169 25771 32262 25816
tri 32169 25726 32215 25771 ne
rect 32215 25770 32262 25771
rect 32308 25771 32399 25816
tri 32399 25771 32444 25817 sw
rect 70802 25812 71000 25870
rect 32308 25770 32444 25771
rect 32215 25726 32444 25770
tri 32444 25726 32489 25771 sw
rect 70802 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
tri 32215 25681 32260 25726 ne
rect 32260 25684 32489 25726
rect 32260 25681 32394 25684
tri 32260 25639 32302 25681 ne
rect 32302 25639 32394 25681
tri 32302 25594 32347 25639 ne
rect 32347 25638 32394 25639
rect 32440 25681 32489 25684
tri 32489 25681 32534 25726 sw
rect 70802 25708 71000 25766
rect 32440 25639 32534 25681
tri 32534 25639 32576 25681 sw
rect 70802 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 32440 25638 32576 25639
rect 32347 25594 32576 25638
tri 32576 25594 32621 25639 sw
rect 70802 25604 71000 25662
tri 32347 25549 32392 25594 ne
rect 32392 25552 32621 25594
rect 32392 25549 32526 25552
tri 32392 25503 32437 25549 ne
rect 32437 25506 32526 25549
rect 32572 25549 32621 25552
tri 32621 25549 32667 25594 sw
rect 70802 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
rect 32572 25506 32667 25549
rect 32437 25503 32667 25506
tri 32667 25503 32712 25549 sw
tri 32437 25497 32444 25503 ne
rect 32444 25500 32712 25503
tri 32712 25500 32715 25503 sw
rect 70802 25500 71000 25558
rect 32444 25497 32715 25500
tri 32444 25452 32489 25497 ne
rect 32489 25455 32715 25497
tri 32715 25455 32760 25500 sw
rect 32489 25452 32760 25455
tri 32489 25407 32534 25452 ne
rect 32534 25420 32760 25452
rect 32534 25407 32658 25420
tri 32534 25365 32576 25407 ne
rect 32576 25374 32658 25407
rect 32704 25410 32760 25420
tri 32760 25410 32805 25455 sw
rect 70802 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
rect 32704 25374 32805 25410
rect 32576 25365 32805 25374
tri 32805 25365 32851 25410 sw
rect 70802 25396 71000 25454
tri 32576 25361 32579 25365 ne
rect 32579 25361 32851 25365
tri 32851 25361 32854 25365 sw
tri 32579 25316 32625 25361 ne
rect 32625 25316 32854 25361
tri 32854 25316 32899 25361 sw
rect 70802 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
tri 32625 25271 32670 25316 ne
rect 32670 25288 32899 25316
rect 32670 25271 32790 25288
tri 32670 25226 32715 25271 ne
rect 32715 25242 32790 25271
rect 32836 25271 32899 25288
tri 32899 25271 32944 25316 sw
rect 70802 25292 71000 25350
rect 32836 25242 32944 25271
rect 32715 25226 32944 25242
tri 32944 25226 32989 25271 sw
rect 70802 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
tri 32715 25181 32760 25226 ne
rect 32760 25181 32989 25226
tri 32989 25181 33035 25226 sw
rect 70802 25188 71000 25246
tri 32760 25135 32805 25181 ne
rect 32805 25156 33035 25181
rect 32805 25135 32922 25156
tri 32805 25090 32851 25135 ne
rect 32851 25110 32922 25135
rect 32968 25135 33035 25156
tri 33035 25135 33080 25181 sw
rect 70802 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
rect 32968 25110 33080 25135
rect 32851 25090 33080 25110
tri 33080 25090 33125 25135 sw
tri 32851 25045 32896 25090 ne
rect 32896 25045 33125 25090
tri 33125 25045 33170 25090 sw
rect 70802 25084 71000 25142
tri 32896 25042 32899 25045 ne
rect 32899 25042 33170 25045
tri 33170 25042 33173 25045 sw
tri 32899 24997 32944 25042 ne
rect 32944 25024 33173 25042
rect 32944 24997 33054 25024
tri 32944 24951 32989 24997 ne
rect 32989 24978 33054 24997
rect 33100 24997 33173 25024
tri 33173 24997 33219 25042 sw
rect 70802 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
rect 33100 24978 33219 24997
rect 32989 24951 33219 24978
tri 33219 24951 33264 24997 sw
rect 70802 24980 71000 25038
tri 32989 24906 33035 24951 ne
rect 33035 24906 33264 24951
tri 33264 24906 33309 24951 sw
rect 70802 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
tri 33035 24861 33080 24906 ne
rect 33080 24892 33309 24906
rect 33080 24861 33186 24892
tri 33080 24816 33125 24861 ne
rect 33125 24846 33186 24861
rect 33232 24861 33309 24892
tri 33309 24861 33354 24906 sw
rect 70802 24876 71000 24934
rect 33232 24846 33354 24861
rect 33125 24816 33354 24846
tri 33354 24816 33399 24861 sw
rect 70802 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
tri 33125 24771 33170 24816 ne
rect 33170 24771 33399 24816
tri 33399 24771 33445 24816 sw
rect 70802 24772 71000 24830
tri 33170 24725 33215 24771 ne
rect 33215 24760 33445 24771
rect 33215 24725 33318 24760
tri 33215 24722 33219 24725 ne
rect 33219 24722 33318 24725
tri 33219 24677 33264 24722 ne
rect 33264 24714 33318 24722
rect 33364 24725 33445 24760
tri 33445 24725 33490 24771 sw
rect 70802 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
rect 33364 24722 33490 24725
tri 33490 24722 33493 24725 sw
rect 33364 24714 33493 24722
rect 33264 24677 33493 24714
tri 33493 24677 33538 24722 sw
tri 33264 24632 33309 24677 ne
rect 33309 24632 33538 24677
tri 33538 24632 33583 24677 sw
rect 70802 24668 71000 24726
tri 33309 24587 33354 24632 ne
rect 33354 24628 33583 24632
rect 33354 24587 33450 24628
tri 33354 24541 33399 24587 ne
rect 33399 24582 33450 24587
rect 33496 24587 33583 24628
tri 33583 24587 33629 24632 sw
rect 70802 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 33496 24582 33629 24587
rect 33399 24541 33629 24582
tri 33629 24541 33674 24587 sw
rect 70802 24564 71000 24622
tri 33399 24496 33445 24541 ne
rect 33445 24496 33674 24541
tri 33674 24496 33719 24541 sw
rect 70802 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
tri 33445 24451 33490 24496 ne
rect 33490 24451 33582 24496
tri 33490 24406 33535 24451 ne
rect 33535 24450 33582 24451
rect 33628 24451 33719 24496
tri 33719 24451 33764 24496 sw
rect 70802 24460 71000 24518
rect 33628 24450 33764 24451
rect 33535 24406 33764 24450
tri 33764 24406 33809 24451 sw
rect 70802 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
tri 33535 24403 33538 24406 ne
rect 33538 24403 33809 24406
tri 33809 24403 33813 24406 sw
tri 33538 24357 33583 24403 ne
rect 33583 24364 33813 24403
rect 33583 24357 33714 24364
tri 33583 24312 33629 24357 ne
rect 33629 24318 33714 24357
rect 33760 24357 33813 24364
tri 33813 24357 33858 24403 sw
rect 33760 24318 33858 24357
rect 33629 24312 33858 24318
tri 33858 24312 33903 24357 sw
rect 70802 24356 71000 24414
tri 33629 24267 33674 24312 ne
rect 33674 24267 33903 24312
tri 33903 24267 33948 24312 sw
rect 70802 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
tri 33674 24222 33719 24267 ne
rect 33719 24232 33948 24267
rect 33719 24222 33846 24232
tri 33719 24177 33764 24222 ne
rect 33764 24186 33846 24222
rect 33892 24222 33948 24232
tri 33948 24222 33993 24267 sw
rect 70802 24252 71000 24310
rect 33892 24186 33993 24222
rect 33764 24177 33993 24186
tri 33993 24177 34039 24222 sw
rect 70802 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
tri 33764 24131 33809 24177 ne
rect 33809 24131 34039 24177
tri 34039 24131 34084 24177 sw
rect 70802 24148 71000 24206
tri 33809 24128 33813 24131 ne
rect 33813 24128 34084 24131
tri 34084 24128 34087 24131 sw
tri 33813 24083 33858 24128 ne
rect 33858 24100 34087 24128
rect 33858 24083 33978 24100
tri 33858 24038 33903 24083 ne
rect 33903 24054 33978 24083
rect 34024 24083 34087 24100
tri 34087 24083 34132 24128 sw
rect 70802 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
rect 34024 24054 34132 24083
rect 33903 24038 34132 24054
tri 34132 24038 34177 24083 sw
rect 70802 24044 71000 24102
tri 33903 23993 33948 24038 ne
rect 33948 23993 34177 24038
tri 34177 23993 34223 24038 sw
rect 70802 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
tri 33948 23947 33993 23993 ne
rect 33993 23968 34223 23993
rect 33993 23947 34110 23968
tri 33993 23902 34039 23947 ne
rect 34039 23922 34110 23947
rect 34156 23947 34223 23968
tri 34223 23947 34268 23993 sw
rect 34156 23922 34268 23947
rect 34039 23902 34268 23922
tri 34268 23902 34313 23947 sw
rect 70802 23940 71000 23998
tri 34039 23857 34084 23902 ne
rect 34084 23857 34313 23902
tri 34313 23857 34358 23902 sw
rect 70802 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
tri 34084 23812 34129 23857 ne
rect 34129 23836 34358 23857
rect 34129 23812 34242 23836
tri 34129 23809 34132 23812 ne
rect 34132 23809 34242 23812
tri 34132 23763 34177 23809 ne
rect 34177 23790 34242 23809
rect 34288 23812 34358 23836
tri 34358 23812 34403 23857 sw
rect 70802 23836 71000 23894
rect 34288 23809 34403 23812
tri 34403 23809 34407 23812 sw
rect 34288 23790 34407 23809
rect 34177 23763 34407 23790
tri 34407 23763 34452 23809 sw
rect 70802 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
tri 34177 23718 34223 23763 ne
rect 34223 23718 34452 23763
tri 34452 23718 34497 23763 sw
rect 70802 23732 71000 23790
tri 34223 23673 34268 23718 ne
rect 34268 23704 34497 23718
rect 34268 23673 34374 23704
tri 34268 23628 34313 23673 ne
rect 34313 23658 34374 23673
rect 34420 23673 34497 23704
tri 34497 23673 34542 23718 sw
rect 70802 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 34420 23658 34542 23673
rect 34313 23628 34542 23658
tri 34542 23628 34587 23673 sw
rect 70802 23628 71000 23686
tri 34313 23583 34358 23628 ne
rect 34358 23583 34587 23628
tri 34587 23583 34633 23628 sw
tri 34358 23537 34403 23583 ne
rect 34403 23572 34633 23583
rect 34403 23537 34506 23572
tri 34403 23492 34449 23537 ne
rect 34449 23526 34506 23537
rect 34552 23537 34633 23572
tri 34633 23537 34678 23583 sw
rect 70802 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
rect 34552 23526 34678 23537
rect 34449 23492 34678 23526
tri 34678 23492 34723 23537 sw
rect 70802 23524 71000 23582
tri 34449 23489 34452 23492 ne
rect 34452 23489 34723 23492
tri 34723 23489 34726 23492 sw
tri 34452 23444 34497 23489 ne
rect 34497 23444 34726 23489
tri 34726 23444 34771 23489 sw
rect 70802 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
tri 34497 23399 34542 23444 ne
rect 34542 23440 34771 23444
rect 34542 23399 34638 23440
tri 34542 23353 34587 23399 ne
rect 34587 23394 34638 23399
rect 34684 23399 34771 23440
tri 34771 23399 34817 23444 sw
rect 70802 23420 71000 23478
rect 34684 23394 34817 23399
rect 34587 23353 34817 23394
tri 34817 23353 34862 23399 sw
rect 70802 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
tri 34587 23308 34633 23353 ne
rect 34633 23308 34862 23353
tri 34862 23308 34907 23353 sw
rect 70802 23316 71000 23374
tri 34633 23263 34678 23308 ne
rect 34678 23263 34770 23308
tri 34678 23218 34723 23263 ne
rect 34723 23262 34770 23263
rect 34816 23263 34907 23308
tri 34907 23263 34952 23308 sw
rect 70802 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
rect 34816 23262 34952 23263
rect 34723 23218 34952 23262
tri 34952 23218 34997 23263 sw
tri 34723 23173 34768 23218 ne
rect 34768 23176 34997 23218
rect 34768 23173 34902 23176
tri 34768 23169 34771 23173 ne
rect 34771 23169 34902 23173
tri 34771 23124 34817 23169 ne
rect 34817 23130 34902 23169
rect 34948 23173 34997 23176
tri 34997 23173 35043 23218 sw
rect 70802 23212 71000 23270
rect 34948 23169 35043 23173
tri 35043 23169 35046 23173 sw
rect 34948 23130 35046 23169
rect 34817 23127 35046 23130
tri 35046 23127 35088 23169 sw
rect 70802 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
rect 34817 23124 35088 23127
tri 34817 23079 34862 23124 ne
rect 34862 23082 35088 23124
tri 35088 23082 35133 23127 sw
rect 70802 23108 71000 23166
rect 34862 23079 35133 23082
tri 34862 23034 34907 23079 ne
rect 34907 23044 35133 23079
rect 34907 23034 35034 23044
tri 34907 23031 34910 23034 ne
rect 34910 23031 35034 23034
tri 34910 22985 34955 23031 ne
rect 34955 22998 35034 23031
rect 35080 23037 35133 23044
tri 35133 23037 35178 23082 sw
rect 70802 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
rect 35080 23031 35178 23037
tri 35178 23031 35185 23037 sw
rect 35080 22998 35185 23031
rect 34955 22985 35185 22998
tri 35185 22985 35230 23031 sw
rect 70802 23004 71000 23062
tri 34955 22940 35001 22985 ne
rect 35001 22940 35230 22985
tri 35230 22940 35275 22985 sw
rect 70802 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
tri 35001 22895 35046 22940 ne
rect 35046 22912 35275 22940
rect 35046 22895 35166 22912
tri 35046 22853 35088 22895 ne
rect 35088 22866 35166 22895
rect 35212 22895 35275 22912
tri 35275 22895 35320 22940 sw
rect 70802 22900 71000 22958
rect 35212 22866 35320 22895
rect 35088 22853 35320 22866
tri 35320 22853 35362 22895 sw
rect 70802 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
tri 35088 22808 35133 22853 ne
rect 35133 22808 35362 22853
tri 35362 22808 35407 22853 sw
tri 35133 22763 35178 22808 ne
rect 35178 22780 35407 22808
rect 35178 22763 35298 22780
tri 35178 22717 35223 22763 ne
rect 35223 22734 35298 22763
rect 35344 22763 35407 22780
tri 35407 22763 35453 22808 sw
rect 70802 22796 71000 22854
rect 35344 22734 35453 22763
rect 35223 22717 35453 22734
tri 35453 22717 35498 22763 sw
rect 70802 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
tri 35223 22711 35230 22717 ne
rect 35230 22711 35498 22717
tri 35498 22711 35504 22717 sw
tri 35230 22666 35275 22711 ne
rect 35275 22666 35504 22711
tri 35504 22666 35549 22711 sw
rect 70802 22692 71000 22750
tri 35275 22621 35320 22666 ne
rect 35320 22648 35549 22666
rect 35320 22621 35430 22648
tri 35320 22575 35365 22621 ne
rect 35365 22602 35430 22621
rect 35476 22621 35549 22648
tri 35549 22621 35595 22666 sw
rect 70802 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 35476 22602 35595 22621
rect 35365 22575 35595 22602
tri 35595 22575 35640 22621 sw
rect 70802 22588 71000 22646
tri 35365 22533 35407 22575 ne
rect 35407 22533 35640 22575
tri 35640 22533 35682 22575 sw
rect 70802 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
tri 35407 22488 35453 22533 ne
rect 35453 22516 35682 22533
rect 35453 22488 35562 22516
tri 35453 22443 35498 22488 ne
rect 35498 22470 35562 22488
rect 35608 22488 35682 22516
tri 35682 22488 35727 22533 sw
rect 35608 22470 35727 22488
rect 35498 22443 35727 22470
tri 35727 22443 35772 22488 sw
rect 70802 22484 71000 22542
tri 35498 22398 35543 22443 ne
rect 35543 22398 35772 22443
tri 35772 22398 35817 22443 sw
rect 70802 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
tri 35543 22391 35549 22398 ne
rect 35549 22391 35817 22398
tri 35817 22391 35824 22398 sw
tri 35549 22346 35595 22391 ne
rect 35595 22384 35824 22391
rect 35595 22346 35694 22384
tri 35595 22301 35640 22346 ne
rect 35640 22338 35694 22346
rect 35740 22346 35824 22384
tri 35824 22346 35869 22391 sw
rect 70802 22380 71000 22438
rect 35740 22338 35869 22346
rect 35640 22301 35869 22338
tri 35869 22301 35914 22346 sw
rect 70802 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
tri 35640 22256 35685 22301 ne
rect 35685 22256 35914 22301
tri 35914 22256 35959 22301 sw
rect 70802 22276 71000 22334
tri 35685 22214 35727 22256 ne
rect 35727 22252 35959 22256
rect 35727 22214 35826 22252
tri 35727 22169 35772 22214 ne
rect 35772 22206 35826 22214
rect 35872 22214 35959 22252
tri 35959 22214 36001 22256 sw
rect 70802 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 35872 22206 36001 22214
rect 35772 22169 36001 22206
tri 36001 22169 36047 22214 sw
rect 70802 22172 71000 22230
tri 35772 22123 35817 22169 ne
rect 35817 22123 36047 22169
tri 36047 22123 36092 22169 sw
rect 70802 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
tri 35817 22078 35863 22123 ne
rect 35863 22120 36092 22123
rect 35863 22078 35958 22120
tri 35863 22072 35869 22078 ne
rect 35869 22074 35958 22078
rect 36004 22078 36092 22120
tri 36092 22078 36137 22123 sw
rect 36004 22074 36137 22078
rect 35869 22072 36137 22074
tri 36137 22072 36143 22078 sw
tri 35869 22027 35914 22072 ne
rect 35914 22033 36143 22072
tri 36143 22033 36182 22072 sw
rect 70802 22068 71000 22126
rect 35914 22027 36182 22033
tri 35914 21981 35959 22027 ne
rect 35959 21988 36182 22027
tri 36182 21988 36227 22033 sw
rect 70802 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
rect 35959 21981 36090 21988
tri 35959 21936 36005 21981 ne
rect 36005 21942 36090 21981
rect 36136 21943 36227 21988
tri 36227 21943 36273 21988 sw
rect 70802 21964 71000 22022
rect 36136 21942 36273 21943
rect 36005 21936 36273 21942
tri 36005 21933 36008 21936 ne
rect 36008 21933 36273 21936
tri 36273 21933 36282 21943 sw
tri 36008 21888 36053 21933 ne
rect 36053 21888 36282 21933
tri 36282 21888 36327 21933 sw
rect 70802 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
tri 36053 21843 36098 21888 ne
rect 36098 21856 36327 21888
rect 36098 21843 36222 21856
tri 36098 21797 36143 21843 ne
rect 36143 21810 36222 21843
rect 36268 21843 36327 21856
tri 36327 21843 36373 21888 sw
rect 70802 21860 71000 21918
rect 36268 21810 36373 21843
rect 36143 21797 36373 21810
tri 36373 21797 36418 21843 sw
rect 70802 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
tri 36143 21759 36182 21797 ne
rect 36182 21759 36418 21797
tri 36418 21759 36457 21797 sw
tri 36182 21713 36227 21759 ne
rect 36227 21724 36457 21759
rect 36227 21713 36354 21724
tri 36227 21668 36273 21713 ne
rect 36273 21678 36354 21713
rect 36400 21713 36457 21724
tri 36457 21713 36502 21759 sw
rect 70802 21756 71000 21814
rect 36400 21678 36502 21713
rect 36273 21668 36502 21678
tri 36502 21668 36547 21713 sw
rect 70802 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
tri 36273 21623 36318 21668 ne
rect 36318 21623 36547 21668
tri 36547 21623 36592 21668 sw
rect 70802 21652 71000 21710
tri 36318 21613 36327 21623 ne
rect 36327 21613 36592 21623
tri 36592 21613 36602 21623 sw
tri 36327 21568 36373 21613 ne
rect 36373 21592 36602 21613
rect 36373 21568 36486 21592
tri 36373 21523 36418 21568 ne
rect 36418 21546 36486 21568
rect 36532 21568 36602 21592
tri 36602 21568 36647 21613 sw
rect 70802 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
rect 36532 21546 36647 21568
rect 36418 21523 36647 21546
tri 36647 21523 36692 21568 sw
rect 70802 21548 71000 21606
tri 36418 21478 36463 21523 ne
rect 36463 21478 36692 21523
tri 36692 21478 36737 21523 sw
rect 70802 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
tri 36463 21439 36502 21478 ne
rect 36502 21460 36737 21478
rect 36502 21439 36618 21460
tri 36502 21394 36547 21439 ne
rect 36547 21414 36618 21439
rect 36664 21439 36737 21460
tri 36737 21439 36776 21478 sw
rect 70802 21444 71000 21502
rect 36664 21414 36776 21439
rect 36547 21394 36776 21414
tri 36776 21394 36821 21439 sw
rect 70802 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
tri 36547 21349 36592 21394 ne
rect 36592 21349 36821 21394
tri 36821 21349 36867 21394 sw
tri 36592 21303 36637 21349 ne
rect 36637 21328 36867 21349
rect 36637 21303 36750 21328
tri 36637 21294 36647 21303 ne
rect 36647 21294 36750 21303
tri 36647 21249 36692 21294 ne
rect 36692 21282 36750 21294
rect 36796 21303 36867 21328
tri 36867 21303 36912 21349 sw
rect 70802 21340 71000 21398
rect 36796 21294 36912 21303
tri 36912 21294 36921 21303 sw
rect 70802 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 36796 21282 36921 21294
rect 36692 21249 36921 21282
tri 36921 21249 36967 21294 sw
tri 36692 21203 36737 21249 ne
rect 36737 21203 36967 21249
tri 36967 21203 37012 21249 sw
rect 70802 21236 71000 21294
tri 36737 21158 36783 21203 ne
rect 36783 21196 37012 21203
rect 36783 21158 36882 21196
tri 36783 21119 36821 21158 ne
rect 36821 21150 36882 21158
rect 36928 21158 37012 21196
tri 37012 21158 37057 21203 sw
rect 70802 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 36928 21150 37057 21158
rect 36821 21119 37057 21150
tri 37057 21119 37096 21158 sw
rect 70802 21132 71000 21190
tri 36821 21074 36867 21119 ne
rect 36867 21074 37096 21119
tri 37096 21074 37141 21119 sw
rect 70802 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
tri 36867 21029 36912 21074 ne
rect 36912 21064 37141 21074
rect 36912 21029 37014 21064
tri 36912 20984 36957 21029 ne
rect 36957 21018 37014 21029
rect 37060 21029 37141 21064
tri 37141 21029 37186 21074 sw
rect 37060 21018 37186 21029
rect 36957 20984 37186 21018
tri 37186 20984 37231 21029 sw
rect 70802 21028 71000 21086
tri 36957 20974 36967 20984 ne
rect 36967 20974 37231 20984
tri 37231 20974 37241 20984 sw
rect 70802 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
tri 36967 20929 37012 20974 ne
rect 37012 20939 37241 20974
tri 37241 20939 37277 20974 sw
rect 37012 20932 37277 20939
rect 37012 20929 37146 20932
tri 37012 20884 37057 20929 ne
rect 37057 20886 37146 20929
rect 37192 20893 37277 20932
tri 37277 20893 37322 20939 sw
rect 70802 20924 71000 20982
rect 37192 20886 37322 20893
rect 37057 20884 37322 20886
tri 37057 20839 37102 20884 ne
rect 37102 20848 37322 20884
tri 37322 20848 37367 20893 sw
rect 70802 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
rect 37102 20839 37367 20848
tri 37102 20835 37105 20839 ne
rect 37105 20835 37367 20839
tri 37367 20835 37380 20848 sw
tri 37105 20790 37151 20835 ne
rect 37151 20800 37380 20835
rect 37151 20790 37278 20800
tri 37151 20745 37196 20790 ne
rect 37196 20754 37278 20790
rect 37324 20790 37380 20800
tri 37380 20790 37425 20835 sw
rect 70802 20820 71000 20878
rect 37324 20754 37425 20790
rect 37196 20745 37425 20754
tri 37425 20745 37470 20790 sw
rect 70802 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
tri 37196 20700 37241 20745 ne
rect 37241 20700 37470 20745
tri 37470 20700 37515 20745 sw
rect 70802 20716 71000 20774
tri 37241 20664 37277 20700 ne
rect 37277 20668 37515 20700
rect 37277 20664 37410 20668
tri 37277 20619 37322 20664 ne
rect 37322 20622 37410 20664
rect 37456 20664 37515 20668
tri 37515 20664 37551 20700 sw
rect 70802 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
rect 37456 20622 37551 20664
rect 37322 20619 37551 20622
tri 37551 20619 37596 20664 sw
tri 37322 20574 37367 20619 ne
rect 37367 20574 37596 20619
tri 37596 20574 37641 20619 sw
rect 70802 20612 71000 20670
tri 37367 20529 37412 20574 ne
rect 37412 20536 37641 20574
rect 37412 20529 37542 20536
tri 37412 20516 37425 20529 ne
rect 37425 20516 37542 20529
tri 37425 20471 37470 20516 ne
rect 37470 20490 37542 20516
rect 37588 20529 37641 20536
tri 37641 20529 37687 20574 sw
rect 70802 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
rect 37588 20516 37687 20529
tri 37687 20516 37699 20529 sw
rect 37588 20490 37699 20516
rect 37470 20471 37699 20490
tri 37699 20471 37745 20516 sw
rect 70802 20508 71000 20566
tri 37470 20425 37515 20471 ne
rect 37515 20425 37745 20471
tri 37745 20425 37790 20471 sw
rect 70802 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
tri 37515 20380 37561 20425 ne
rect 37561 20404 37790 20425
rect 37561 20380 37674 20404
tri 37561 20345 37596 20380 ne
rect 37596 20358 37674 20380
rect 37720 20380 37790 20404
tri 37790 20380 37835 20425 sw
rect 70802 20404 71000 20462
rect 37720 20358 37835 20380
rect 37596 20345 37835 20358
tri 37835 20345 37871 20380 sw
rect 70802 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
tri 37596 20299 37641 20345 ne
rect 37641 20299 37871 20345
tri 37871 20299 37916 20345 sw
rect 70802 20300 71000 20358
tri 37641 20254 37687 20299 ne
rect 37687 20272 37916 20299
rect 37687 20254 37806 20272
tri 37687 20209 37732 20254 ne
rect 37732 20226 37806 20254
rect 37852 20254 37916 20272
tri 37916 20254 37961 20299 sw
rect 70802 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 37852 20226 37961 20254
rect 37732 20209 37961 20226
tri 37961 20209 38006 20254 sw
tri 37732 20196 37745 20209 ne
rect 37745 20196 38006 20209
tri 38006 20196 38019 20209 sw
rect 70802 20196 71000 20254
tri 37745 20151 37790 20196 ne
rect 37790 20151 38019 20196
tri 38019 20151 38064 20196 sw
tri 37790 20106 37835 20151 ne
rect 37835 20140 38064 20151
rect 37835 20106 37938 20140
tri 37835 20061 37880 20106 ne
rect 37880 20094 37938 20106
rect 37984 20106 38064 20140
tri 38064 20106 38109 20151 sw
rect 70802 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
rect 37984 20094 38109 20106
rect 37880 20061 38109 20094
tri 38109 20061 38155 20106 sw
rect 70802 20092 71000 20150
tri 37880 20025 37916 20061 ne
rect 37916 20025 38155 20061
tri 38155 20025 38190 20061 sw
rect 70802 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
tri 37916 19980 37961 20025 ne
rect 37961 20008 38190 20025
rect 37961 19980 38070 20008
tri 37961 19935 38006 19980 ne
rect 38006 19962 38070 19980
rect 38116 19980 38190 20008
tri 38190 19980 38235 20025 sw
rect 70802 19988 71000 20046
rect 38116 19962 38235 19980
rect 38006 19935 38235 19962
tri 38235 19935 38281 19980 sw
rect 70802 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
tri 38006 19889 38051 19935 ne
rect 38051 19889 38281 19935
tri 38281 19889 38326 19935 sw
tri 38051 19877 38064 19889 ne
rect 38064 19877 38326 19889
tri 38326 19877 38339 19889 sw
rect 70802 19884 71000 19942
tri 38064 19831 38109 19877 ne
rect 38109 19876 38339 19877
rect 38109 19831 38202 19876
tri 38109 19786 38155 19831 ne
rect 38155 19830 38202 19831
rect 38248 19844 38339 19876
tri 38339 19844 38371 19877 sw
rect 38248 19830 38371 19844
rect 38155 19799 38371 19830
tri 38371 19799 38416 19844 sw
rect 70802 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
rect 38155 19786 38416 19799
tri 38155 19741 38200 19786 ne
rect 38200 19754 38416 19786
tri 38416 19754 38461 19799 sw
rect 70802 19780 71000 19838
rect 38200 19744 38461 19754
rect 38200 19741 38334 19744
tri 38200 19738 38203 19741 ne
rect 38203 19738 38334 19741
tri 38203 19693 38248 19738 ne
rect 38248 19698 38334 19738
rect 38380 19738 38461 19744
tri 38461 19738 38477 19754 sw
rect 38380 19698 38477 19738
rect 38248 19693 38477 19698
tri 38477 19693 38523 19738 sw
rect 70802 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
tri 38248 19647 38293 19693 ne
rect 38293 19647 38523 19693
tri 38523 19647 38568 19693 sw
rect 70802 19676 71000 19734
tri 38293 19602 38339 19647 ne
rect 38339 19612 38568 19647
rect 38339 19602 38466 19612
tri 38339 19570 38371 19602 ne
rect 38371 19570 38466 19602
tri 38371 19525 38416 19570 ne
rect 38416 19566 38466 19570
rect 38512 19602 38568 19612
tri 38568 19602 38613 19647 sw
rect 70802 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
rect 38512 19570 38613 19602
tri 38613 19570 38645 19602 sw
rect 70802 19572 71000 19630
rect 38512 19566 38645 19570
rect 38416 19525 38645 19566
tri 38645 19525 38691 19570 sw
rect 70802 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
tri 38416 19479 38461 19525 ne
rect 38461 19480 38691 19525
rect 38461 19479 38598 19480
tri 38461 19434 38507 19479 ne
rect 38507 19434 38598 19479
rect 38644 19479 38691 19480
tri 38691 19479 38736 19525 sw
rect 38644 19434 38736 19479
tri 38736 19434 38781 19479 sw
rect 70802 19468 71000 19526
tri 38507 19418 38523 19434 ne
rect 38523 19418 38781 19434
tri 38781 19418 38797 19434 sw
rect 70802 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
tri 38523 19373 38568 19418 ne
rect 38568 19373 38797 19418
tri 38797 19373 38842 19418 sw
tri 38568 19328 38613 19373 ne
rect 38613 19348 38842 19373
rect 38613 19328 38730 19348
tri 38613 19283 38658 19328 ne
rect 38658 19302 38730 19328
rect 38776 19328 38842 19348
tri 38842 19328 38887 19373 sw
rect 70802 19364 71000 19422
rect 38776 19302 38887 19328
rect 38658 19283 38887 19302
tri 38887 19283 38933 19328 sw
rect 70802 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
tri 38658 19250 38691 19283 ne
rect 38691 19250 38933 19283
tri 38933 19250 38965 19283 sw
rect 70802 19260 71000 19318
tri 38691 19205 38736 19250 ne
rect 38736 19216 38965 19250
rect 38736 19205 38862 19216
tri 38736 19160 38781 19205 ne
rect 38781 19170 38862 19205
rect 38908 19205 38965 19216
tri 38965 19205 39010 19250 sw
rect 70802 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 38908 19170 39010 19205
rect 38781 19160 39010 19170
tri 39010 19160 39055 19205 sw
tri 38781 19115 38826 19160 ne
rect 38826 19115 39055 19160
tri 39055 19115 39101 19160 sw
rect 70802 19156 71000 19214
tri 38826 19099 38842 19115 ne
rect 38842 19099 39101 19115
tri 39101 19099 39117 19115 sw
rect 70802 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
tri 38842 19053 38887 19099 ne
rect 38887 19084 39117 19099
rect 38887 19053 38994 19084
tri 38887 19008 38933 19053 ne
rect 38933 19038 38994 19053
rect 39040 19053 39117 19084
tri 39117 19053 39162 19099 sw
rect 39040 19038 39162 19053
rect 38933 19008 39162 19038
tri 39162 19008 39207 19053 sw
rect 70802 19052 71000 19110
tri 38933 18963 38978 19008 ne
rect 38978 18963 39207 19008
tri 39207 18963 39252 19008 sw
rect 70802 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
tri 38978 18931 39010 18963 ne
rect 39010 18952 39252 18963
rect 39010 18931 39126 18952
tri 39010 18885 39055 18931 ne
rect 39055 18906 39126 18931
rect 39172 18931 39252 18952
tri 39252 18931 39285 18963 sw
rect 70802 18948 71000 19006
rect 39172 18906 39285 18931
rect 39055 18885 39285 18906
tri 39285 18885 39330 18931 sw
rect 70802 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
tri 39055 18840 39101 18885 ne
rect 39101 18840 39330 18885
tri 39330 18840 39375 18885 sw
rect 70802 18844 71000 18902
tri 39101 18795 39146 18840 ne
rect 39146 18820 39375 18840
rect 39146 18795 39258 18820
tri 39146 18779 39162 18795 ne
rect 39162 18779 39258 18795
tri 39162 18734 39207 18779 ne
rect 39207 18774 39258 18779
rect 39304 18795 39375 18820
tri 39375 18795 39420 18840 sw
rect 70802 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 39304 18779 39420 18795
tri 39420 18779 39436 18795 sw
rect 39304 18774 39436 18779
rect 39207 18750 39436 18774
tri 39436 18750 39465 18779 sw
rect 39207 18734 39465 18750
tri 39207 18689 39252 18734 ne
rect 39252 18705 39465 18734
tri 39465 18705 39511 18750 sw
rect 70802 18740 71000 18798
rect 39252 18689 39511 18705
tri 39252 18643 39297 18689 ne
rect 39297 18688 39511 18689
rect 39297 18643 39390 18688
tri 39297 18640 39301 18643 ne
rect 39301 18642 39390 18643
rect 39436 18659 39511 18688
tri 39511 18659 39556 18705 sw
rect 70802 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
rect 39436 18642 39556 18659
rect 39301 18640 39556 18642
tri 39556 18640 39575 18659 sw
tri 39301 18595 39346 18640 ne
rect 39346 18595 39575 18640
tri 39575 18595 39620 18640 sw
rect 70802 18636 71000 18694
tri 39346 18550 39391 18595 ne
rect 39391 18556 39620 18595
rect 39391 18550 39522 18556
tri 39391 18505 39436 18550 ne
rect 39436 18510 39522 18550
rect 39568 18550 39620 18556
tri 39620 18550 39665 18595 sw
rect 70802 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
rect 39568 18510 39665 18550
rect 39436 18505 39665 18510
tri 39665 18505 39711 18550 sw
rect 70802 18532 71000 18590
tri 39436 18475 39465 18505 ne
rect 39465 18475 39711 18505
tri 39711 18475 39740 18505 sw
rect 70802 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
tri 39465 18430 39511 18475 ne
rect 39511 18430 39740 18475
tri 39740 18430 39785 18475 sw
tri 39511 18385 39556 18430 ne
rect 39556 18424 39785 18430
rect 39556 18385 39654 18424
tri 39556 18340 39601 18385 ne
rect 39601 18378 39654 18385
rect 39700 18385 39785 18424
tri 39785 18385 39830 18430 sw
rect 70802 18428 71000 18486
rect 39700 18378 39830 18385
rect 39601 18340 39830 18378
tri 39830 18340 39875 18385 sw
rect 70802 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
tri 39601 18321 39620 18340 ne
rect 39620 18321 39875 18340
tri 39875 18321 39895 18340 sw
rect 70802 18324 71000 18382
tri 39620 18275 39665 18321 ne
rect 39665 18292 39895 18321
rect 39665 18275 39786 18292
tri 39665 18230 39711 18275 ne
rect 39711 18246 39786 18275
rect 39832 18275 39895 18292
tri 39895 18275 39940 18321 sw
rect 70802 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
rect 39832 18246 39940 18275
rect 39711 18230 39940 18246
tri 39940 18230 39985 18275 sw
tri 39711 18185 39756 18230 ne
rect 39756 18185 39985 18230
tri 39985 18185 40030 18230 sw
rect 70802 18220 71000 18278
tri 39756 18156 39785 18185 ne
rect 39785 18160 40030 18185
rect 39785 18156 39918 18160
tri 39785 18111 39830 18156 ne
rect 39830 18114 39918 18156
rect 39964 18156 40030 18160
tri 40030 18156 40059 18185 sw
rect 70802 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
rect 39964 18114 40059 18156
rect 39830 18111 40059 18114
tri 40059 18111 40105 18156 sw
rect 70802 18116 71000 18174
tri 39830 18065 39875 18111 ne
rect 39875 18065 40105 18111
tri 40105 18065 40150 18111 sw
rect 70802 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
tri 39875 18020 39921 18065 ne
rect 39921 18028 40150 18065
rect 39921 18020 40050 18028
tri 39921 18001 39940 18020 ne
rect 39940 18001 40050 18020
tri 39940 17956 39985 18001 ne
rect 39985 17982 40050 18001
rect 40096 18020 40150 18028
tri 40150 18020 40195 18065 sw
rect 40096 18001 40195 18020
tri 40195 18001 40214 18020 sw
rect 70802 18012 71000 18070
rect 40096 17982 40214 18001
rect 39985 17956 40214 17982
tri 40214 17956 40259 18001 sw
rect 70802 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
tri 39985 17911 40030 17956 ne
rect 40030 17911 40259 17956
tri 40259 17911 40305 17956 sw
tri 40030 17865 40075 17911 ne
rect 40075 17896 40305 17911
rect 40075 17865 40182 17896
tri 40075 17836 40105 17865 ne
rect 40105 17850 40182 17865
rect 40228 17865 40305 17896
tri 40305 17865 40350 17911 sw
rect 70802 17908 71000 17966
rect 40228 17850 40350 17865
rect 40105 17836 40350 17850
tri 40350 17836 40379 17865 sw
rect 70802 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
tri 40105 17791 40150 17836 ne
rect 40150 17791 40379 17836
tri 40379 17791 40424 17836 sw
rect 70802 17804 71000 17862
tri 40150 17746 40195 17791 ne
rect 40195 17764 40424 17791
rect 40195 17746 40314 17764
tri 40195 17701 40240 17746 ne
rect 40240 17718 40314 17746
rect 40360 17746 40424 17764
tri 40424 17746 40469 17791 sw
rect 70802 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 40360 17718 40469 17746
rect 40240 17701 40469 17718
tri 40469 17701 40515 17746 sw
tri 40240 17681 40259 17701 ne
rect 40259 17681 40515 17701
tri 40515 17681 40534 17701 sw
rect 70802 17700 71000 17758
tri 40259 17636 40305 17681 ne
rect 40305 17655 40534 17681
tri 40534 17655 40560 17681 sw
rect 40305 17636 40560 17655
tri 40305 17591 40350 17636 ne
rect 40350 17632 40560 17636
rect 40350 17591 40446 17632
tri 40350 17546 40395 17591 ne
rect 40395 17586 40446 17591
rect 40492 17610 40560 17632
tri 40560 17610 40605 17655 sw
rect 70802 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
rect 40492 17586 40605 17610
rect 40395 17565 40605 17586
tri 40605 17565 40650 17610 sw
rect 70802 17596 71000 17654
rect 40395 17546 40650 17565
tri 40395 17543 40398 17546 ne
rect 40398 17543 40650 17546
tri 40650 17543 40673 17565 sw
rect 70802 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
tri 40398 17497 40443 17543 ne
rect 40443 17500 40673 17543
rect 40443 17497 40578 17500
tri 40443 17452 40489 17497 ne
rect 40489 17454 40578 17497
rect 40624 17497 40673 17500
tri 40673 17497 40718 17543 sw
rect 40624 17454 40718 17497
rect 40489 17452 40718 17454
tri 40718 17452 40763 17497 sw
rect 70802 17492 71000 17550
tri 40489 17407 40534 17452 ne
rect 40534 17407 40763 17452
tri 40763 17407 40808 17452 sw
rect 70802 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
tri 40534 17381 40560 17407 ne
rect 40560 17381 40808 17407
tri 40808 17381 40834 17407 sw
rect 70802 17388 71000 17446
tri 40560 17336 40605 17381 ne
rect 40605 17368 40834 17381
rect 40605 17336 40710 17368
tri 40605 17291 40650 17336 ne
rect 40650 17322 40710 17336
rect 40756 17336 40834 17368
tri 40834 17336 40879 17381 sw
rect 70802 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 40756 17322 40879 17336
rect 40650 17291 40879 17322
tri 40879 17291 40925 17336 sw
tri 40650 17245 40695 17291 ne
rect 40695 17245 40925 17291
tri 40925 17245 40970 17291 sw
rect 70802 17284 71000 17342
tri 40695 17223 40718 17245 ne
rect 40718 17236 40970 17245
rect 40718 17223 40842 17236
tri 40718 17178 40763 17223 ne
rect 40763 17190 40842 17223
rect 40888 17223 40970 17236
tri 40970 17223 40992 17245 sw
rect 70802 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
rect 40888 17190 40992 17223
rect 40763 17178 40992 17190
tri 40992 17178 41037 17223 sw
rect 70802 17180 71000 17238
tri 40763 17133 40808 17178 ne
rect 40808 17133 41037 17178
tri 41037 17133 41083 17178 sw
rect 70802 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
tri 40808 17087 40853 17133 ne
rect 40853 17104 41083 17133
rect 40853 17087 40974 17104
tri 40853 17061 40879 17087 ne
rect 40879 17061 40974 17087
tri 40879 17016 40925 17061 ne
rect 40925 17058 40974 17061
rect 41020 17087 41083 17104
tri 41083 17087 41128 17133 sw
rect 41020 17061 41128 17087
tri 41128 17061 41154 17087 sw
rect 70802 17076 71000 17134
rect 41020 17058 41154 17061
rect 40925 17016 41154 17058
tri 41154 17016 41199 17061 sw
rect 70802 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
tri 40925 16971 40970 17016 ne
rect 40970 16972 41199 17016
rect 40970 16971 41106 16972
tri 40970 16926 41015 16971 ne
rect 41015 16926 41106 16971
rect 41152 16971 41199 16972
tri 41199 16971 41244 17016 sw
rect 70802 16972 71000 17030
rect 41152 16926 41244 16971
tri 41244 16926 41289 16971 sw
rect 70802 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
tri 41015 16903 41037 16926 ne
rect 41037 16903 41289 16926
tri 41289 16903 41312 16926 sw
tri 41037 16858 41083 16903 ne
rect 41083 16858 41312 16903
tri 41312 16858 41357 16903 sw
rect 70802 16868 71000 16926
tri 41083 16813 41128 16858 ne
rect 41128 16840 41357 16858
rect 41128 16813 41238 16840
tri 41128 16768 41173 16813 ne
rect 41173 16794 41238 16813
rect 41284 16813 41357 16840
tri 41357 16813 41402 16858 sw
rect 70802 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 41284 16794 41402 16813
rect 41173 16768 41402 16794
tri 41402 16768 41447 16813 sw
tri 41173 16742 41199 16768 ne
rect 41199 16742 41447 16768
tri 41447 16742 41473 16768 sw
rect 70802 16764 71000 16822
tri 41199 16697 41244 16742 ne
rect 41244 16708 41473 16742
rect 41244 16697 41370 16708
tri 41244 16651 41289 16697 ne
rect 41289 16662 41370 16697
rect 41416 16697 41473 16708
tri 41473 16697 41519 16742 sw
rect 70802 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
rect 41416 16662 41519 16697
rect 41289 16651 41519 16662
tri 41519 16651 41564 16697 sw
rect 70802 16660 71000 16718
tri 41289 16606 41335 16651 ne
rect 41335 16606 41564 16651
tri 41564 16606 41609 16651 sw
rect 70802 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
tri 41335 16584 41357 16606 ne
rect 41357 16584 41609 16606
tri 41609 16584 41631 16606 sw
tri 41357 16539 41402 16584 ne
rect 41402 16576 41631 16584
rect 41402 16539 41502 16576
tri 41402 16493 41447 16539 ne
rect 41447 16530 41502 16539
rect 41548 16561 41631 16576
tri 41631 16561 41654 16584 sw
rect 41548 16530 41654 16561
rect 41447 16516 41654 16530
tri 41654 16516 41699 16561 sw
rect 70802 16556 71000 16614
rect 41447 16493 41699 16516
tri 41447 16448 41493 16493 ne
rect 41493 16471 41699 16493
tri 41699 16471 41745 16516 sw
rect 70802 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
rect 41493 16448 41745 16471
tri 41493 16445 41496 16448 ne
rect 41496 16445 41745 16448
tri 41745 16445 41770 16471 sw
rect 70802 16452 71000 16510
tri 41496 16400 41541 16445 ne
rect 41541 16444 41770 16445
rect 41541 16400 41634 16444
tri 41541 16355 41586 16400 ne
rect 41586 16398 41634 16400
rect 41680 16400 41770 16444
tri 41770 16400 41815 16445 sw
rect 70802 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
rect 41680 16398 41815 16400
rect 41586 16355 41815 16398
tri 41815 16355 41861 16400 sw
tri 41586 16309 41631 16355 ne
rect 41631 16312 41861 16355
rect 41631 16309 41766 16312
tri 41631 16287 41654 16309 ne
rect 41654 16287 41766 16309
tri 41654 16241 41699 16287 ne
rect 41699 16266 41766 16287
rect 41812 16309 41861 16312
tri 41861 16309 41906 16355 sw
rect 70802 16348 71000 16406
rect 41812 16287 41906 16309
tri 41906 16287 41929 16309 sw
rect 70802 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 41812 16266 41929 16287
rect 41699 16241 41929 16266
tri 41929 16241 41974 16287 sw
rect 70802 16244 71000 16302
tri 41699 16196 41745 16241 ne
rect 41745 16196 41974 16241
tri 41974 16196 42019 16241 sw
rect 70802 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
tri 41745 16151 41790 16196 ne
rect 41790 16180 42019 16196
rect 41790 16151 41898 16180
tri 41790 16125 41815 16151 ne
rect 41815 16134 41898 16151
rect 41944 16151 42019 16180
tri 42019 16151 42064 16196 sw
rect 41944 16134 42064 16151
rect 41815 16125 42064 16134
tri 42064 16125 42090 16151 sw
rect 70802 16140 71000 16198
tri 41815 16080 41861 16125 ne
rect 41861 16080 42090 16125
tri 42090 16080 42135 16125 sw
rect 70802 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
tri 41861 16035 41906 16080 ne
rect 41906 16048 42135 16080
rect 41906 16035 42030 16048
tri 41906 15990 41951 16035 ne
rect 41951 16002 42030 16035
rect 42076 16035 42135 16048
tri 42135 16035 42180 16080 sw
rect 70802 16036 71000 16094
rect 42076 16002 42180 16035
rect 41951 15990 42180 16002
tri 42180 15990 42225 16035 sw
rect 70802 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
tri 41951 15967 41974 15990 ne
rect 41974 15967 42225 15990
tri 42225 15967 42248 15990 sw
tri 41974 15922 42019 15967 ne
rect 42019 15922 42248 15967
tri 42248 15922 42293 15967 sw
rect 70802 15932 71000 15990
tri 42019 15877 42064 15922 ne
rect 42064 15916 42293 15922
rect 42064 15877 42162 15916
tri 42064 15831 42109 15877 ne
rect 42109 15870 42162 15877
rect 42208 15877 42293 15916
tri 42293 15877 42339 15922 sw
rect 70802 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
rect 42208 15870 42339 15877
rect 42109 15831 42339 15870
tri 42339 15831 42384 15877 sw
tri 42109 15806 42135 15831 ne
rect 42135 15806 42384 15831
tri 42384 15806 42409 15831 sw
rect 70802 15828 71000 15886
tri 42135 15761 42180 15806 ne
rect 42180 15784 42409 15806
rect 42180 15761 42294 15784
tri 42180 15715 42225 15761 ne
rect 42225 15738 42294 15761
rect 42340 15761 42409 15784
tri 42409 15761 42455 15806 sw
rect 70802 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 42340 15738 42455 15761
rect 42225 15715 42455 15738
tri 42455 15715 42500 15761 sw
rect 70802 15724 71000 15782
tri 42225 15670 42271 15715 ne
rect 42271 15670 42500 15715
tri 42500 15670 42545 15715 sw
rect 70802 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
tri 42271 15647 42293 15670 ne
rect 42293 15652 42545 15670
rect 42293 15647 42426 15652
tri 42293 15602 42339 15647 ne
rect 42339 15606 42426 15647
rect 42472 15647 42545 15652
tri 42545 15647 42568 15670 sw
rect 42472 15606 42568 15647
rect 42339 15602 42568 15606
tri 42568 15602 42613 15647 sw
rect 70802 15620 71000 15678
tri 42339 15557 42384 15602 ne
rect 42384 15557 42613 15602
tri 42613 15557 42658 15602 sw
rect 70802 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
tri 42384 15512 42429 15557 ne
rect 42429 15520 42658 15557
rect 42429 15512 42558 15520
tri 42429 15486 42455 15512 ne
rect 42455 15486 42558 15512
tri 42455 15441 42500 15486 ne
rect 42500 15474 42558 15486
rect 42604 15512 42658 15520
tri 42658 15512 42703 15557 sw
rect 70802 15516 71000 15574
rect 42604 15486 42703 15512
tri 42703 15486 42729 15512 sw
rect 42604 15474 42729 15486
rect 42500 15467 42729 15474
tri 42729 15467 42749 15486 sw
rect 70802 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
rect 42500 15441 42749 15467
tri 42500 15396 42545 15441 ne
rect 42545 15421 42749 15441
tri 42749 15421 42794 15467 sw
rect 42545 15396 42794 15421
tri 42545 15351 42590 15396 ne
rect 42590 15388 42794 15396
rect 42590 15351 42690 15388
tri 42590 15347 42593 15351 ne
rect 42593 15347 42690 15351
tri 42593 15302 42639 15347 ne
rect 42639 15342 42690 15347
rect 42736 15376 42794 15388
tri 42794 15376 42839 15421 sw
rect 70802 15412 71000 15470
rect 42736 15347 42839 15376
tri 42839 15347 42868 15376 sw
rect 70802 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 42736 15342 42868 15347
rect 42639 15302 42868 15342
tri 42868 15302 42913 15347 sw
rect 70802 15308 71000 15366
tri 42639 15257 42684 15302 ne
rect 42684 15257 42913 15302
tri 42913 15257 42958 15302 sw
rect 70802 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
tri 42684 15212 42729 15257 ne
rect 42729 15256 42958 15257
rect 42729 15212 42822 15256
tri 42729 15192 42749 15212 ne
rect 42749 15210 42822 15212
rect 42868 15212 42958 15256
tri 42958 15212 43003 15257 sw
rect 42868 15210 43003 15212
rect 42749 15192 43003 15210
tri 43003 15192 43023 15212 sw
rect 70802 15204 71000 15262
tri 42749 15147 42794 15192 ne
rect 42794 15147 43023 15192
tri 43023 15147 43068 15192 sw
rect 70802 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
tri 42794 15102 42839 15147 ne
rect 42839 15124 43068 15147
rect 42839 15102 42954 15124
tri 42839 15057 42884 15102 ne
rect 42884 15078 42954 15102
rect 43000 15102 43068 15124
tri 43068 15102 43113 15147 sw
rect 43000 15078 43113 15102
rect 42884 15057 43113 15078
tri 43113 15057 43159 15102 sw
rect 70802 15100 71000 15158
tri 42884 15028 42913 15057 ne
rect 42913 15028 43159 15057
tri 43159 15028 43187 15057 sw
rect 70802 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
tri 42913 14983 42958 15028 ne
rect 42958 14992 43187 15028
rect 42958 14983 43086 14992
tri 42958 14937 43003 14983 ne
rect 43003 14946 43086 14983
rect 43132 14983 43187 14992
tri 43187 14983 43233 15028 sw
rect 70802 14996 71000 15054
rect 43132 14946 43233 14983
rect 43003 14937 43233 14946
tri 43233 14937 43278 14983 sw
rect 70802 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
tri 43003 14892 43049 14937 ne
rect 43049 14892 43278 14937
tri 43278 14892 43323 14937 sw
rect 70802 14892 71000 14950
tri 43049 14873 43068 14892 ne
rect 43068 14873 43323 14892
tri 43323 14873 43343 14892 sw
tri 43068 14827 43113 14873 ne
rect 43113 14860 43343 14873
rect 43113 14827 43218 14860
tri 43113 14782 43159 14827 ne
rect 43159 14814 43218 14827
rect 43264 14827 43343 14860
tri 43343 14827 43388 14873 sw
rect 70802 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
rect 43264 14814 43388 14827
rect 43159 14782 43388 14814
tri 43388 14782 43433 14827 sw
rect 70802 14788 71000 14846
tri 43159 14737 43204 14782 ne
rect 43204 14737 43433 14782
tri 43433 14737 43478 14782 sw
rect 70802 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
tri 43204 14708 43233 14737 ne
rect 43233 14728 43478 14737
rect 43233 14708 43350 14728
tri 43233 14663 43278 14708 ne
rect 43278 14682 43350 14708
rect 43396 14708 43478 14728
tri 43478 14708 43507 14737 sw
rect 43396 14682 43507 14708
rect 43278 14663 43507 14682
tri 43507 14663 43552 14708 sw
rect 70802 14684 71000 14742
tri 43278 14618 43323 14663 ne
rect 43323 14618 43552 14663
tri 43552 14618 43597 14663 sw
rect 70802 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
tri 43323 14573 43368 14618 ne
rect 43368 14596 43597 14618
rect 43368 14573 43482 14596
tri 43368 14553 43388 14573 ne
rect 43388 14553 43482 14573
tri 43388 14508 43433 14553 ne
rect 43433 14550 43482 14553
rect 43528 14573 43597 14596
tri 43597 14573 43643 14618 sw
rect 70802 14580 71000 14638
rect 43528 14553 43643 14573
tri 43643 14553 43662 14573 sw
rect 43528 14550 43662 14553
rect 43433 14508 43662 14550
tri 43662 14508 43707 14553 sw
rect 70802 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
tri 43433 14463 43478 14508 ne
rect 43478 14464 43707 14508
rect 43478 14463 43614 14464
tri 43478 14417 43523 14463 ne
rect 43523 14418 43614 14463
rect 43660 14463 43707 14464
tri 43707 14463 43753 14508 sw
rect 70802 14476 71000 14534
rect 43660 14418 43753 14463
rect 43523 14417 43753 14418
tri 43753 14417 43798 14463 sw
rect 70802 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
tri 43523 14389 43552 14417 ne
rect 43552 14389 43798 14417
tri 43798 14389 43827 14417 sw
tri 43552 14343 43597 14389 ne
rect 43597 14372 43827 14389
tri 43827 14372 43843 14389 sw
rect 70802 14372 71000 14430
rect 43597 14343 43843 14372
tri 43597 14298 43643 14343 ne
rect 43643 14332 43843 14343
rect 43643 14298 43746 14332
tri 43643 14253 43688 14298 ne
rect 43688 14286 43746 14298
rect 43792 14327 43843 14332
tri 43843 14327 43888 14372 sw
rect 43792 14286 43888 14327
rect 43688 14282 43888 14286
tri 43888 14282 43933 14327 sw
rect 70802 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 43688 14253 43933 14282
tri 43688 14250 43691 14253 ne
rect 43691 14250 43933 14253
tri 43933 14250 43965 14282 sw
rect 70802 14268 71000 14326
tri 43691 14205 43736 14250 ne
rect 43736 14205 43965 14250
tri 43965 14205 44011 14250 sw
rect 70802 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
tri 43736 14159 43781 14205 ne
rect 43781 14200 44011 14205
rect 43781 14159 43878 14200
tri 43781 14114 43827 14159 ne
rect 43827 14154 43878 14159
rect 43924 14159 44011 14200
tri 44011 14159 44056 14205 sw
rect 70802 14164 71000 14222
rect 43924 14154 44056 14159
rect 43827 14114 44056 14154
tri 44056 14114 44101 14159 sw
rect 70802 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
tri 43827 14098 43843 14114 ne
rect 43843 14098 44101 14114
tri 44101 14098 44117 14114 sw
tri 43843 14053 43888 14098 ne
rect 43888 14068 44117 14098
rect 43888 14053 44010 14068
tri 43888 14007 43933 14053 ne
rect 43933 14022 44010 14053
rect 44056 14053 44117 14068
tri 44117 14053 44163 14098 sw
rect 70802 14060 71000 14118
rect 44056 14022 44163 14053
rect 43933 14007 44163 14022
tri 44163 14007 44208 14053 sw
rect 70802 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
tri 43933 13962 43979 14007 ne
rect 43979 13962 44208 14007
tri 44208 13962 44253 14007 sw
tri 43979 13930 44011 13962 ne
rect 44011 13936 44253 13962
rect 44011 13930 44142 13936
tri 44011 13885 44056 13930 ne
rect 44056 13890 44142 13930
rect 44188 13930 44253 13936
tri 44253 13930 44285 13962 sw
rect 70802 13956 71000 14014
rect 44188 13890 44285 13930
rect 44056 13885 44285 13890
tri 44285 13885 44330 13930 sw
rect 70802 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
tri 44056 13840 44101 13885 ne
rect 44101 13840 44330 13885
tri 44330 13840 44375 13885 sw
rect 70802 13852 71000 13910
tri 44101 13795 44146 13840 ne
rect 44146 13804 44375 13840
rect 44146 13795 44274 13804
tri 44146 13778 44163 13795 ne
rect 44163 13778 44274 13795
tri 44163 13733 44208 13778 ne
rect 44208 13758 44274 13778
rect 44320 13795 44375 13804
tri 44375 13795 44421 13840 sw
rect 70802 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
rect 44320 13778 44421 13795
tri 44421 13778 44437 13795 sw
rect 44320 13758 44437 13778
rect 44208 13733 44437 13758
tri 44437 13733 44482 13778 sw
rect 70802 13748 71000 13806
tri 44208 13688 44253 13733 ne
rect 44253 13688 44482 13733
tri 44482 13688 44527 13733 sw
rect 70802 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
tri 44253 13643 44298 13688 ne
rect 44298 13672 44527 13688
rect 44298 13643 44406 13672
tri 44298 13611 44330 13643 ne
rect 44330 13626 44406 13643
rect 44452 13643 44527 13672
tri 44527 13643 44573 13688 sw
rect 70802 13644 71000 13702
rect 44452 13626 44573 13643
rect 44330 13611 44573 13626
tri 44573 13611 44605 13643 sw
tri 44330 13565 44375 13611 ne
rect 44375 13565 44605 13611
tri 44605 13565 44650 13611 sw
rect 70802 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
tri 44375 13520 44421 13565 ne
rect 44421 13540 44650 13565
rect 44421 13520 44538 13540
tri 44421 13475 44466 13520 ne
rect 44466 13494 44538 13520
rect 44584 13520 44650 13540
tri 44650 13520 44695 13565 sw
rect 70802 13540 71000 13598
rect 44584 13494 44695 13520
rect 44466 13475 44695 13494
tri 44695 13475 44740 13520 sw
rect 70802 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
tri 44466 13459 44482 13475 ne
rect 44482 13459 44740 13475
tri 44740 13459 44757 13475 sw
tri 44482 13413 44527 13459 ne
rect 44527 13413 44757 13459
tri 44757 13413 44802 13459 sw
rect 70802 13436 71000 13494
tri 44527 13368 44573 13413 ne
rect 44573 13408 44802 13413
rect 44573 13368 44670 13408
tri 44573 13323 44618 13368 ne
rect 44618 13362 44670 13368
rect 44716 13368 44802 13408
tri 44802 13368 44847 13413 sw
rect 70802 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 44716 13362 44847 13368
rect 44618 13323 44847 13362
tri 44847 13323 44892 13368 sw
tri 44618 13291 44650 13323 ne
rect 44650 13291 44892 13323
tri 44892 13291 44924 13323 sw
rect 70802 13291 71000 13390
tri 44650 13246 44695 13291 ne
rect 44695 13269 71000 13291
rect 44695 13256 45088 13269
rect 44695 13246 44850 13256
tri 44695 13201 44740 13246 ne
rect 44740 13210 44850 13246
rect 44896 13223 45088 13256
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 44896 13210 71000 13223
rect 44740 13201 71000 13210
tri 44740 13155 44785 13201 ne
rect 44785 13165 71000 13201
rect 44785 13155 45088 13165
tri 44785 13110 44831 13155 ne
rect 44831 13119 45088 13155
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
rect 44831 13110 71000 13119
tri 44831 13097 44844 13110 ne
rect 44844 13097 71000 13110
<< psubdiffcont >>
rect 13119 70929 13165 70975
rect 13223 70929 13269 70975
rect 13377 70929 13423 70975
rect 13481 70929 13527 70975
rect 13585 70929 13631 70975
rect 13689 70929 13735 70975
rect 13793 70929 13839 70975
rect 13897 70929 13943 70975
rect 14001 70929 14047 70975
rect 14105 70929 14151 70975
rect 14209 70929 14255 70975
rect 14313 70929 14359 70975
rect 14417 70929 14463 70975
rect 14521 70929 14567 70975
rect 14625 70929 14671 70975
rect 14729 70929 14775 70975
rect 14833 70929 14879 70975
rect 14937 70929 14983 70975
rect 15041 70929 15087 70975
rect 15145 70929 15191 70975
rect 15249 70929 15295 70975
rect 15353 70929 15399 70975
rect 15457 70929 15503 70975
rect 15561 70929 15607 70975
rect 15665 70929 15711 70975
rect 15769 70929 15815 70975
rect 15873 70929 15919 70975
rect 15977 70929 16023 70975
rect 16081 70929 16127 70975
rect 16185 70929 16231 70975
rect 16289 70929 16335 70975
rect 16393 70929 16439 70975
rect 16497 70929 16543 70975
rect 16601 70929 16647 70975
rect 16705 70929 16751 70975
rect 16809 70929 16855 70975
rect 16913 70929 16959 70975
rect 17017 70929 17063 70975
rect 17121 70929 17167 70975
rect 17225 70929 17271 70975
rect 17329 70929 17375 70975
rect 17433 70929 17479 70975
rect 17537 70929 17583 70975
rect 17641 70929 17687 70975
rect 17745 70929 17791 70975
rect 17849 70929 17895 70975
rect 17953 70929 17999 70975
rect 18057 70929 18103 70975
rect 18161 70929 18207 70975
rect 18265 70929 18311 70975
rect 18369 70929 18415 70975
rect 18473 70929 18519 70975
rect 18577 70929 18623 70975
rect 18681 70929 18727 70975
rect 18785 70929 18831 70975
rect 18889 70929 18935 70975
rect 18993 70929 19039 70975
rect 19097 70929 19143 70975
rect 19201 70929 19247 70975
rect 19305 70929 19351 70975
rect 19409 70929 19455 70975
rect 19513 70929 19559 70975
rect 19617 70929 19663 70975
rect 19721 70929 19767 70975
rect 19825 70929 19871 70975
rect 19929 70929 19975 70975
rect 20033 70929 20079 70975
rect 20137 70929 20183 70975
rect 20241 70929 20287 70975
rect 20345 70929 20391 70975
rect 20449 70929 20495 70975
rect 20553 70929 20599 70975
rect 20657 70929 20703 70975
rect 20761 70929 20807 70975
rect 20865 70929 20911 70975
rect 20969 70929 21015 70975
rect 21073 70929 21119 70975
rect 21177 70929 21223 70975
rect 21281 70929 21327 70975
rect 21385 70929 21431 70975
rect 21489 70929 21535 70975
rect 21593 70929 21639 70975
rect 21697 70929 21743 70975
rect 21801 70929 21847 70975
rect 21905 70929 21951 70975
rect 22009 70929 22055 70975
rect 22113 70929 22159 70975
rect 22217 70929 22263 70975
rect 22321 70929 22367 70975
rect 22425 70929 22471 70975
rect 22529 70929 22575 70975
rect 22633 70929 22679 70975
rect 22737 70929 22783 70975
rect 22841 70929 22887 70975
rect 22945 70929 22991 70975
rect 23049 70929 23095 70975
rect 23153 70929 23199 70975
rect 23257 70929 23303 70975
rect 23361 70929 23407 70975
rect 23465 70929 23511 70975
rect 23569 70929 23615 70975
rect 23673 70929 23719 70975
rect 23777 70929 23823 70975
rect 23881 70929 23927 70975
rect 23985 70929 24031 70975
rect 24089 70929 24135 70975
rect 24193 70929 24239 70975
rect 24297 70929 24343 70975
rect 24401 70929 24447 70975
rect 24505 70929 24551 70975
rect 24609 70929 24655 70975
rect 24713 70929 24759 70975
rect 24817 70929 24863 70975
rect 24921 70929 24967 70975
rect 25025 70929 25071 70975
rect 25129 70929 25175 70975
rect 25233 70929 25279 70975
rect 25337 70929 25383 70975
rect 25441 70929 25487 70975
rect 25545 70929 25591 70975
rect 25649 70929 25695 70975
rect 25753 70929 25799 70975
rect 25857 70929 25903 70975
rect 25961 70929 26007 70975
rect 26065 70929 26111 70975
rect 26169 70929 26215 70975
rect 26273 70929 26319 70975
rect 26377 70929 26423 70975
rect 26481 70929 26527 70975
rect 26585 70929 26631 70975
rect 26689 70929 26735 70975
rect 26793 70929 26839 70975
rect 26897 70929 26943 70975
rect 27001 70929 27047 70975
rect 27105 70929 27151 70975
rect 27209 70929 27255 70975
rect 27313 70929 27359 70975
rect 27417 70929 27463 70975
rect 27521 70929 27567 70975
rect 27625 70929 27671 70975
rect 27729 70929 27775 70975
rect 27833 70929 27879 70975
rect 27937 70929 27983 70975
rect 28041 70929 28087 70975
rect 28145 70929 28191 70975
rect 28249 70929 28295 70975
rect 28353 70929 28399 70975
rect 28457 70929 28503 70975
rect 28561 70929 28607 70975
rect 28665 70929 28711 70975
rect 28769 70929 28815 70975
rect 28873 70929 28919 70975
rect 28977 70929 29023 70975
rect 29081 70929 29127 70975
rect 29185 70929 29231 70975
rect 29289 70929 29335 70975
rect 29393 70929 29439 70975
rect 29497 70929 29543 70975
rect 29601 70929 29647 70975
rect 29705 70929 29751 70975
rect 29809 70929 29855 70975
rect 29913 70929 29959 70975
rect 30017 70929 30063 70975
rect 30121 70929 30167 70975
rect 30225 70929 30271 70975
rect 30329 70929 30375 70975
rect 30433 70929 30479 70975
rect 30537 70929 30583 70975
rect 30641 70929 30687 70975
rect 30745 70929 30791 70975
rect 30849 70929 30895 70975
rect 30953 70929 30999 70975
rect 31057 70929 31103 70975
rect 31161 70929 31207 70975
rect 31265 70929 31311 70975
rect 31369 70929 31415 70975
rect 31473 70929 31519 70975
rect 31577 70929 31623 70975
rect 31681 70929 31727 70975
rect 31785 70929 31831 70975
rect 31889 70929 31935 70975
rect 31993 70929 32039 70975
rect 32097 70929 32143 70975
rect 32201 70929 32247 70975
rect 32305 70929 32351 70975
rect 32409 70929 32455 70975
rect 32513 70929 32559 70975
rect 32617 70929 32663 70975
rect 32721 70929 32767 70975
rect 32825 70929 32871 70975
rect 32929 70929 32975 70975
rect 33033 70929 33079 70975
rect 33137 70929 33183 70975
rect 33241 70929 33287 70975
rect 33345 70929 33391 70975
rect 33449 70929 33495 70975
rect 33553 70929 33599 70975
rect 33657 70929 33703 70975
rect 33761 70929 33807 70975
rect 33865 70929 33911 70975
rect 33969 70929 34015 70975
rect 34073 70929 34119 70975
rect 34177 70929 34223 70975
rect 34281 70929 34327 70975
rect 34385 70929 34431 70975
rect 34489 70929 34535 70975
rect 34593 70929 34639 70975
rect 34697 70929 34743 70975
rect 34801 70929 34847 70975
rect 34905 70929 34951 70975
rect 35009 70929 35055 70975
rect 35113 70929 35159 70975
rect 35217 70929 35263 70975
rect 35321 70929 35367 70975
rect 35425 70929 35471 70975
rect 35529 70929 35575 70975
rect 35633 70929 35679 70975
rect 35737 70929 35783 70975
rect 35841 70929 35887 70975
rect 35945 70929 35991 70975
rect 36049 70929 36095 70975
rect 36153 70929 36199 70975
rect 36257 70929 36303 70975
rect 36361 70929 36407 70975
rect 36465 70929 36511 70975
rect 36569 70929 36615 70975
rect 36673 70929 36719 70975
rect 36777 70929 36823 70975
rect 36881 70929 36927 70975
rect 36985 70929 37031 70975
rect 37089 70929 37135 70975
rect 37193 70929 37239 70975
rect 37297 70929 37343 70975
rect 37401 70929 37447 70975
rect 37505 70929 37551 70975
rect 37609 70929 37655 70975
rect 37713 70929 37759 70975
rect 37817 70929 37863 70975
rect 37921 70929 37967 70975
rect 38025 70929 38071 70975
rect 38129 70929 38175 70975
rect 38233 70929 38279 70975
rect 38337 70929 38383 70975
rect 38441 70929 38487 70975
rect 38545 70929 38591 70975
rect 38649 70929 38695 70975
rect 38753 70929 38799 70975
rect 38857 70929 38903 70975
rect 38961 70929 39007 70975
rect 39065 70929 39111 70975
rect 39169 70929 39215 70975
rect 39273 70929 39319 70975
rect 39377 70929 39423 70975
rect 39481 70929 39527 70975
rect 39585 70929 39631 70975
rect 39689 70929 39735 70975
rect 39793 70929 39839 70975
rect 39897 70929 39943 70975
rect 40001 70929 40047 70975
rect 40105 70929 40151 70975
rect 40209 70929 40255 70975
rect 40313 70929 40359 70975
rect 40417 70929 40463 70975
rect 40521 70929 40567 70975
rect 40625 70929 40671 70975
rect 40729 70929 40775 70975
rect 40833 70929 40879 70975
rect 40937 70929 40983 70975
rect 41041 70929 41087 70975
rect 41145 70929 41191 70975
rect 41249 70929 41295 70975
rect 41353 70929 41399 70975
rect 41457 70929 41503 70975
rect 41561 70929 41607 70975
rect 41665 70929 41711 70975
rect 41769 70929 41815 70975
rect 41873 70929 41919 70975
rect 41977 70929 42023 70975
rect 42081 70929 42127 70975
rect 42185 70929 42231 70975
rect 42289 70929 42335 70975
rect 42393 70929 42439 70975
rect 42497 70929 42543 70975
rect 42601 70929 42647 70975
rect 42705 70929 42751 70975
rect 42809 70929 42855 70975
rect 42913 70929 42959 70975
rect 43017 70929 43063 70975
rect 43121 70929 43167 70975
rect 43225 70929 43271 70975
rect 43329 70929 43375 70975
rect 43433 70929 43479 70975
rect 43537 70929 43583 70975
rect 43641 70929 43687 70975
rect 43745 70929 43791 70975
rect 43849 70929 43895 70975
rect 43953 70929 43999 70975
rect 44057 70929 44103 70975
rect 44161 70929 44207 70975
rect 44265 70929 44311 70975
rect 44369 70929 44415 70975
rect 44473 70929 44519 70975
rect 44577 70929 44623 70975
rect 44681 70929 44727 70975
rect 44785 70929 44831 70975
rect 44889 70929 44935 70975
rect 44993 70929 45039 70975
rect 45097 70929 45143 70975
rect 45201 70929 45247 70975
rect 45305 70929 45351 70975
rect 45409 70929 45455 70975
rect 45513 70929 45559 70975
rect 45617 70929 45663 70975
rect 45721 70929 45767 70975
rect 45825 70929 45871 70975
rect 45929 70929 45975 70975
rect 46033 70929 46079 70975
rect 46137 70929 46183 70975
rect 46241 70929 46287 70975
rect 46345 70929 46391 70975
rect 46449 70929 46495 70975
rect 46553 70929 46599 70975
rect 46657 70929 46703 70975
rect 46761 70929 46807 70975
rect 46865 70929 46911 70975
rect 46969 70929 47015 70975
rect 47073 70929 47119 70975
rect 47177 70929 47223 70975
rect 47281 70929 47327 70975
rect 47385 70929 47431 70975
rect 47489 70929 47535 70975
rect 47593 70929 47639 70975
rect 47697 70929 47743 70975
rect 47801 70929 47847 70975
rect 47905 70929 47951 70975
rect 48009 70929 48055 70975
rect 48113 70929 48159 70975
rect 48217 70929 48263 70975
rect 48321 70929 48367 70975
rect 48425 70929 48471 70975
rect 48529 70929 48575 70975
rect 48633 70929 48679 70975
rect 48737 70929 48783 70975
rect 48841 70929 48887 70975
rect 48945 70929 48991 70975
rect 49049 70929 49095 70975
rect 49153 70929 49199 70975
rect 49257 70929 49303 70975
rect 49361 70929 49407 70975
rect 49465 70929 49511 70975
rect 49569 70929 49615 70975
rect 49673 70929 49719 70975
rect 49777 70929 49823 70975
rect 49881 70929 49927 70975
rect 49985 70929 50031 70975
rect 50089 70929 50135 70975
rect 50193 70929 50239 70975
rect 50297 70929 50343 70975
rect 50401 70929 50447 70975
rect 50505 70929 50551 70975
rect 50609 70929 50655 70975
rect 50713 70929 50759 70975
rect 50817 70929 50863 70975
rect 50921 70929 50967 70975
rect 51025 70929 51071 70975
rect 51129 70929 51175 70975
rect 51233 70929 51279 70975
rect 51337 70929 51383 70975
rect 51441 70929 51487 70975
rect 51545 70929 51591 70975
rect 51649 70929 51695 70975
rect 51753 70929 51799 70975
rect 51857 70929 51903 70975
rect 51961 70929 52007 70975
rect 52065 70929 52111 70975
rect 52169 70929 52215 70975
rect 52273 70929 52319 70975
rect 52377 70929 52423 70975
rect 52481 70929 52527 70975
rect 52585 70929 52631 70975
rect 52689 70929 52735 70975
rect 52793 70929 52839 70975
rect 52897 70929 52943 70975
rect 53001 70929 53047 70975
rect 53105 70929 53151 70975
rect 53209 70929 53255 70975
rect 53313 70929 53359 70975
rect 53417 70929 53463 70975
rect 53521 70929 53567 70975
rect 53625 70929 53671 70975
rect 53729 70929 53775 70975
rect 53833 70929 53879 70975
rect 53937 70929 53983 70975
rect 54041 70929 54087 70975
rect 54145 70929 54191 70975
rect 54249 70929 54295 70975
rect 54353 70929 54399 70975
rect 54457 70929 54503 70975
rect 54561 70929 54607 70975
rect 54665 70929 54711 70975
rect 54769 70929 54815 70975
rect 54873 70929 54919 70975
rect 54977 70929 55023 70975
rect 55081 70929 55127 70975
rect 55185 70929 55231 70975
rect 55289 70929 55335 70975
rect 55393 70929 55439 70975
rect 55497 70929 55543 70975
rect 55601 70929 55647 70975
rect 55705 70929 55751 70975
rect 55809 70929 55855 70975
rect 55913 70929 55959 70975
rect 56017 70929 56063 70975
rect 56121 70929 56167 70975
rect 56225 70929 56271 70975
rect 56329 70929 56375 70975
rect 56433 70929 56479 70975
rect 56537 70929 56583 70975
rect 56641 70929 56687 70975
rect 56745 70929 56791 70975
rect 56849 70929 56895 70975
rect 56953 70929 56999 70975
rect 57057 70929 57103 70975
rect 57161 70929 57207 70975
rect 57265 70929 57311 70975
rect 57369 70929 57415 70975
rect 57473 70929 57519 70975
rect 57577 70929 57623 70975
rect 57681 70929 57727 70975
rect 57785 70929 57831 70975
rect 57889 70929 57935 70975
rect 57993 70929 58039 70975
rect 58097 70929 58143 70975
rect 58201 70929 58247 70975
rect 58305 70929 58351 70975
rect 58409 70929 58455 70975
rect 58513 70929 58559 70975
rect 58617 70929 58663 70975
rect 58721 70929 58767 70975
rect 58825 70929 58871 70975
rect 58929 70929 58975 70975
rect 59033 70929 59079 70975
rect 59137 70929 59183 70975
rect 59241 70929 59287 70975
rect 59345 70929 59391 70975
rect 59449 70929 59495 70975
rect 59553 70929 59599 70975
rect 59657 70929 59703 70975
rect 59761 70929 59807 70975
rect 59865 70929 59911 70975
rect 59969 70929 60015 70975
rect 60073 70929 60119 70975
rect 60177 70929 60223 70975
rect 60281 70929 60327 70975
rect 60385 70929 60431 70975
rect 60489 70929 60535 70975
rect 60593 70929 60639 70975
rect 60697 70929 60743 70975
rect 60801 70929 60847 70975
rect 60905 70929 60951 70975
rect 61009 70929 61055 70975
rect 61113 70929 61159 70975
rect 61217 70929 61263 70975
rect 61321 70929 61367 70975
rect 61425 70929 61471 70975
rect 61529 70929 61575 70975
rect 61633 70929 61679 70975
rect 61737 70929 61783 70975
rect 61841 70929 61887 70975
rect 61945 70929 61991 70975
rect 62049 70929 62095 70975
rect 62153 70929 62199 70975
rect 62257 70929 62303 70975
rect 62361 70929 62407 70975
rect 62465 70929 62511 70975
rect 62569 70929 62615 70975
rect 62673 70929 62719 70975
rect 62777 70929 62823 70975
rect 62881 70929 62927 70975
rect 62985 70929 63031 70975
rect 63089 70929 63135 70975
rect 63193 70929 63239 70975
rect 63297 70929 63343 70975
rect 63401 70929 63447 70975
rect 63505 70929 63551 70975
rect 63609 70929 63655 70975
rect 63713 70929 63759 70975
rect 63817 70929 63863 70975
rect 63921 70929 63967 70975
rect 64025 70929 64071 70975
rect 64129 70929 64175 70975
rect 64233 70929 64279 70975
rect 64337 70929 64383 70975
rect 64441 70929 64487 70975
rect 64545 70929 64591 70975
rect 64649 70929 64695 70975
rect 64753 70929 64799 70975
rect 64857 70929 64903 70975
rect 64961 70929 65007 70975
rect 65065 70929 65111 70975
rect 65169 70929 65215 70975
rect 65273 70929 65319 70975
rect 65377 70929 65423 70975
rect 65481 70929 65527 70975
rect 65585 70929 65631 70975
rect 65689 70929 65735 70975
rect 65793 70929 65839 70975
rect 65897 70929 65943 70975
rect 66001 70929 66047 70975
rect 66105 70929 66151 70975
rect 66209 70929 66255 70975
rect 66313 70929 66359 70975
rect 66417 70929 66463 70975
rect 66521 70929 66567 70975
rect 66625 70929 66671 70975
rect 66729 70929 66775 70975
rect 66833 70929 66879 70975
rect 66937 70929 66983 70975
rect 67041 70929 67087 70975
rect 67145 70929 67191 70975
rect 67249 70929 67295 70975
rect 67353 70929 67399 70975
rect 67457 70929 67503 70975
rect 67561 70929 67607 70975
rect 67665 70929 67711 70975
rect 67769 70929 67815 70975
rect 67873 70929 67919 70975
rect 67977 70929 68023 70975
rect 68081 70929 68127 70975
rect 68185 70929 68231 70975
rect 68289 70929 68335 70975
rect 68393 70929 68439 70975
rect 68497 70929 68543 70975
rect 68601 70929 68647 70975
rect 68705 70929 68751 70975
rect 68809 70929 68855 70975
rect 68913 70929 68959 70975
rect 69017 70929 69063 70975
rect 69121 70929 69167 70975
rect 69225 70929 69271 70975
rect 69329 70929 69375 70975
rect 69433 70929 69479 70975
rect 69537 70929 69583 70975
rect 69641 70929 69687 70975
rect 69745 70929 69791 70975
rect 69849 70929 69895 70975
rect 13119 70825 13165 70871
rect 13223 70825 13269 70871
rect 13377 70825 13423 70871
rect 13481 70825 13527 70871
rect 13585 70825 13631 70871
rect 13689 70825 13735 70871
rect 13793 70825 13839 70871
rect 13897 70825 13943 70871
rect 14001 70825 14047 70871
rect 14105 70825 14151 70871
rect 14209 70825 14255 70871
rect 14313 70825 14359 70871
rect 14417 70825 14463 70871
rect 14521 70825 14567 70871
rect 14625 70825 14671 70871
rect 14729 70825 14775 70871
rect 14833 70825 14879 70871
rect 14937 70825 14983 70871
rect 15041 70825 15087 70871
rect 15145 70825 15191 70871
rect 15249 70825 15295 70871
rect 15353 70825 15399 70871
rect 15457 70825 15503 70871
rect 15561 70825 15607 70871
rect 15665 70825 15711 70871
rect 15769 70825 15815 70871
rect 15873 70825 15919 70871
rect 15977 70825 16023 70871
rect 16081 70825 16127 70871
rect 16185 70825 16231 70871
rect 16289 70825 16335 70871
rect 16393 70825 16439 70871
rect 16497 70825 16543 70871
rect 16601 70825 16647 70871
rect 16705 70825 16751 70871
rect 16809 70825 16855 70871
rect 16913 70825 16959 70871
rect 17017 70825 17063 70871
rect 17121 70825 17167 70871
rect 17225 70825 17271 70871
rect 17329 70825 17375 70871
rect 17433 70825 17479 70871
rect 17537 70825 17583 70871
rect 17641 70825 17687 70871
rect 17745 70825 17791 70871
rect 17849 70825 17895 70871
rect 17953 70825 17999 70871
rect 18057 70825 18103 70871
rect 18161 70825 18207 70871
rect 18265 70825 18311 70871
rect 18369 70825 18415 70871
rect 18473 70825 18519 70871
rect 18577 70825 18623 70871
rect 18681 70825 18727 70871
rect 18785 70825 18831 70871
rect 18889 70825 18935 70871
rect 18993 70825 19039 70871
rect 19097 70825 19143 70871
rect 19201 70825 19247 70871
rect 19305 70825 19351 70871
rect 19409 70825 19455 70871
rect 19513 70825 19559 70871
rect 19617 70825 19663 70871
rect 19721 70825 19767 70871
rect 19825 70825 19871 70871
rect 19929 70825 19975 70871
rect 20033 70825 20079 70871
rect 20137 70825 20183 70871
rect 20241 70825 20287 70871
rect 20345 70825 20391 70871
rect 20449 70825 20495 70871
rect 20553 70825 20599 70871
rect 20657 70825 20703 70871
rect 20761 70825 20807 70871
rect 20865 70825 20911 70871
rect 20969 70825 21015 70871
rect 21073 70825 21119 70871
rect 21177 70825 21223 70871
rect 21281 70825 21327 70871
rect 21385 70825 21431 70871
rect 21489 70825 21535 70871
rect 21593 70825 21639 70871
rect 21697 70825 21743 70871
rect 21801 70825 21847 70871
rect 21905 70825 21951 70871
rect 22009 70825 22055 70871
rect 22113 70825 22159 70871
rect 22217 70825 22263 70871
rect 22321 70825 22367 70871
rect 22425 70825 22471 70871
rect 22529 70825 22575 70871
rect 22633 70825 22679 70871
rect 22737 70825 22783 70871
rect 22841 70825 22887 70871
rect 22945 70825 22991 70871
rect 23049 70825 23095 70871
rect 23153 70825 23199 70871
rect 23257 70825 23303 70871
rect 23361 70825 23407 70871
rect 23465 70825 23511 70871
rect 23569 70825 23615 70871
rect 23673 70825 23719 70871
rect 23777 70825 23823 70871
rect 23881 70825 23927 70871
rect 23985 70825 24031 70871
rect 24089 70825 24135 70871
rect 24193 70825 24239 70871
rect 24297 70825 24343 70871
rect 24401 70825 24447 70871
rect 24505 70825 24551 70871
rect 24609 70825 24655 70871
rect 24713 70825 24759 70871
rect 24817 70825 24863 70871
rect 24921 70825 24967 70871
rect 25025 70825 25071 70871
rect 25129 70825 25175 70871
rect 25233 70825 25279 70871
rect 25337 70825 25383 70871
rect 25441 70825 25487 70871
rect 25545 70825 25591 70871
rect 25649 70825 25695 70871
rect 25753 70825 25799 70871
rect 25857 70825 25903 70871
rect 25961 70825 26007 70871
rect 26065 70825 26111 70871
rect 26169 70825 26215 70871
rect 26273 70825 26319 70871
rect 26377 70825 26423 70871
rect 26481 70825 26527 70871
rect 26585 70825 26631 70871
rect 26689 70825 26735 70871
rect 26793 70825 26839 70871
rect 26897 70825 26943 70871
rect 27001 70825 27047 70871
rect 27105 70825 27151 70871
rect 27209 70825 27255 70871
rect 27313 70825 27359 70871
rect 27417 70825 27463 70871
rect 27521 70825 27567 70871
rect 27625 70825 27671 70871
rect 27729 70825 27775 70871
rect 27833 70825 27879 70871
rect 27937 70825 27983 70871
rect 28041 70825 28087 70871
rect 28145 70825 28191 70871
rect 28249 70825 28295 70871
rect 28353 70825 28399 70871
rect 28457 70825 28503 70871
rect 28561 70825 28607 70871
rect 28665 70825 28711 70871
rect 28769 70825 28815 70871
rect 28873 70825 28919 70871
rect 28977 70825 29023 70871
rect 29081 70825 29127 70871
rect 29185 70825 29231 70871
rect 29289 70825 29335 70871
rect 29393 70825 29439 70871
rect 29497 70825 29543 70871
rect 29601 70825 29647 70871
rect 29705 70825 29751 70871
rect 29809 70825 29855 70871
rect 29913 70825 29959 70871
rect 30017 70825 30063 70871
rect 30121 70825 30167 70871
rect 30225 70825 30271 70871
rect 30329 70825 30375 70871
rect 30433 70825 30479 70871
rect 30537 70825 30583 70871
rect 30641 70825 30687 70871
rect 30745 70825 30791 70871
rect 30849 70825 30895 70871
rect 30953 70825 30999 70871
rect 31057 70825 31103 70871
rect 31161 70825 31207 70871
rect 31265 70825 31311 70871
rect 31369 70825 31415 70871
rect 31473 70825 31519 70871
rect 31577 70825 31623 70871
rect 31681 70825 31727 70871
rect 31785 70825 31831 70871
rect 31889 70825 31935 70871
rect 31993 70825 32039 70871
rect 32097 70825 32143 70871
rect 32201 70825 32247 70871
rect 32305 70825 32351 70871
rect 32409 70825 32455 70871
rect 32513 70825 32559 70871
rect 32617 70825 32663 70871
rect 32721 70825 32767 70871
rect 32825 70825 32871 70871
rect 32929 70825 32975 70871
rect 33033 70825 33079 70871
rect 33137 70825 33183 70871
rect 33241 70825 33287 70871
rect 33345 70825 33391 70871
rect 33449 70825 33495 70871
rect 33553 70825 33599 70871
rect 33657 70825 33703 70871
rect 33761 70825 33807 70871
rect 33865 70825 33911 70871
rect 33969 70825 34015 70871
rect 34073 70825 34119 70871
rect 34177 70825 34223 70871
rect 34281 70825 34327 70871
rect 34385 70825 34431 70871
rect 34489 70825 34535 70871
rect 34593 70825 34639 70871
rect 34697 70825 34743 70871
rect 34801 70825 34847 70871
rect 34905 70825 34951 70871
rect 35009 70825 35055 70871
rect 35113 70825 35159 70871
rect 35217 70825 35263 70871
rect 35321 70825 35367 70871
rect 35425 70825 35471 70871
rect 35529 70825 35575 70871
rect 35633 70825 35679 70871
rect 35737 70825 35783 70871
rect 35841 70825 35887 70871
rect 35945 70825 35991 70871
rect 36049 70825 36095 70871
rect 36153 70825 36199 70871
rect 36257 70825 36303 70871
rect 36361 70825 36407 70871
rect 36465 70825 36511 70871
rect 36569 70825 36615 70871
rect 36673 70825 36719 70871
rect 36777 70825 36823 70871
rect 36881 70825 36927 70871
rect 36985 70825 37031 70871
rect 37089 70825 37135 70871
rect 37193 70825 37239 70871
rect 37297 70825 37343 70871
rect 37401 70825 37447 70871
rect 37505 70825 37551 70871
rect 37609 70825 37655 70871
rect 37713 70825 37759 70871
rect 37817 70825 37863 70871
rect 37921 70825 37967 70871
rect 38025 70825 38071 70871
rect 38129 70825 38175 70871
rect 38233 70825 38279 70871
rect 38337 70825 38383 70871
rect 38441 70825 38487 70871
rect 38545 70825 38591 70871
rect 38649 70825 38695 70871
rect 38753 70825 38799 70871
rect 38857 70825 38903 70871
rect 38961 70825 39007 70871
rect 39065 70825 39111 70871
rect 39169 70825 39215 70871
rect 39273 70825 39319 70871
rect 39377 70825 39423 70871
rect 39481 70825 39527 70871
rect 39585 70825 39631 70871
rect 39689 70825 39735 70871
rect 39793 70825 39839 70871
rect 39897 70825 39943 70871
rect 40001 70825 40047 70871
rect 40105 70825 40151 70871
rect 40209 70825 40255 70871
rect 40313 70825 40359 70871
rect 40417 70825 40463 70871
rect 40521 70825 40567 70871
rect 40625 70825 40671 70871
rect 40729 70825 40775 70871
rect 40833 70825 40879 70871
rect 40937 70825 40983 70871
rect 41041 70825 41087 70871
rect 41145 70825 41191 70871
rect 41249 70825 41295 70871
rect 41353 70825 41399 70871
rect 41457 70825 41503 70871
rect 41561 70825 41607 70871
rect 41665 70825 41711 70871
rect 41769 70825 41815 70871
rect 41873 70825 41919 70871
rect 41977 70825 42023 70871
rect 42081 70825 42127 70871
rect 42185 70825 42231 70871
rect 42289 70825 42335 70871
rect 42393 70825 42439 70871
rect 42497 70825 42543 70871
rect 42601 70825 42647 70871
rect 42705 70825 42751 70871
rect 42809 70825 42855 70871
rect 42913 70825 42959 70871
rect 43017 70825 43063 70871
rect 43121 70825 43167 70871
rect 43225 70825 43271 70871
rect 43329 70825 43375 70871
rect 43433 70825 43479 70871
rect 43537 70825 43583 70871
rect 43641 70825 43687 70871
rect 43745 70825 43791 70871
rect 43849 70825 43895 70871
rect 43953 70825 43999 70871
rect 44057 70825 44103 70871
rect 44161 70825 44207 70871
rect 44265 70825 44311 70871
rect 44369 70825 44415 70871
rect 44473 70825 44519 70871
rect 44577 70825 44623 70871
rect 44681 70825 44727 70871
rect 44785 70825 44831 70871
rect 44889 70825 44935 70871
rect 44993 70825 45039 70871
rect 45097 70825 45143 70871
rect 45201 70825 45247 70871
rect 45305 70825 45351 70871
rect 45409 70825 45455 70871
rect 45513 70825 45559 70871
rect 45617 70825 45663 70871
rect 45721 70825 45767 70871
rect 45825 70825 45871 70871
rect 45929 70825 45975 70871
rect 46033 70825 46079 70871
rect 46137 70825 46183 70871
rect 46241 70825 46287 70871
rect 46345 70825 46391 70871
rect 46449 70825 46495 70871
rect 46553 70825 46599 70871
rect 46657 70825 46703 70871
rect 46761 70825 46807 70871
rect 46865 70825 46911 70871
rect 46969 70825 47015 70871
rect 47073 70825 47119 70871
rect 47177 70825 47223 70871
rect 47281 70825 47327 70871
rect 47385 70825 47431 70871
rect 47489 70825 47535 70871
rect 47593 70825 47639 70871
rect 47697 70825 47743 70871
rect 47801 70825 47847 70871
rect 47905 70825 47951 70871
rect 48009 70825 48055 70871
rect 48113 70825 48159 70871
rect 48217 70825 48263 70871
rect 48321 70825 48367 70871
rect 48425 70825 48471 70871
rect 48529 70825 48575 70871
rect 48633 70825 48679 70871
rect 48737 70825 48783 70871
rect 48841 70825 48887 70871
rect 48945 70825 48991 70871
rect 49049 70825 49095 70871
rect 49153 70825 49199 70871
rect 49257 70825 49303 70871
rect 49361 70825 49407 70871
rect 49465 70825 49511 70871
rect 49569 70825 49615 70871
rect 49673 70825 49719 70871
rect 49777 70825 49823 70871
rect 49881 70825 49927 70871
rect 49985 70825 50031 70871
rect 50089 70825 50135 70871
rect 50193 70825 50239 70871
rect 50297 70825 50343 70871
rect 50401 70825 50447 70871
rect 50505 70825 50551 70871
rect 50609 70825 50655 70871
rect 50713 70825 50759 70871
rect 50817 70825 50863 70871
rect 50921 70825 50967 70871
rect 51025 70825 51071 70871
rect 51129 70825 51175 70871
rect 51233 70825 51279 70871
rect 51337 70825 51383 70871
rect 51441 70825 51487 70871
rect 51545 70825 51591 70871
rect 51649 70825 51695 70871
rect 51753 70825 51799 70871
rect 51857 70825 51903 70871
rect 51961 70825 52007 70871
rect 52065 70825 52111 70871
rect 52169 70825 52215 70871
rect 52273 70825 52319 70871
rect 52377 70825 52423 70871
rect 52481 70825 52527 70871
rect 52585 70825 52631 70871
rect 52689 70825 52735 70871
rect 52793 70825 52839 70871
rect 52897 70825 52943 70871
rect 53001 70825 53047 70871
rect 53105 70825 53151 70871
rect 53209 70825 53255 70871
rect 53313 70825 53359 70871
rect 53417 70825 53463 70871
rect 53521 70825 53567 70871
rect 53625 70825 53671 70871
rect 53729 70825 53775 70871
rect 53833 70825 53879 70871
rect 53937 70825 53983 70871
rect 54041 70825 54087 70871
rect 54145 70825 54191 70871
rect 54249 70825 54295 70871
rect 54353 70825 54399 70871
rect 54457 70825 54503 70871
rect 54561 70825 54607 70871
rect 54665 70825 54711 70871
rect 54769 70825 54815 70871
rect 54873 70825 54919 70871
rect 54977 70825 55023 70871
rect 55081 70825 55127 70871
rect 55185 70825 55231 70871
rect 55289 70825 55335 70871
rect 55393 70825 55439 70871
rect 55497 70825 55543 70871
rect 55601 70825 55647 70871
rect 55705 70825 55751 70871
rect 55809 70825 55855 70871
rect 55913 70825 55959 70871
rect 56017 70825 56063 70871
rect 56121 70825 56167 70871
rect 56225 70825 56271 70871
rect 56329 70825 56375 70871
rect 56433 70825 56479 70871
rect 56537 70825 56583 70871
rect 56641 70825 56687 70871
rect 56745 70825 56791 70871
rect 56849 70825 56895 70871
rect 56953 70825 56999 70871
rect 57057 70825 57103 70871
rect 57161 70825 57207 70871
rect 57265 70825 57311 70871
rect 57369 70825 57415 70871
rect 57473 70825 57519 70871
rect 57577 70825 57623 70871
rect 57681 70825 57727 70871
rect 57785 70825 57831 70871
rect 57889 70825 57935 70871
rect 57993 70825 58039 70871
rect 58097 70825 58143 70871
rect 58201 70825 58247 70871
rect 58305 70825 58351 70871
rect 58409 70825 58455 70871
rect 58513 70825 58559 70871
rect 58617 70825 58663 70871
rect 58721 70825 58767 70871
rect 58825 70825 58871 70871
rect 58929 70825 58975 70871
rect 59033 70825 59079 70871
rect 59137 70825 59183 70871
rect 59241 70825 59287 70871
rect 59345 70825 59391 70871
rect 59449 70825 59495 70871
rect 59553 70825 59599 70871
rect 59657 70825 59703 70871
rect 59761 70825 59807 70871
rect 59865 70825 59911 70871
rect 59969 70825 60015 70871
rect 60073 70825 60119 70871
rect 60177 70825 60223 70871
rect 60281 70825 60327 70871
rect 60385 70825 60431 70871
rect 60489 70825 60535 70871
rect 60593 70825 60639 70871
rect 60697 70825 60743 70871
rect 60801 70825 60847 70871
rect 60905 70825 60951 70871
rect 61009 70825 61055 70871
rect 61113 70825 61159 70871
rect 61217 70825 61263 70871
rect 61321 70825 61367 70871
rect 61425 70825 61471 70871
rect 61529 70825 61575 70871
rect 61633 70825 61679 70871
rect 61737 70825 61783 70871
rect 61841 70825 61887 70871
rect 61945 70825 61991 70871
rect 62049 70825 62095 70871
rect 62153 70825 62199 70871
rect 62257 70825 62303 70871
rect 62361 70825 62407 70871
rect 62465 70825 62511 70871
rect 62569 70825 62615 70871
rect 62673 70825 62719 70871
rect 62777 70825 62823 70871
rect 62881 70825 62927 70871
rect 62985 70825 63031 70871
rect 63089 70825 63135 70871
rect 63193 70825 63239 70871
rect 63297 70825 63343 70871
rect 63401 70825 63447 70871
rect 63505 70825 63551 70871
rect 63609 70825 63655 70871
rect 63713 70825 63759 70871
rect 63817 70825 63863 70871
rect 63921 70825 63967 70871
rect 64025 70825 64071 70871
rect 64129 70825 64175 70871
rect 64233 70825 64279 70871
rect 64337 70825 64383 70871
rect 64441 70825 64487 70871
rect 64545 70825 64591 70871
rect 64649 70825 64695 70871
rect 64753 70825 64799 70871
rect 64857 70825 64903 70871
rect 64961 70825 65007 70871
rect 65065 70825 65111 70871
rect 65169 70825 65215 70871
rect 65273 70825 65319 70871
rect 65377 70825 65423 70871
rect 65481 70825 65527 70871
rect 65585 70825 65631 70871
rect 65689 70825 65735 70871
rect 65793 70825 65839 70871
rect 65897 70825 65943 70871
rect 66001 70825 66047 70871
rect 66105 70825 66151 70871
rect 66209 70825 66255 70871
rect 66313 70825 66359 70871
rect 66417 70825 66463 70871
rect 66521 70825 66567 70871
rect 66625 70825 66671 70871
rect 66729 70825 66775 70871
rect 66833 70825 66879 70871
rect 66937 70825 66983 70871
rect 67041 70825 67087 70871
rect 67145 70825 67191 70871
rect 67249 70825 67295 70871
rect 67353 70825 67399 70871
rect 67457 70825 67503 70871
rect 67561 70825 67607 70871
rect 67665 70825 67711 70871
rect 67769 70825 67815 70871
rect 67873 70825 67919 70871
rect 67977 70825 68023 70871
rect 68081 70825 68127 70871
rect 68185 70825 68231 70871
rect 68289 70825 68335 70871
rect 68393 70825 68439 70871
rect 68497 70825 68543 70871
rect 68601 70825 68647 70871
rect 68705 70825 68751 70871
rect 68809 70825 68855 70871
rect 68913 70825 68959 70871
rect 69017 70825 69063 70871
rect 69121 70825 69167 70871
rect 69225 70825 69271 70871
rect 69329 70825 69375 70871
rect 69433 70825 69479 70871
rect 69537 70825 69583 70871
rect 69641 70825 69687 70871
rect 69745 70825 69791 70871
rect 69849 70825 69895 70871
rect 13119 70721 13165 70767
rect 13223 70721 13269 70767
rect 13119 70617 13165 70663
rect 13223 70617 13269 70663
rect 13119 70513 13165 70559
rect 13223 70513 13269 70559
rect 13119 70409 13165 70455
rect 13223 70409 13269 70455
rect 13119 70305 13165 70351
rect 13223 70305 13269 70351
rect 13119 70201 13165 70247
rect 13223 70201 13269 70247
rect 13119 70097 13165 70143
rect 13223 70097 13269 70143
rect 13119 69993 13165 70039
rect 13223 69993 13269 70039
rect 13119 69889 13165 69935
rect 13223 69889 13269 69935
rect 13119 69785 13165 69831
rect 13223 69785 13269 69831
rect 69796 70674 69842 70720
rect 69900 70674 69946 70720
rect 69796 70570 69842 70616
rect 69900 70570 69946 70616
rect 69796 70466 69842 70512
rect 69900 70466 69946 70512
rect 69796 70362 69842 70408
rect 69900 70362 69946 70408
rect 69796 70258 69842 70304
rect 69900 70258 69946 70304
rect 69796 70154 69842 70200
rect 69900 70154 69946 70200
rect 69796 70050 69842 70096
rect 69900 70050 69946 70096
rect 69796 69900 69842 69946
rect 69900 69900 69946 69946
rect 70004 69900 70050 69946
rect 70108 69900 70154 69946
rect 70212 69900 70258 69946
rect 70316 69900 70362 69946
rect 70420 69900 70466 69946
rect 70524 69900 70570 69946
rect 70628 69900 70674 69946
rect 70824 69862 70870 69908
rect 70928 69862 70974 69908
rect 69796 69796 69842 69842
rect 69900 69796 69946 69842
rect 70004 69796 70050 69842
rect 70108 69796 70154 69842
rect 70212 69796 70258 69842
rect 70316 69796 70362 69842
rect 70420 69796 70466 69842
rect 70524 69796 70570 69842
rect 70628 69796 70674 69842
rect 13119 69681 13165 69727
rect 13223 69681 13269 69727
rect 13119 69577 13165 69623
rect 13223 69577 13269 69623
rect 13119 69473 13165 69519
rect 13223 69473 13269 69519
rect 13119 69369 13165 69415
rect 13223 69369 13269 69415
rect 13119 69265 13165 69311
rect 13223 69265 13269 69311
rect 13119 69161 13165 69207
rect 13223 69161 13269 69207
rect 13119 69057 13165 69103
rect 13223 69057 13269 69103
rect 13119 68953 13165 68999
rect 13223 68953 13269 68999
rect 13119 68849 13165 68895
rect 13223 68849 13269 68895
rect 13119 68745 13165 68791
rect 13223 68745 13269 68791
rect 13119 68641 13165 68687
rect 13223 68641 13269 68687
rect 13119 68537 13165 68583
rect 13223 68537 13269 68583
rect 13119 68433 13165 68479
rect 13223 68433 13269 68479
rect 13119 68329 13165 68375
rect 13223 68329 13269 68375
rect 13119 68225 13165 68271
rect 13223 68225 13269 68271
rect 13119 68121 13165 68167
rect 13223 68121 13269 68167
rect 13119 68017 13165 68063
rect 13223 68017 13269 68063
rect 13119 67913 13165 67959
rect 13223 67913 13269 67959
rect 13119 67809 13165 67855
rect 13223 67809 13269 67855
rect 13119 67705 13165 67751
rect 13223 67705 13269 67751
rect 13119 67601 13165 67647
rect 13223 67601 13269 67647
rect 13119 67497 13165 67543
rect 13223 67497 13269 67543
rect 13119 67393 13165 67439
rect 13223 67393 13269 67439
rect 13119 67289 13165 67335
rect 13223 67289 13269 67335
rect 13119 67185 13165 67231
rect 13223 67185 13269 67231
rect 13119 67081 13165 67127
rect 13223 67081 13269 67127
rect 13119 66977 13165 67023
rect 13223 66977 13269 67023
rect 13119 66873 13165 66919
rect 13223 66873 13269 66919
rect 13119 66769 13165 66815
rect 13223 66769 13269 66815
rect 13119 66665 13165 66711
rect 13223 66665 13269 66711
rect 13119 66561 13165 66607
rect 13223 66561 13269 66607
rect 13119 66457 13165 66503
rect 13223 66457 13269 66503
rect 13119 66353 13165 66399
rect 13223 66353 13269 66399
rect 13119 66249 13165 66295
rect 13223 66249 13269 66295
rect 13119 66145 13165 66191
rect 13223 66145 13269 66191
rect 13119 66041 13165 66087
rect 13223 66041 13269 66087
rect 13119 65937 13165 65983
rect 13223 65937 13269 65983
rect 13119 65833 13165 65879
rect 13223 65833 13269 65879
rect 13119 65729 13165 65775
rect 13223 65729 13269 65775
rect 13119 65625 13165 65671
rect 13223 65625 13269 65671
rect 13119 65521 13165 65567
rect 13223 65521 13269 65567
rect 13119 65417 13165 65463
rect 13223 65417 13269 65463
rect 13119 65313 13165 65359
rect 13223 65313 13269 65359
rect 13119 65209 13165 65255
rect 13223 65209 13269 65255
rect 13119 65105 13165 65151
rect 13223 65105 13269 65151
rect 13119 65001 13165 65047
rect 13223 65001 13269 65047
rect 13119 64897 13165 64943
rect 13223 64897 13269 64943
rect 13119 64793 13165 64839
rect 13223 64793 13269 64839
rect 13119 64689 13165 64735
rect 13223 64689 13269 64735
rect 13119 64585 13165 64631
rect 13223 64585 13269 64631
rect 13119 64481 13165 64527
rect 13223 64481 13269 64527
rect 13119 64377 13165 64423
rect 13223 64377 13269 64423
rect 13119 64273 13165 64319
rect 13223 64273 13269 64319
rect 13119 64169 13165 64215
rect 13223 64169 13269 64215
rect 13119 64065 13165 64111
rect 13223 64065 13269 64111
rect 13119 63961 13165 64007
rect 13223 63961 13269 64007
rect 13119 63857 13165 63903
rect 13223 63857 13269 63903
rect 13119 63753 13165 63799
rect 13223 63753 13269 63799
rect 13119 63649 13165 63695
rect 13223 63649 13269 63695
rect 13119 63545 13165 63591
rect 13223 63545 13269 63591
rect 13119 63441 13165 63487
rect 13223 63441 13269 63487
rect 13119 63337 13165 63383
rect 13223 63337 13269 63383
rect 13119 63233 13165 63279
rect 13223 63233 13269 63279
rect 13119 63129 13165 63175
rect 13223 63129 13269 63175
rect 13119 63025 13165 63071
rect 13223 63025 13269 63071
rect 13119 62921 13165 62967
rect 13223 62921 13269 62967
rect 13119 62817 13165 62863
rect 13223 62817 13269 62863
rect 13119 62713 13165 62759
rect 13223 62713 13269 62759
rect 13119 62609 13165 62655
rect 13223 62609 13269 62655
rect 13119 62505 13165 62551
rect 13223 62505 13269 62551
rect 13119 62401 13165 62447
rect 13223 62401 13269 62447
rect 13119 62297 13165 62343
rect 13223 62297 13269 62343
rect 13119 62193 13165 62239
rect 13223 62193 13269 62239
rect 13119 62089 13165 62135
rect 13223 62089 13269 62135
rect 13119 61985 13165 62031
rect 13223 61985 13269 62031
rect 13119 61881 13165 61927
rect 13223 61881 13269 61927
rect 13119 61777 13165 61823
rect 13223 61777 13269 61823
rect 13119 61673 13165 61719
rect 13223 61673 13269 61719
rect 13119 61569 13165 61615
rect 13223 61569 13269 61615
rect 13119 61465 13165 61511
rect 13223 61465 13269 61511
rect 13119 61361 13165 61407
rect 13223 61361 13269 61407
rect 13119 61257 13165 61303
rect 13223 61257 13269 61303
rect 13119 61153 13165 61199
rect 13223 61153 13269 61199
rect 13119 61049 13165 61095
rect 13223 61049 13269 61095
rect 13119 60945 13165 60991
rect 13223 60945 13269 60991
rect 13119 60841 13165 60887
rect 13223 60841 13269 60887
rect 13119 60737 13165 60783
rect 13223 60737 13269 60783
rect 13119 60633 13165 60679
rect 13223 60633 13269 60679
rect 13119 60529 13165 60575
rect 13223 60529 13269 60575
rect 13119 60425 13165 60471
rect 13223 60425 13269 60471
rect 13119 60321 13165 60367
rect 13223 60321 13269 60367
rect 13119 60217 13165 60263
rect 13223 60217 13269 60263
rect 13119 60113 13165 60159
rect 13223 60113 13269 60159
rect 13119 60009 13165 60055
rect 13223 60009 13269 60055
rect 13119 59905 13165 59951
rect 13223 59905 13269 59951
rect 13119 59801 13165 59847
rect 13223 59801 13269 59847
rect 13119 59697 13165 59743
rect 13223 59697 13269 59743
rect 13119 59593 13165 59639
rect 13223 59593 13269 59639
rect 13119 59489 13165 59535
rect 13223 59489 13269 59535
rect 13119 59385 13165 59431
rect 13223 59385 13269 59431
rect 13119 59281 13165 59327
rect 13223 59281 13269 59327
rect 13119 59177 13165 59223
rect 13223 59177 13269 59223
rect 13119 59073 13165 59119
rect 13223 59073 13269 59119
rect 13119 58969 13165 59015
rect 13223 58969 13269 59015
rect 13119 58865 13165 58911
rect 13223 58865 13269 58911
rect 13119 58761 13165 58807
rect 13223 58761 13269 58807
rect 13119 58657 13165 58703
rect 13223 58657 13269 58703
rect 13119 58553 13165 58599
rect 13223 58553 13269 58599
rect 13119 58449 13165 58495
rect 13223 58449 13269 58495
rect 13119 58345 13165 58391
rect 13223 58345 13269 58391
rect 13119 58241 13165 58287
rect 13223 58241 13269 58287
rect 13119 58137 13165 58183
rect 13223 58137 13269 58183
rect 13119 58033 13165 58079
rect 13223 58033 13269 58079
rect 13119 57929 13165 57975
rect 13223 57929 13269 57975
rect 13119 57825 13165 57871
rect 13223 57825 13269 57871
rect 13119 57721 13165 57767
rect 13223 57721 13269 57767
rect 13119 57617 13165 57663
rect 13223 57617 13269 57663
rect 13119 57513 13165 57559
rect 13223 57513 13269 57559
rect 13119 57409 13165 57455
rect 13223 57409 13269 57455
rect 13119 57305 13165 57351
rect 13223 57305 13269 57351
rect 13119 57201 13165 57247
rect 13223 57201 13269 57247
rect 13119 57097 13165 57143
rect 13223 57097 13269 57143
rect 13119 56993 13165 57039
rect 13223 56993 13269 57039
rect 13119 56889 13165 56935
rect 13223 56889 13269 56935
rect 13119 56785 13165 56831
rect 13223 56785 13269 56831
rect 13119 56681 13165 56727
rect 13223 56681 13269 56727
rect 13119 56577 13165 56623
rect 13223 56577 13269 56623
rect 13119 56473 13165 56519
rect 13223 56473 13269 56519
rect 13119 56369 13165 56415
rect 13223 56369 13269 56415
rect 13119 56265 13165 56311
rect 13223 56265 13269 56311
rect 13119 56161 13165 56207
rect 13223 56161 13269 56207
rect 13119 56057 13165 56103
rect 13223 56057 13269 56103
rect 13119 55953 13165 55999
rect 13223 55953 13269 55999
rect 13119 55849 13165 55895
rect 13223 55849 13269 55895
rect 13119 55745 13165 55791
rect 13223 55745 13269 55791
rect 13119 55641 13165 55687
rect 13223 55641 13269 55687
rect 13119 55537 13165 55583
rect 13223 55537 13269 55583
rect 13119 55433 13165 55479
rect 13223 55433 13269 55479
rect 13119 55329 13165 55375
rect 13223 55329 13269 55375
rect 13119 55225 13165 55271
rect 13223 55225 13269 55271
rect 13119 55121 13165 55167
rect 13223 55121 13269 55167
rect 13119 55017 13165 55063
rect 13223 55017 13269 55063
rect 13119 54913 13165 54959
rect 13223 54913 13269 54959
rect 13119 54809 13165 54855
rect 13223 54809 13269 54855
rect 13119 54705 13165 54751
rect 13223 54705 13269 54751
rect 13119 54601 13165 54647
rect 13223 54601 13269 54647
rect 13119 54497 13165 54543
rect 13223 54497 13269 54543
rect 13119 54393 13165 54439
rect 13223 54393 13269 54439
rect 13119 54289 13165 54335
rect 13223 54289 13269 54335
rect 13119 54185 13165 54231
rect 13223 54185 13269 54231
rect 13119 54081 13165 54127
rect 13223 54081 13269 54127
rect 13119 53977 13165 54023
rect 13223 53977 13269 54023
rect 13119 53873 13165 53919
rect 13223 53873 13269 53919
rect 13119 53769 13165 53815
rect 13223 53769 13269 53815
rect 13119 53665 13165 53711
rect 13223 53665 13269 53711
rect 13119 53561 13165 53607
rect 13223 53561 13269 53607
rect 13119 53457 13165 53503
rect 13223 53457 13269 53503
rect 13119 53353 13165 53399
rect 13223 53353 13269 53399
rect 13119 53249 13165 53295
rect 13223 53249 13269 53295
rect 13119 53145 13165 53191
rect 13223 53145 13269 53191
rect 13119 53041 13165 53087
rect 13223 53041 13269 53087
rect 13119 52937 13165 52983
rect 13223 52937 13269 52983
rect 13119 52833 13165 52879
rect 13223 52833 13269 52879
rect 13119 52729 13165 52775
rect 13223 52729 13269 52775
rect 13119 52625 13165 52671
rect 13223 52625 13269 52671
rect 13119 52521 13165 52567
rect 13223 52521 13269 52567
rect 13119 52417 13165 52463
rect 13223 52417 13269 52463
rect 13119 52313 13165 52359
rect 13223 52313 13269 52359
rect 13119 52209 13165 52255
rect 13223 52209 13269 52255
rect 13119 52105 13165 52151
rect 13223 52105 13269 52151
rect 13119 52001 13165 52047
rect 13223 52001 13269 52047
rect 13119 51897 13165 51943
rect 13223 51897 13269 51943
rect 13119 51793 13165 51839
rect 13223 51793 13269 51839
rect 13119 51689 13165 51735
rect 13223 51689 13269 51735
rect 13119 51585 13165 51631
rect 13223 51585 13269 51631
rect 13119 51481 13165 51527
rect 13223 51481 13269 51527
rect 13119 51377 13165 51423
rect 13223 51377 13269 51423
rect 13119 51273 13165 51319
rect 13223 51273 13269 51319
rect 13119 51169 13165 51215
rect 13223 51169 13269 51215
rect 13119 51065 13165 51111
rect 13223 51065 13269 51111
rect 13119 50961 13165 51007
rect 13223 50961 13269 51007
rect 13119 50857 13165 50903
rect 13223 50857 13269 50903
rect 13119 50753 13165 50799
rect 13223 50753 13269 50799
rect 13119 50649 13165 50695
rect 13223 50649 13269 50695
rect 13119 50545 13165 50591
rect 13223 50545 13269 50591
rect 13119 50441 13165 50487
rect 13223 50441 13269 50487
rect 13119 50337 13165 50383
rect 13223 50337 13269 50383
rect 13119 50233 13165 50279
rect 13223 50233 13269 50279
rect 13119 50129 13165 50175
rect 13223 50129 13269 50175
rect 13119 50025 13165 50071
rect 13223 50025 13269 50071
rect 13119 49921 13165 49967
rect 13223 49921 13269 49967
rect 13119 49817 13165 49863
rect 13223 49817 13269 49863
rect 13119 49713 13165 49759
rect 13223 49713 13269 49759
rect 13119 49609 13165 49655
rect 13223 49609 13269 49655
rect 13119 49505 13165 49551
rect 13223 49505 13269 49551
rect 13119 49401 13165 49447
rect 13223 49401 13269 49447
rect 13119 49297 13165 49343
rect 13223 49297 13269 49343
rect 13119 49193 13165 49239
rect 13223 49193 13269 49239
rect 13119 49089 13165 49135
rect 13223 49089 13269 49135
rect 13119 48985 13165 49031
rect 13223 48985 13269 49031
rect 13119 48881 13165 48927
rect 13223 48881 13269 48927
rect 13119 48777 13165 48823
rect 13223 48777 13269 48823
rect 13119 48673 13165 48719
rect 13223 48673 13269 48719
rect 13119 48569 13165 48615
rect 13223 48569 13269 48615
rect 13119 48465 13165 48511
rect 13223 48465 13269 48511
rect 13119 48361 13165 48407
rect 13223 48361 13269 48407
rect 13119 48257 13165 48303
rect 13223 48257 13269 48303
rect 13119 48153 13165 48199
rect 13223 48153 13269 48199
rect 13119 48049 13165 48095
rect 13223 48049 13269 48095
rect 13119 47945 13165 47991
rect 13223 47945 13269 47991
rect 13119 47841 13165 47887
rect 13223 47841 13269 47887
rect 13119 47737 13165 47783
rect 13223 47737 13269 47783
rect 13119 47633 13165 47679
rect 13223 47633 13269 47679
rect 13119 47529 13165 47575
rect 13223 47529 13269 47575
rect 13119 47425 13165 47471
rect 13223 47425 13269 47471
rect 13119 47321 13165 47367
rect 13223 47321 13269 47367
rect 13119 47217 13165 47263
rect 13223 47217 13269 47263
rect 13119 47113 13165 47159
rect 13223 47113 13269 47159
rect 13119 47009 13165 47055
rect 13223 47009 13269 47055
rect 13119 46905 13165 46951
rect 13223 46905 13269 46951
rect 13119 46801 13165 46847
rect 13223 46801 13269 46847
rect 13119 46697 13165 46743
rect 13223 46697 13269 46743
rect 13119 46593 13165 46639
rect 13223 46593 13269 46639
rect 13119 46489 13165 46535
rect 13223 46489 13269 46535
rect 13119 46385 13165 46431
rect 13223 46385 13269 46431
rect 13119 46281 13165 46327
rect 13223 46281 13269 46327
rect 13119 46177 13165 46223
rect 13223 46177 13269 46223
rect 13119 46073 13165 46119
rect 13223 46073 13269 46119
rect 13119 45969 13165 46015
rect 13223 45969 13269 46015
rect 13119 45865 13165 45911
rect 13223 45865 13269 45911
rect 13119 45761 13165 45807
rect 13223 45761 13269 45807
rect 13119 45657 13165 45703
rect 13223 45657 13269 45703
rect 13119 45553 13165 45599
rect 13223 45553 13269 45599
rect 13119 45449 13165 45495
rect 13223 45449 13269 45495
rect 13119 45345 13165 45391
rect 13223 45345 13269 45391
rect 13119 45241 13165 45287
rect 13223 45241 13269 45287
rect 13119 45137 13165 45183
rect 13223 45137 13269 45183
rect 13119 45033 13165 45079
rect 13223 45033 13269 45079
rect 70824 69758 70870 69804
rect 70928 69758 70974 69804
rect 70824 69654 70870 69700
rect 70928 69654 70974 69700
rect 70824 69550 70870 69596
rect 70928 69550 70974 69596
rect 70824 69446 70870 69492
rect 70928 69446 70974 69492
rect 70824 69342 70870 69388
rect 70928 69342 70974 69388
rect 70824 69238 70870 69284
rect 70928 69238 70974 69284
rect 70824 69134 70870 69180
rect 70928 69134 70974 69180
rect 70824 69030 70870 69076
rect 70928 69030 70974 69076
rect 70824 68926 70870 68972
rect 70928 68926 70974 68972
rect 70824 68822 70870 68868
rect 70928 68822 70974 68868
rect 70824 68718 70870 68764
rect 70928 68718 70974 68764
rect 70824 68614 70870 68660
rect 70928 68614 70974 68660
rect 70824 68510 70870 68556
rect 70928 68510 70974 68556
rect 70824 68406 70870 68452
rect 70928 68406 70974 68452
rect 70824 68302 70870 68348
rect 70928 68302 70974 68348
rect 70824 68198 70870 68244
rect 70928 68198 70974 68244
rect 70824 68094 70870 68140
rect 70928 68094 70974 68140
rect 70824 67990 70870 68036
rect 70928 67990 70974 68036
rect 70824 67886 70870 67932
rect 70928 67886 70974 67932
rect 70824 67782 70870 67828
rect 70928 67782 70974 67828
rect 70824 67678 70870 67724
rect 70928 67678 70974 67724
rect 70824 67574 70870 67620
rect 70928 67574 70974 67620
rect 70824 67470 70870 67516
rect 70928 67470 70974 67516
rect 70824 67366 70870 67412
rect 70928 67366 70974 67412
rect 70824 67262 70870 67308
rect 70928 67262 70974 67308
rect 70824 67158 70870 67204
rect 70928 67158 70974 67204
rect 70824 67054 70870 67100
rect 70928 67054 70974 67100
rect 70824 66950 70870 66996
rect 70928 66950 70974 66996
rect 70824 66846 70870 66892
rect 70928 66846 70974 66892
rect 70824 66742 70870 66788
rect 70928 66742 70974 66788
rect 70824 66638 70870 66684
rect 70928 66638 70974 66684
rect 70824 66534 70870 66580
rect 70928 66534 70974 66580
rect 70824 66430 70870 66476
rect 70928 66430 70974 66476
rect 70824 66326 70870 66372
rect 70928 66326 70974 66372
rect 70824 66222 70870 66268
rect 70928 66222 70974 66268
rect 70824 66118 70870 66164
rect 70928 66118 70974 66164
rect 70824 66014 70870 66060
rect 70928 66014 70974 66060
rect 70824 65910 70870 65956
rect 70928 65910 70974 65956
rect 70824 65806 70870 65852
rect 70928 65806 70974 65852
rect 70824 65702 70870 65748
rect 70928 65702 70974 65748
rect 70824 65598 70870 65644
rect 70928 65598 70974 65644
rect 70824 65494 70870 65540
rect 70928 65494 70974 65540
rect 70824 65390 70870 65436
rect 70928 65390 70974 65436
rect 70824 65286 70870 65332
rect 70928 65286 70974 65332
rect 70824 65182 70870 65228
rect 70928 65182 70974 65228
rect 70824 65078 70870 65124
rect 70928 65078 70974 65124
rect 70824 64974 70870 65020
rect 70928 64974 70974 65020
rect 70824 64870 70870 64916
rect 70928 64870 70974 64916
rect 70824 64766 70870 64812
rect 70928 64766 70974 64812
rect 70824 64662 70870 64708
rect 70928 64662 70974 64708
rect 70824 64558 70870 64604
rect 70928 64558 70974 64604
rect 70824 64454 70870 64500
rect 70928 64454 70974 64500
rect 70824 64350 70870 64396
rect 70928 64350 70974 64396
rect 70824 64246 70870 64292
rect 70928 64246 70974 64292
rect 70824 64142 70870 64188
rect 70928 64142 70974 64188
rect 70824 64038 70870 64084
rect 70928 64038 70974 64084
rect 70824 63934 70870 63980
rect 70928 63934 70974 63980
rect 70824 63830 70870 63876
rect 70928 63830 70974 63876
rect 70824 63726 70870 63772
rect 70928 63726 70974 63772
rect 70824 63622 70870 63668
rect 70928 63622 70974 63668
rect 70824 63518 70870 63564
rect 70928 63518 70974 63564
rect 70824 63414 70870 63460
rect 70928 63414 70974 63460
rect 70824 63310 70870 63356
rect 70928 63310 70974 63356
rect 70824 63206 70870 63252
rect 70928 63206 70974 63252
rect 70824 63102 70870 63148
rect 70928 63102 70974 63148
rect 70824 62998 70870 63044
rect 70928 62998 70974 63044
rect 70824 62894 70870 62940
rect 70928 62894 70974 62940
rect 70824 62790 70870 62836
rect 70928 62790 70974 62836
rect 70824 62686 70870 62732
rect 70928 62686 70974 62732
rect 70824 62582 70870 62628
rect 70928 62582 70974 62628
rect 70824 62478 70870 62524
rect 70928 62478 70974 62524
rect 70824 62374 70870 62420
rect 70928 62374 70974 62420
rect 70824 62270 70870 62316
rect 70928 62270 70974 62316
rect 70824 62166 70870 62212
rect 70928 62166 70974 62212
rect 70824 62062 70870 62108
rect 70928 62062 70974 62108
rect 70824 61958 70870 62004
rect 70928 61958 70974 62004
rect 70824 61854 70870 61900
rect 70928 61854 70974 61900
rect 70824 61750 70870 61796
rect 70928 61750 70974 61796
rect 70824 61646 70870 61692
rect 70928 61646 70974 61692
rect 70824 61542 70870 61588
rect 70928 61542 70974 61588
rect 70824 61438 70870 61484
rect 70928 61438 70974 61484
rect 70824 61334 70870 61380
rect 70928 61334 70974 61380
rect 70824 61230 70870 61276
rect 70928 61230 70974 61276
rect 70824 61126 70870 61172
rect 70928 61126 70974 61172
rect 70824 61022 70870 61068
rect 70928 61022 70974 61068
rect 70824 60918 70870 60964
rect 70928 60918 70974 60964
rect 70824 60814 70870 60860
rect 70928 60814 70974 60860
rect 70824 60710 70870 60756
rect 70928 60710 70974 60756
rect 70824 60606 70870 60652
rect 70928 60606 70974 60652
rect 70824 60502 70870 60548
rect 70928 60502 70974 60548
rect 70824 60398 70870 60444
rect 70928 60398 70974 60444
rect 70824 60294 70870 60340
rect 70928 60294 70974 60340
rect 70824 60190 70870 60236
rect 70928 60190 70974 60236
rect 70824 60086 70870 60132
rect 70928 60086 70974 60132
rect 70824 59982 70870 60028
rect 70928 59982 70974 60028
rect 70824 59878 70870 59924
rect 70928 59878 70974 59924
rect 70824 59774 70870 59820
rect 70928 59774 70974 59820
rect 70824 59670 70870 59716
rect 70928 59670 70974 59716
rect 70824 59566 70870 59612
rect 70928 59566 70974 59612
rect 70824 59462 70870 59508
rect 70928 59462 70974 59508
rect 70824 59358 70870 59404
rect 70928 59358 70974 59404
rect 70824 59254 70870 59300
rect 70928 59254 70974 59300
rect 70824 59150 70870 59196
rect 70928 59150 70974 59196
rect 70824 59046 70870 59092
rect 70928 59046 70974 59092
rect 70824 58942 70870 58988
rect 70928 58942 70974 58988
rect 70824 58838 70870 58884
rect 70928 58838 70974 58884
rect 70824 58734 70870 58780
rect 70928 58734 70974 58780
rect 70824 58630 70870 58676
rect 70928 58630 70974 58676
rect 70824 58526 70870 58572
rect 70928 58526 70974 58572
rect 70824 58422 70870 58468
rect 70928 58422 70974 58468
rect 70824 58318 70870 58364
rect 70928 58318 70974 58364
rect 70824 58214 70870 58260
rect 70928 58214 70974 58260
rect 70824 58110 70870 58156
rect 70928 58110 70974 58156
rect 70824 58006 70870 58052
rect 70928 58006 70974 58052
rect 70824 57902 70870 57948
rect 70928 57902 70974 57948
rect 70824 57798 70870 57844
rect 70928 57798 70974 57844
rect 70824 57694 70870 57740
rect 70928 57694 70974 57740
rect 70824 57590 70870 57636
rect 70928 57590 70974 57636
rect 70824 57486 70870 57532
rect 70928 57486 70974 57532
rect 70824 57382 70870 57428
rect 70928 57382 70974 57428
rect 70824 57278 70870 57324
rect 70928 57278 70974 57324
rect 70824 57174 70870 57220
rect 70928 57174 70974 57220
rect 70824 57070 70870 57116
rect 70928 57070 70974 57116
rect 70824 56966 70870 57012
rect 70928 56966 70974 57012
rect 70824 56862 70870 56908
rect 70928 56862 70974 56908
rect 70824 56758 70870 56804
rect 70928 56758 70974 56804
rect 70824 56654 70870 56700
rect 70928 56654 70974 56700
rect 70824 56550 70870 56596
rect 70928 56550 70974 56596
rect 70824 56446 70870 56492
rect 70928 56446 70974 56492
rect 70824 56342 70870 56388
rect 70928 56342 70974 56388
rect 70824 56238 70870 56284
rect 70928 56238 70974 56284
rect 70824 56134 70870 56180
rect 70928 56134 70974 56180
rect 70824 56030 70870 56076
rect 70928 56030 70974 56076
rect 70824 55926 70870 55972
rect 70928 55926 70974 55972
rect 70824 55822 70870 55868
rect 70928 55822 70974 55868
rect 70824 55718 70870 55764
rect 70928 55718 70974 55764
rect 70824 55614 70870 55660
rect 70928 55614 70974 55660
rect 70824 55510 70870 55556
rect 70928 55510 70974 55556
rect 70824 55406 70870 55452
rect 70928 55406 70974 55452
rect 70824 55302 70870 55348
rect 70928 55302 70974 55348
rect 70824 55198 70870 55244
rect 70928 55198 70974 55244
rect 70824 55094 70870 55140
rect 70928 55094 70974 55140
rect 70824 54990 70870 55036
rect 70928 54990 70974 55036
rect 70824 54886 70870 54932
rect 70928 54886 70974 54932
rect 70824 54782 70870 54828
rect 70928 54782 70974 54828
rect 70824 54678 70870 54724
rect 70928 54678 70974 54724
rect 70824 54574 70870 54620
rect 70928 54574 70974 54620
rect 70824 54470 70870 54516
rect 70928 54470 70974 54516
rect 70824 54366 70870 54412
rect 70928 54366 70974 54412
rect 70824 54262 70870 54308
rect 70928 54262 70974 54308
rect 70824 54158 70870 54204
rect 70928 54158 70974 54204
rect 70824 54054 70870 54100
rect 70928 54054 70974 54100
rect 70824 53950 70870 53996
rect 70928 53950 70974 53996
rect 70824 53846 70870 53892
rect 70928 53846 70974 53892
rect 70824 53742 70870 53788
rect 70928 53742 70974 53788
rect 70824 53638 70870 53684
rect 70928 53638 70974 53684
rect 70824 53534 70870 53580
rect 70928 53534 70974 53580
rect 70824 53430 70870 53476
rect 70928 53430 70974 53476
rect 70824 53326 70870 53372
rect 70928 53326 70974 53372
rect 70824 53222 70870 53268
rect 70928 53222 70974 53268
rect 70824 53118 70870 53164
rect 70928 53118 70974 53164
rect 70824 53014 70870 53060
rect 70928 53014 70974 53060
rect 70824 52910 70870 52956
rect 70928 52910 70974 52956
rect 70824 52806 70870 52852
rect 70928 52806 70974 52852
rect 70824 52702 70870 52748
rect 70928 52702 70974 52748
rect 70824 52598 70870 52644
rect 70928 52598 70974 52644
rect 70824 52494 70870 52540
rect 70928 52494 70974 52540
rect 70824 52390 70870 52436
rect 70928 52390 70974 52436
rect 70824 52286 70870 52332
rect 70928 52286 70974 52332
rect 70824 52182 70870 52228
rect 70928 52182 70974 52228
rect 70824 52078 70870 52124
rect 70928 52078 70974 52124
rect 70824 51974 70870 52020
rect 70928 51974 70974 52020
rect 70824 51870 70870 51916
rect 70928 51870 70974 51916
rect 70824 51766 70870 51812
rect 70928 51766 70974 51812
rect 70824 51662 70870 51708
rect 70928 51662 70974 51708
rect 70824 51558 70870 51604
rect 70928 51558 70974 51604
rect 70824 51454 70870 51500
rect 70928 51454 70974 51500
rect 70824 51350 70870 51396
rect 70928 51350 70974 51396
rect 70824 51246 70870 51292
rect 70928 51246 70974 51292
rect 70824 51142 70870 51188
rect 70928 51142 70974 51188
rect 70824 51038 70870 51084
rect 70928 51038 70974 51084
rect 70824 50934 70870 50980
rect 70928 50934 70974 50980
rect 70824 50830 70870 50876
rect 70928 50830 70974 50876
rect 70824 50726 70870 50772
rect 70928 50726 70974 50772
rect 70824 50622 70870 50668
rect 70928 50622 70974 50668
rect 70824 50518 70870 50564
rect 70928 50518 70974 50564
rect 70824 50414 70870 50460
rect 70928 50414 70974 50460
rect 70824 50310 70870 50356
rect 70928 50310 70974 50356
rect 70824 50206 70870 50252
rect 70928 50206 70974 50252
rect 70824 50102 70870 50148
rect 70928 50102 70974 50148
rect 70824 49998 70870 50044
rect 70928 49998 70974 50044
rect 70824 49894 70870 49940
rect 70928 49894 70974 49940
rect 70824 49790 70870 49836
rect 70928 49790 70974 49836
rect 70824 49686 70870 49732
rect 70928 49686 70974 49732
rect 70824 49582 70870 49628
rect 70928 49582 70974 49628
rect 70824 49478 70870 49524
rect 70928 49478 70974 49524
rect 70824 49374 70870 49420
rect 70928 49374 70974 49420
rect 70824 49270 70870 49316
rect 70928 49270 70974 49316
rect 70824 49166 70870 49212
rect 70928 49166 70974 49212
rect 70824 49062 70870 49108
rect 70928 49062 70974 49108
rect 70824 48958 70870 49004
rect 70928 48958 70974 49004
rect 70824 48854 70870 48900
rect 70928 48854 70974 48900
rect 70824 48750 70870 48796
rect 70928 48750 70974 48796
rect 70824 48646 70870 48692
rect 70928 48646 70974 48692
rect 70824 48542 70870 48588
rect 70928 48542 70974 48588
rect 70824 48438 70870 48484
rect 70928 48438 70974 48484
rect 70824 48334 70870 48380
rect 70928 48334 70974 48380
rect 70824 48230 70870 48276
rect 70928 48230 70974 48276
rect 70824 48126 70870 48172
rect 70928 48126 70974 48172
rect 70824 48022 70870 48068
rect 70928 48022 70974 48068
rect 70824 47918 70870 47964
rect 70928 47918 70974 47964
rect 70824 47814 70870 47860
rect 70928 47814 70974 47860
rect 70824 47710 70870 47756
rect 70928 47710 70974 47756
rect 70824 47606 70870 47652
rect 70928 47606 70974 47652
rect 70824 47502 70870 47548
rect 70928 47502 70974 47548
rect 70824 47398 70870 47444
rect 70928 47398 70974 47444
rect 70824 47294 70870 47340
rect 70928 47294 70974 47340
rect 70824 47190 70870 47236
rect 70928 47190 70974 47236
rect 70824 47086 70870 47132
rect 70928 47086 70974 47132
rect 70824 46982 70870 47028
rect 70928 46982 70974 47028
rect 70824 46878 70870 46924
rect 70928 46878 70974 46924
rect 70824 46774 70870 46820
rect 70928 46774 70974 46820
rect 70824 46670 70870 46716
rect 70928 46670 70974 46716
rect 70824 46566 70870 46612
rect 70928 46566 70974 46612
rect 70824 46462 70870 46508
rect 70928 46462 70974 46508
rect 70824 46358 70870 46404
rect 70928 46358 70974 46404
rect 70824 46254 70870 46300
rect 70928 46254 70974 46300
rect 70824 46150 70870 46196
rect 70928 46150 70974 46196
rect 70824 46046 70870 46092
rect 70928 46046 70974 46092
rect 70824 45942 70870 45988
rect 70928 45942 70974 45988
rect 70824 45838 70870 45884
rect 70928 45838 70974 45884
rect 70824 45734 70870 45780
rect 70928 45734 70974 45780
rect 70824 45630 70870 45676
rect 70928 45630 70974 45676
rect 70824 45526 70870 45572
rect 70928 45526 70974 45572
rect 70824 45422 70870 45468
rect 70928 45422 70974 45468
rect 70824 45318 70870 45364
rect 70928 45318 70974 45364
rect 70824 45214 70870 45260
rect 70928 45214 70974 45260
rect 70824 45110 70870 45156
rect 70928 45110 70974 45156
rect 70824 45006 70870 45052
rect 70928 45006 70974 45052
rect 70824 44902 70870 44948
rect 70928 44902 70974 44948
rect 13254 44778 13300 44824
rect 70824 44798 70870 44844
rect 70928 44798 70974 44844
rect 13386 44646 13432 44692
rect 70824 44694 70870 44740
rect 70928 44694 70974 44740
rect 70824 44590 70870 44636
rect 70928 44590 70974 44636
rect 13518 44514 13564 44560
rect 70824 44486 70870 44532
rect 70928 44486 70974 44532
rect 13650 44382 13696 44428
rect 70824 44382 70870 44428
rect 70928 44382 70974 44428
rect 13782 44250 13828 44296
rect 70824 44278 70870 44324
rect 70928 44278 70974 44324
rect 13914 44118 13960 44164
rect 70824 44174 70870 44220
rect 70928 44174 70974 44220
rect 70824 44070 70870 44116
rect 70928 44070 70974 44116
rect 14046 43986 14092 44032
rect 70824 43966 70870 44012
rect 70928 43966 70974 44012
rect 14178 43854 14224 43900
rect 70824 43862 70870 43908
rect 70928 43862 70974 43908
rect 14310 43722 14356 43768
rect 70824 43758 70870 43804
rect 70928 43758 70974 43804
rect 70824 43654 70870 43700
rect 70928 43654 70974 43700
rect 14442 43590 14488 43636
rect 70824 43550 70870 43596
rect 70928 43550 70974 43596
rect 14574 43458 14620 43504
rect 70824 43446 70870 43492
rect 70928 43446 70974 43492
rect 14706 43326 14752 43372
rect 70824 43342 70870 43388
rect 70928 43342 70974 43388
rect 14838 43194 14884 43240
rect 70824 43238 70870 43284
rect 70928 43238 70974 43284
rect 14970 43062 15016 43108
rect 70824 43134 70870 43180
rect 70928 43134 70974 43180
rect 70824 43030 70870 43076
rect 70928 43030 70974 43076
rect 15102 42930 15148 42976
rect 70824 42926 70870 42972
rect 70928 42926 70974 42972
rect 15234 42798 15280 42844
rect 70824 42822 70870 42868
rect 70928 42822 70974 42868
rect 15366 42666 15412 42712
rect 70824 42718 70870 42764
rect 70928 42718 70974 42764
rect 70824 42614 70870 42660
rect 70928 42614 70974 42660
rect 15498 42534 15544 42580
rect 70824 42510 70870 42556
rect 70928 42510 70974 42556
rect 15630 42402 15676 42448
rect 70824 42406 70870 42452
rect 70928 42406 70974 42452
rect 15762 42270 15808 42316
rect 70824 42302 70870 42348
rect 70928 42302 70974 42348
rect 70824 42198 70870 42244
rect 70928 42198 70974 42244
rect 15894 42138 15940 42184
rect 70824 42094 70870 42140
rect 70928 42094 70974 42140
rect 16026 42006 16072 42052
rect 70824 41990 70870 42036
rect 70928 41990 70974 42036
rect 16158 41874 16204 41920
rect 70824 41886 70870 41932
rect 70928 41886 70974 41932
rect 16290 41742 16336 41788
rect 70824 41782 70870 41828
rect 70928 41782 70974 41828
rect 16422 41610 16468 41656
rect 70824 41678 70870 41724
rect 70928 41678 70974 41724
rect 70824 41574 70870 41620
rect 70928 41574 70974 41620
rect 16554 41478 16600 41524
rect 70824 41470 70870 41516
rect 70928 41470 70974 41516
rect 16686 41346 16732 41392
rect 70824 41366 70870 41412
rect 70928 41366 70974 41412
rect 16818 41214 16864 41260
rect 70824 41262 70870 41308
rect 70928 41262 70974 41308
rect 70824 41158 70870 41204
rect 70928 41158 70974 41204
rect 16950 41082 16996 41128
rect 70824 41054 70870 41100
rect 70928 41054 70974 41100
rect 17082 40950 17128 40996
rect 70824 40950 70870 40996
rect 70928 40950 70974 40996
rect 17214 40818 17260 40864
rect 70824 40846 70870 40892
rect 70928 40846 70974 40892
rect 17346 40686 17392 40732
rect 70824 40742 70870 40788
rect 70928 40742 70974 40788
rect 70824 40638 70870 40684
rect 70928 40638 70974 40684
rect 17478 40554 17524 40600
rect 70824 40534 70870 40580
rect 70928 40534 70974 40580
rect 17610 40422 17656 40468
rect 70824 40430 70870 40476
rect 70928 40430 70974 40476
rect 17742 40290 17788 40336
rect 70824 40326 70870 40372
rect 70928 40326 70974 40372
rect 17874 40158 17920 40204
rect 70824 40222 70870 40268
rect 70928 40222 70974 40268
rect 70824 40118 70870 40164
rect 70928 40118 70974 40164
rect 18006 40026 18052 40072
rect 70824 40014 70870 40060
rect 70928 40014 70974 40060
rect 18138 39894 18184 39940
rect 70824 39910 70870 39956
rect 70928 39910 70974 39956
rect 18270 39762 18316 39808
rect 70824 39806 70870 39852
rect 70928 39806 70974 39852
rect 70824 39702 70870 39748
rect 70928 39702 70974 39748
rect 18402 39630 18448 39676
rect 70824 39598 70870 39644
rect 70928 39598 70974 39644
rect 18534 39498 18580 39544
rect 70824 39494 70870 39540
rect 70928 39494 70974 39540
rect 18666 39366 18712 39412
rect 70824 39390 70870 39436
rect 70928 39390 70974 39436
rect 18798 39234 18844 39280
rect 70824 39286 70870 39332
rect 70928 39286 70974 39332
rect 70824 39182 70870 39228
rect 70928 39182 70974 39228
rect 18930 39102 18976 39148
rect 70824 39078 70870 39124
rect 70928 39078 70974 39124
rect 19062 38970 19108 39016
rect 70824 38974 70870 39020
rect 70928 38974 70974 39020
rect 19194 38838 19240 38884
rect 70824 38870 70870 38916
rect 70928 38870 70974 38916
rect 70824 38766 70870 38812
rect 70928 38766 70974 38812
rect 19326 38706 19372 38752
rect 70824 38662 70870 38708
rect 70928 38662 70974 38708
rect 19458 38574 19504 38620
rect 70824 38558 70870 38604
rect 70928 38558 70974 38604
rect 19590 38442 19636 38488
rect 70824 38454 70870 38500
rect 70928 38454 70974 38500
rect 19722 38310 19768 38356
rect 70824 38350 70870 38396
rect 70928 38350 70974 38396
rect 19854 38178 19900 38224
rect 70824 38246 70870 38292
rect 70928 38246 70974 38292
rect 70824 38142 70870 38188
rect 70928 38142 70974 38188
rect 19986 38046 20032 38092
rect 70824 38038 70870 38084
rect 70928 38038 70974 38084
rect 20118 37914 20164 37960
rect 70824 37934 70870 37980
rect 70928 37934 70974 37980
rect 20250 37782 20296 37828
rect 70824 37830 70870 37876
rect 70928 37830 70974 37876
rect 70824 37726 70870 37772
rect 70928 37726 70974 37772
rect 20382 37650 20428 37696
rect 70824 37622 70870 37668
rect 70928 37622 70974 37668
rect 20514 37518 20560 37564
rect 70824 37518 70870 37564
rect 70928 37518 70974 37564
rect 20646 37386 20692 37432
rect 70824 37414 70870 37460
rect 70928 37414 70974 37460
rect 70824 37310 70870 37356
rect 70928 37310 70974 37356
rect 20778 37254 20824 37300
rect 20910 37122 20956 37168
rect 70824 37206 70870 37252
rect 70928 37206 70974 37252
rect 70824 37102 70870 37148
rect 70928 37102 70974 37148
rect 21042 36990 21088 37036
rect 70824 36998 70870 37044
rect 70928 36998 70974 37044
rect 21174 36858 21220 36904
rect 70824 36894 70870 36940
rect 70928 36894 70974 36940
rect 21306 36726 21352 36772
rect 70824 36790 70870 36836
rect 70928 36790 70974 36836
rect 70824 36686 70870 36732
rect 70928 36686 70974 36732
rect 21438 36594 21484 36640
rect 70824 36582 70870 36628
rect 70928 36582 70974 36628
rect 21570 36462 21616 36508
rect 70824 36478 70870 36524
rect 70928 36478 70974 36524
rect 21702 36330 21748 36376
rect 70824 36374 70870 36420
rect 70928 36374 70974 36420
rect 70824 36270 70870 36316
rect 70928 36270 70974 36316
rect 21834 36198 21880 36244
rect 70824 36166 70870 36212
rect 70928 36166 70974 36212
rect 21966 36066 22012 36112
rect 70824 36062 70870 36108
rect 70928 36062 70974 36108
rect 22098 35934 22144 35980
rect 70824 35958 70870 36004
rect 70928 35958 70974 36004
rect 70824 35854 70870 35900
rect 70928 35854 70974 35900
rect 22230 35802 22276 35848
rect 70824 35750 70870 35796
rect 70928 35750 70974 35796
rect 22362 35670 22408 35716
rect 70824 35646 70870 35692
rect 70928 35646 70974 35692
rect 22494 35538 22540 35584
rect 70824 35542 70870 35588
rect 70928 35542 70974 35588
rect 22626 35406 22672 35452
rect 70824 35438 70870 35484
rect 70928 35438 70974 35484
rect 70824 35334 70870 35380
rect 70928 35334 70974 35380
rect 22758 35274 22804 35320
rect 70824 35230 70870 35276
rect 70928 35230 70974 35276
rect 22890 35142 22936 35188
rect 70824 35126 70870 35172
rect 70928 35126 70974 35172
rect 23022 35010 23068 35056
rect 70824 35022 70870 35068
rect 70928 35022 70974 35068
rect 23154 34878 23200 34924
rect 70824 34918 70870 34964
rect 70928 34918 70974 34964
rect 70824 34814 70870 34860
rect 70928 34814 70974 34860
rect 23286 34746 23332 34792
rect 70824 34710 70870 34756
rect 70928 34710 70974 34756
rect 23418 34614 23464 34660
rect 70824 34606 70870 34652
rect 70928 34606 70974 34652
rect 23550 34482 23596 34528
rect 70824 34502 70870 34548
rect 70928 34502 70974 34548
rect 23682 34350 23728 34396
rect 70824 34398 70870 34444
rect 70928 34398 70974 34444
rect 70824 34294 70870 34340
rect 70928 34294 70974 34340
rect 23814 34218 23860 34264
rect 70824 34190 70870 34236
rect 70928 34190 70974 34236
rect 23946 34086 23992 34132
rect 70824 34086 70870 34132
rect 70928 34086 70974 34132
rect 24078 33954 24124 34000
rect 70824 33982 70870 34028
rect 70928 33982 70974 34028
rect 70824 33878 70870 33924
rect 70928 33878 70974 33924
rect 24210 33822 24256 33868
rect 70824 33774 70870 33820
rect 70928 33774 70974 33820
rect 24342 33690 24388 33736
rect 70824 33670 70870 33716
rect 70928 33670 70974 33716
rect 24474 33558 24520 33604
rect 70824 33566 70870 33612
rect 70928 33566 70974 33612
rect 24606 33426 24652 33472
rect 70824 33462 70870 33508
rect 70928 33462 70974 33508
rect 70824 33358 70870 33404
rect 70928 33358 70974 33404
rect 24738 33294 24784 33340
rect 70824 33254 70870 33300
rect 70928 33254 70974 33300
rect 24870 33162 24916 33208
rect 70824 33150 70870 33196
rect 70928 33150 70974 33196
rect 25002 33030 25048 33076
rect 70824 33046 70870 33092
rect 70928 33046 70974 33092
rect 25134 32898 25180 32944
rect 70824 32942 70870 32988
rect 70928 32942 70974 32988
rect 70824 32838 70870 32884
rect 70928 32838 70974 32884
rect 25266 32766 25312 32812
rect 70824 32734 70870 32780
rect 70928 32734 70974 32780
rect 25398 32634 25444 32680
rect 70824 32630 70870 32676
rect 70928 32630 70974 32676
rect 25530 32502 25576 32548
rect 70824 32526 70870 32572
rect 70928 32526 70974 32572
rect 25662 32370 25708 32416
rect 70824 32422 70870 32468
rect 70928 32422 70974 32468
rect 70824 32318 70870 32364
rect 70928 32318 70974 32364
rect 25794 32238 25840 32284
rect 70824 32214 70870 32260
rect 70928 32214 70974 32260
rect 25926 32106 25972 32152
rect 70824 32110 70870 32156
rect 70928 32110 70974 32156
rect 26058 31974 26104 32020
rect 70824 32006 70870 32052
rect 70928 32006 70974 32052
rect 26190 31842 26236 31888
rect 70824 31902 70870 31948
rect 70928 31902 70974 31948
rect 70824 31798 70870 31844
rect 70928 31798 70974 31844
rect 26322 31710 26368 31756
rect 70824 31694 70870 31740
rect 70928 31694 70974 31740
rect 26454 31578 26500 31624
rect 70824 31590 70870 31636
rect 70928 31590 70974 31636
rect 26586 31446 26632 31492
rect 70824 31486 70870 31532
rect 70928 31486 70974 31532
rect 26718 31314 26764 31360
rect 70824 31382 70870 31428
rect 70928 31382 70974 31428
rect 70824 31278 70870 31324
rect 70928 31278 70974 31324
rect 26850 31182 26896 31228
rect 70824 31174 70870 31220
rect 70928 31174 70974 31220
rect 26982 31050 27028 31096
rect 70824 31070 70870 31116
rect 70928 31070 70974 31116
rect 27114 30918 27160 30964
rect 70824 30966 70870 31012
rect 70928 30966 70974 31012
rect 70824 30862 70870 30908
rect 70928 30862 70974 30908
rect 27246 30786 27292 30832
rect 70824 30758 70870 30804
rect 70928 30758 70974 30804
rect 27378 30654 27424 30700
rect 70824 30654 70870 30700
rect 70928 30654 70974 30700
rect 27510 30522 27556 30568
rect 70824 30550 70870 30596
rect 70928 30550 70974 30596
rect 27642 30390 27688 30436
rect 70824 30446 70870 30492
rect 70928 30446 70974 30492
rect 70824 30342 70870 30388
rect 70928 30342 70974 30388
rect 27774 30258 27820 30304
rect 70824 30238 70870 30284
rect 70928 30238 70974 30284
rect 27906 30126 27952 30172
rect 70824 30134 70870 30180
rect 70928 30134 70974 30180
rect 28038 29994 28084 30040
rect 70824 30030 70870 30076
rect 70928 30030 70974 30076
rect 28170 29862 28216 29908
rect 70824 29926 70870 29972
rect 70928 29926 70974 29972
rect 70824 29822 70870 29868
rect 70928 29822 70974 29868
rect 28302 29730 28348 29776
rect 70824 29718 70870 29764
rect 70928 29718 70974 29764
rect 28434 29598 28480 29644
rect 70824 29614 70870 29660
rect 70928 29614 70974 29660
rect 28566 29466 28612 29512
rect 70824 29510 70870 29556
rect 70928 29510 70974 29556
rect 28698 29334 28744 29380
rect 70824 29406 70870 29452
rect 70928 29406 70974 29452
rect 70824 29302 70870 29348
rect 70928 29302 70974 29348
rect 28830 29202 28876 29248
rect 70824 29198 70870 29244
rect 70928 29198 70974 29244
rect 28962 29070 29008 29116
rect 70824 29094 70870 29140
rect 70928 29094 70974 29140
rect 29094 28938 29140 28984
rect 70824 28990 70870 29036
rect 70928 28990 70974 29036
rect 29226 28806 29272 28852
rect 70824 28886 70870 28932
rect 70928 28886 70974 28932
rect 70824 28782 70870 28828
rect 70928 28782 70974 28828
rect 29358 28674 29404 28720
rect 70824 28678 70870 28724
rect 70928 28678 70974 28724
rect 29490 28542 29536 28588
rect 70824 28574 70870 28620
rect 70928 28574 70974 28620
rect 29622 28410 29668 28456
rect 70824 28470 70870 28516
rect 70928 28470 70974 28516
rect 70824 28366 70870 28412
rect 70928 28366 70974 28412
rect 29754 28278 29800 28324
rect 70824 28262 70870 28308
rect 70928 28262 70974 28308
rect 29886 28146 29932 28192
rect 70824 28158 70870 28204
rect 70928 28158 70974 28204
rect 30018 28014 30064 28060
rect 70824 28054 70870 28100
rect 70928 28054 70974 28100
rect 30150 27882 30196 27928
rect 70824 27950 70870 27996
rect 70928 27950 70974 27996
rect 70824 27846 70870 27892
rect 70928 27846 70974 27892
rect 30282 27750 30328 27796
rect 70824 27742 70870 27788
rect 70928 27742 70974 27788
rect 30414 27618 30460 27664
rect 70824 27638 70870 27684
rect 70928 27638 70974 27684
rect 30546 27486 30592 27532
rect 70824 27534 70870 27580
rect 70928 27534 70974 27580
rect 70824 27430 70870 27476
rect 70928 27430 70974 27476
rect 30678 27354 30724 27400
rect 70824 27326 70870 27372
rect 70928 27326 70974 27372
rect 30810 27222 30856 27268
rect 70824 27222 70870 27268
rect 70928 27222 70974 27268
rect 30942 27090 30988 27136
rect 70824 27118 70870 27164
rect 70928 27118 70974 27164
rect 70824 27014 70870 27060
rect 70928 27014 70974 27060
rect 31074 26958 31120 27004
rect 31206 26826 31252 26872
rect 70824 26910 70870 26956
rect 70928 26910 70974 26956
rect 70824 26806 70870 26852
rect 70928 26806 70974 26852
rect 31338 26694 31384 26740
rect 70824 26702 70870 26748
rect 70928 26702 70974 26748
rect 31470 26562 31516 26608
rect 70824 26598 70870 26644
rect 70928 26598 70974 26644
rect 31602 26430 31648 26476
rect 70824 26494 70870 26540
rect 70928 26494 70974 26540
rect 70824 26390 70870 26436
rect 70928 26390 70974 26436
rect 31734 26298 31780 26344
rect 70824 26286 70870 26332
rect 70928 26286 70974 26332
rect 31866 26166 31912 26212
rect 70824 26182 70870 26228
rect 70928 26182 70974 26228
rect 31998 26034 32044 26080
rect 70824 26078 70870 26124
rect 70928 26078 70974 26124
rect 70824 25974 70870 26020
rect 70928 25974 70974 26020
rect 32130 25902 32176 25948
rect 70824 25870 70870 25916
rect 70928 25870 70974 25916
rect 32262 25770 32308 25816
rect 70824 25766 70870 25812
rect 70928 25766 70974 25812
rect 32394 25638 32440 25684
rect 70824 25662 70870 25708
rect 70928 25662 70974 25708
rect 32526 25506 32572 25552
rect 70824 25558 70870 25604
rect 70928 25558 70974 25604
rect 32658 25374 32704 25420
rect 70824 25454 70870 25500
rect 70928 25454 70974 25500
rect 70824 25350 70870 25396
rect 70928 25350 70974 25396
rect 32790 25242 32836 25288
rect 70824 25246 70870 25292
rect 70928 25246 70974 25292
rect 32922 25110 32968 25156
rect 70824 25142 70870 25188
rect 70928 25142 70974 25188
rect 33054 24978 33100 25024
rect 70824 25038 70870 25084
rect 70928 25038 70974 25084
rect 70824 24934 70870 24980
rect 70928 24934 70974 24980
rect 33186 24846 33232 24892
rect 70824 24830 70870 24876
rect 70928 24830 70974 24876
rect 33318 24714 33364 24760
rect 70824 24726 70870 24772
rect 70928 24726 70974 24772
rect 33450 24582 33496 24628
rect 70824 24622 70870 24668
rect 70928 24622 70974 24668
rect 70824 24518 70870 24564
rect 70928 24518 70974 24564
rect 33582 24450 33628 24496
rect 70824 24414 70870 24460
rect 70928 24414 70974 24460
rect 33714 24318 33760 24364
rect 70824 24310 70870 24356
rect 70928 24310 70974 24356
rect 33846 24186 33892 24232
rect 70824 24206 70870 24252
rect 70928 24206 70974 24252
rect 33978 24054 34024 24100
rect 70824 24102 70870 24148
rect 70928 24102 70974 24148
rect 70824 23998 70870 24044
rect 70928 23998 70974 24044
rect 34110 23922 34156 23968
rect 70824 23894 70870 23940
rect 70928 23894 70974 23940
rect 34242 23790 34288 23836
rect 70824 23790 70870 23836
rect 70928 23790 70974 23836
rect 34374 23658 34420 23704
rect 70824 23686 70870 23732
rect 70928 23686 70974 23732
rect 34506 23526 34552 23572
rect 70824 23582 70870 23628
rect 70928 23582 70974 23628
rect 70824 23478 70870 23524
rect 70928 23478 70974 23524
rect 34638 23394 34684 23440
rect 70824 23374 70870 23420
rect 70928 23374 70974 23420
rect 34770 23262 34816 23308
rect 70824 23270 70870 23316
rect 70928 23270 70974 23316
rect 34902 23130 34948 23176
rect 70824 23166 70870 23212
rect 70928 23166 70974 23212
rect 35034 22998 35080 23044
rect 70824 23062 70870 23108
rect 70928 23062 70974 23108
rect 70824 22958 70870 23004
rect 70928 22958 70974 23004
rect 35166 22866 35212 22912
rect 70824 22854 70870 22900
rect 70928 22854 70974 22900
rect 35298 22734 35344 22780
rect 70824 22750 70870 22796
rect 70928 22750 70974 22796
rect 35430 22602 35476 22648
rect 70824 22646 70870 22692
rect 70928 22646 70974 22692
rect 70824 22542 70870 22588
rect 70928 22542 70974 22588
rect 35562 22470 35608 22516
rect 70824 22438 70870 22484
rect 70928 22438 70974 22484
rect 35694 22338 35740 22384
rect 70824 22334 70870 22380
rect 70928 22334 70974 22380
rect 35826 22206 35872 22252
rect 70824 22230 70870 22276
rect 70928 22230 70974 22276
rect 70824 22126 70870 22172
rect 70928 22126 70974 22172
rect 35958 22074 36004 22120
rect 70824 22022 70870 22068
rect 70928 22022 70974 22068
rect 36090 21942 36136 21988
rect 70824 21918 70870 21964
rect 70928 21918 70974 21964
rect 36222 21810 36268 21856
rect 70824 21814 70870 21860
rect 70928 21814 70974 21860
rect 36354 21678 36400 21724
rect 70824 21710 70870 21756
rect 70928 21710 70974 21756
rect 36486 21546 36532 21592
rect 70824 21606 70870 21652
rect 70928 21606 70974 21652
rect 70824 21502 70870 21548
rect 70928 21502 70974 21548
rect 36618 21414 36664 21460
rect 70824 21398 70870 21444
rect 70928 21398 70974 21444
rect 36750 21282 36796 21328
rect 70824 21294 70870 21340
rect 70928 21294 70974 21340
rect 36882 21150 36928 21196
rect 70824 21190 70870 21236
rect 70928 21190 70974 21236
rect 70824 21086 70870 21132
rect 70928 21086 70974 21132
rect 37014 21018 37060 21064
rect 70824 20982 70870 21028
rect 70928 20982 70974 21028
rect 37146 20886 37192 20932
rect 70824 20878 70870 20924
rect 70928 20878 70974 20924
rect 37278 20754 37324 20800
rect 70824 20774 70870 20820
rect 70928 20774 70974 20820
rect 37410 20622 37456 20668
rect 70824 20670 70870 20716
rect 70928 20670 70974 20716
rect 37542 20490 37588 20536
rect 70824 20566 70870 20612
rect 70928 20566 70974 20612
rect 70824 20462 70870 20508
rect 70928 20462 70974 20508
rect 37674 20358 37720 20404
rect 70824 20358 70870 20404
rect 70928 20358 70974 20404
rect 37806 20226 37852 20272
rect 70824 20254 70870 20300
rect 70928 20254 70974 20300
rect 37938 20094 37984 20140
rect 70824 20150 70870 20196
rect 70928 20150 70974 20196
rect 70824 20046 70870 20092
rect 70928 20046 70974 20092
rect 38070 19962 38116 20008
rect 70824 19942 70870 19988
rect 70928 19942 70974 19988
rect 38202 19830 38248 19876
rect 70824 19838 70870 19884
rect 70928 19838 70974 19884
rect 38334 19698 38380 19744
rect 70824 19734 70870 19780
rect 70928 19734 70974 19780
rect 38466 19566 38512 19612
rect 70824 19630 70870 19676
rect 70928 19630 70974 19676
rect 70824 19526 70870 19572
rect 70928 19526 70974 19572
rect 38598 19434 38644 19480
rect 70824 19422 70870 19468
rect 70928 19422 70974 19468
rect 38730 19302 38776 19348
rect 70824 19318 70870 19364
rect 70928 19318 70974 19364
rect 38862 19170 38908 19216
rect 70824 19214 70870 19260
rect 70928 19214 70974 19260
rect 70824 19110 70870 19156
rect 70928 19110 70974 19156
rect 38994 19038 39040 19084
rect 70824 19006 70870 19052
rect 70928 19006 70974 19052
rect 39126 18906 39172 18952
rect 70824 18902 70870 18948
rect 70928 18902 70974 18948
rect 39258 18774 39304 18820
rect 70824 18798 70870 18844
rect 70928 18798 70974 18844
rect 39390 18642 39436 18688
rect 70824 18694 70870 18740
rect 70928 18694 70974 18740
rect 39522 18510 39568 18556
rect 70824 18590 70870 18636
rect 70928 18590 70974 18636
rect 70824 18486 70870 18532
rect 70928 18486 70974 18532
rect 39654 18378 39700 18424
rect 70824 18382 70870 18428
rect 70928 18382 70974 18428
rect 39786 18246 39832 18292
rect 70824 18278 70870 18324
rect 70928 18278 70974 18324
rect 39918 18114 39964 18160
rect 70824 18174 70870 18220
rect 70928 18174 70974 18220
rect 70824 18070 70870 18116
rect 70928 18070 70974 18116
rect 40050 17982 40096 18028
rect 70824 17966 70870 18012
rect 70928 17966 70974 18012
rect 40182 17850 40228 17896
rect 70824 17862 70870 17908
rect 70928 17862 70974 17908
rect 40314 17718 40360 17764
rect 70824 17758 70870 17804
rect 70928 17758 70974 17804
rect 40446 17586 40492 17632
rect 70824 17654 70870 17700
rect 70928 17654 70974 17700
rect 70824 17550 70870 17596
rect 70928 17550 70974 17596
rect 40578 17454 40624 17500
rect 70824 17446 70870 17492
rect 70928 17446 70974 17492
rect 40710 17322 40756 17368
rect 70824 17342 70870 17388
rect 70928 17342 70974 17388
rect 40842 17190 40888 17236
rect 70824 17238 70870 17284
rect 70928 17238 70974 17284
rect 70824 17134 70870 17180
rect 70928 17134 70974 17180
rect 40974 17058 41020 17104
rect 70824 17030 70870 17076
rect 70928 17030 70974 17076
rect 41106 16926 41152 16972
rect 70824 16926 70870 16972
rect 70928 16926 70974 16972
rect 41238 16794 41284 16840
rect 70824 16822 70870 16868
rect 70928 16822 70974 16868
rect 41370 16662 41416 16708
rect 70824 16718 70870 16764
rect 70928 16718 70974 16764
rect 70824 16614 70870 16660
rect 70928 16614 70974 16660
rect 41502 16530 41548 16576
rect 70824 16510 70870 16556
rect 70928 16510 70974 16556
rect 41634 16398 41680 16444
rect 70824 16406 70870 16452
rect 70928 16406 70974 16452
rect 41766 16266 41812 16312
rect 70824 16302 70870 16348
rect 70928 16302 70974 16348
rect 70824 16198 70870 16244
rect 70928 16198 70974 16244
rect 41898 16134 41944 16180
rect 70824 16094 70870 16140
rect 70928 16094 70974 16140
rect 42030 16002 42076 16048
rect 70824 15990 70870 16036
rect 70928 15990 70974 16036
rect 42162 15870 42208 15916
rect 70824 15886 70870 15932
rect 70928 15886 70974 15932
rect 42294 15738 42340 15784
rect 70824 15782 70870 15828
rect 70928 15782 70974 15828
rect 70824 15678 70870 15724
rect 70928 15678 70974 15724
rect 42426 15606 42472 15652
rect 70824 15574 70870 15620
rect 70928 15574 70974 15620
rect 42558 15474 42604 15520
rect 70824 15470 70870 15516
rect 70928 15470 70974 15516
rect 42690 15342 42736 15388
rect 70824 15366 70870 15412
rect 70928 15366 70974 15412
rect 70824 15262 70870 15308
rect 70928 15262 70974 15308
rect 42822 15210 42868 15256
rect 70824 15158 70870 15204
rect 70928 15158 70974 15204
rect 42954 15078 43000 15124
rect 70824 15054 70870 15100
rect 70928 15054 70974 15100
rect 43086 14946 43132 14992
rect 70824 14950 70870 14996
rect 70928 14950 70974 14996
rect 43218 14814 43264 14860
rect 70824 14846 70870 14892
rect 70928 14846 70974 14892
rect 70824 14742 70870 14788
rect 70928 14742 70974 14788
rect 43350 14682 43396 14728
rect 70824 14638 70870 14684
rect 70928 14638 70974 14684
rect 43482 14550 43528 14596
rect 70824 14534 70870 14580
rect 70928 14534 70974 14580
rect 43614 14418 43660 14464
rect 70824 14430 70870 14476
rect 70928 14430 70974 14476
rect 43746 14286 43792 14332
rect 70824 14326 70870 14372
rect 70928 14326 70974 14372
rect 70824 14222 70870 14268
rect 70928 14222 70974 14268
rect 43878 14154 43924 14200
rect 70824 14118 70870 14164
rect 70928 14118 70974 14164
rect 44010 14022 44056 14068
rect 70824 14014 70870 14060
rect 70928 14014 70974 14060
rect 44142 13890 44188 13936
rect 70824 13910 70870 13956
rect 70928 13910 70974 13956
rect 44274 13758 44320 13804
rect 70824 13806 70870 13852
rect 70928 13806 70974 13852
rect 70824 13702 70870 13748
rect 70928 13702 70974 13748
rect 44406 13626 44452 13672
rect 70824 13598 70870 13644
rect 70928 13598 70974 13644
rect 44538 13494 44584 13540
rect 70824 13494 70870 13540
rect 70928 13494 70974 13540
rect 44670 13362 44716 13408
rect 70824 13390 70870 13436
rect 70928 13390 70974 13436
rect 44850 13210 44896 13256
rect 45088 13223 45134 13269
rect 45192 13223 45238 13269
rect 45296 13223 45342 13269
rect 45400 13223 45446 13269
rect 45504 13223 45550 13269
rect 45608 13223 45654 13269
rect 45712 13223 45758 13269
rect 45816 13223 45862 13269
rect 45920 13223 45966 13269
rect 46024 13223 46070 13269
rect 46128 13223 46174 13269
rect 46232 13223 46278 13269
rect 46336 13223 46382 13269
rect 46440 13223 46486 13269
rect 46544 13223 46590 13269
rect 46648 13223 46694 13269
rect 46752 13223 46798 13269
rect 46856 13223 46902 13269
rect 46960 13223 47006 13269
rect 47064 13223 47110 13269
rect 47168 13223 47214 13269
rect 47272 13223 47318 13269
rect 47376 13223 47422 13269
rect 47480 13223 47526 13269
rect 47584 13223 47630 13269
rect 47688 13223 47734 13269
rect 47792 13223 47838 13269
rect 47896 13223 47942 13269
rect 48000 13223 48046 13269
rect 48104 13223 48150 13269
rect 48208 13223 48254 13269
rect 48312 13223 48358 13269
rect 48416 13223 48462 13269
rect 48520 13223 48566 13269
rect 48624 13223 48670 13269
rect 48728 13223 48774 13269
rect 48832 13223 48878 13269
rect 48936 13223 48982 13269
rect 49040 13223 49086 13269
rect 49144 13223 49190 13269
rect 49248 13223 49294 13269
rect 49352 13223 49398 13269
rect 49456 13223 49502 13269
rect 49560 13223 49606 13269
rect 49664 13223 49710 13269
rect 49768 13223 49814 13269
rect 49872 13223 49918 13269
rect 49976 13223 50022 13269
rect 50080 13223 50126 13269
rect 50184 13223 50230 13269
rect 50288 13223 50334 13269
rect 50392 13223 50438 13269
rect 50496 13223 50542 13269
rect 50600 13223 50646 13269
rect 50704 13223 50750 13269
rect 50808 13223 50854 13269
rect 50912 13223 50958 13269
rect 51016 13223 51062 13269
rect 51120 13223 51166 13269
rect 51224 13223 51270 13269
rect 51328 13223 51374 13269
rect 51432 13223 51478 13269
rect 51536 13223 51582 13269
rect 51640 13223 51686 13269
rect 51744 13223 51790 13269
rect 51848 13223 51894 13269
rect 51952 13223 51998 13269
rect 52056 13223 52102 13269
rect 52160 13223 52206 13269
rect 52264 13223 52310 13269
rect 52368 13223 52414 13269
rect 52472 13223 52518 13269
rect 52576 13223 52622 13269
rect 52680 13223 52726 13269
rect 52784 13223 52830 13269
rect 52888 13223 52934 13269
rect 52992 13223 53038 13269
rect 53096 13223 53142 13269
rect 53200 13223 53246 13269
rect 53304 13223 53350 13269
rect 53408 13223 53454 13269
rect 53512 13223 53558 13269
rect 53616 13223 53662 13269
rect 53720 13223 53766 13269
rect 53824 13223 53870 13269
rect 53928 13223 53974 13269
rect 54032 13223 54078 13269
rect 54136 13223 54182 13269
rect 54240 13223 54286 13269
rect 54344 13223 54390 13269
rect 54448 13223 54494 13269
rect 54552 13223 54598 13269
rect 54656 13223 54702 13269
rect 54760 13223 54806 13269
rect 54864 13223 54910 13269
rect 54968 13223 55014 13269
rect 55072 13223 55118 13269
rect 55176 13223 55222 13269
rect 55280 13223 55326 13269
rect 55384 13223 55430 13269
rect 55488 13223 55534 13269
rect 55592 13223 55638 13269
rect 55696 13223 55742 13269
rect 55800 13223 55846 13269
rect 55904 13223 55950 13269
rect 56008 13223 56054 13269
rect 56112 13223 56158 13269
rect 56216 13223 56262 13269
rect 56320 13223 56366 13269
rect 56424 13223 56470 13269
rect 56528 13223 56574 13269
rect 56632 13223 56678 13269
rect 56736 13223 56782 13269
rect 56840 13223 56886 13269
rect 56944 13223 56990 13269
rect 57048 13223 57094 13269
rect 57152 13223 57198 13269
rect 57256 13223 57302 13269
rect 57360 13223 57406 13269
rect 57464 13223 57510 13269
rect 57568 13223 57614 13269
rect 57672 13223 57718 13269
rect 57776 13223 57822 13269
rect 57880 13223 57926 13269
rect 57984 13223 58030 13269
rect 58088 13223 58134 13269
rect 58192 13223 58238 13269
rect 58296 13223 58342 13269
rect 58400 13223 58446 13269
rect 58504 13223 58550 13269
rect 58608 13223 58654 13269
rect 58712 13223 58758 13269
rect 58816 13223 58862 13269
rect 58920 13223 58966 13269
rect 59024 13223 59070 13269
rect 59128 13223 59174 13269
rect 59232 13223 59278 13269
rect 59336 13223 59382 13269
rect 59440 13223 59486 13269
rect 59544 13223 59590 13269
rect 59648 13223 59694 13269
rect 59752 13223 59798 13269
rect 59856 13223 59902 13269
rect 59960 13223 60006 13269
rect 60064 13223 60110 13269
rect 60168 13223 60214 13269
rect 60272 13223 60318 13269
rect 60376 13223 60422 13269
rect 60480 13223 60526 13269
rect 60584 13223 60630 13269
rect 60688 13223 60734 13269
rect 60792 13223 60838 13269
rect 60896 13223 60942 13269
rect 61000 13223 61046 13269
rect 61104 13223 61150 13269
rect 61208 13223 61254 13269
rect 61312 13223 61358 13269
rect 61416 13223 61462 13269
rect 61520 13223 61566 13269
rect 61624 13223 61670 13269
rect 61728 13223 61774 13269
rect 61832 13223 61878 13269
rect 61936 13223 61982 13269
rect 62040 13223 62086 13269
rect 62144 13223 62190 13269
rect 62248 13223 62294 13269
rect 62352 13223 62398 13269
rect 62456 13223 62502 13269
rect 62560 13223 62606 13269
rect 62664 13223 62710 13269
rect 62768 13223 62814 13269
rect 62872 13223 62918 13269
rect 62976 13223 63022 13269
rect 63080 13223 63126 13269
rect 63184 13223 63230 13269
rect 63288 13223 63334 13269
rect 63392 13223 63438 13269
rect 63496 13223 63542 13269
rect 63600 13223 63646 13269
rect 63704 13223 63750 13269
rect 63808 13223 63854 13269
rect 63912 13223 63958 13269
rect 64016 13223 64062 13269
rect 64120 13223 64166 13269
rect 64224 13223 64270 13269
rect 64328 13223 64374 13269
rect 64432 13223 64478 13269
rect 64536 13223 64582 13269
rect 64640 13223 64686 13269
rect 64744 13223 64790 13269
rect 64848 13223 64894 13269
rect 64952 13223 64998 13269
rect 65056 13223 65102 13269
rect 65160 13223 65206 13269
rect 65264 13223 65310 13269
rect 65368 13223 65414 13269
rect 65472 13223 65518 13269
rect 65576 13223 65622 13269
rect 65680 13223 65726 13269
rect 65784 13223 65830 13269
rect 65888 13223 65934 13269
rect 65992 13223 66038 13269
rect 66096 13223 66142 13269
rect 66200 13223 66246 13269
rect 66304 13223 66350 13269
rect 66408 13223 66454 13269
rect 66512 13223 66558 13269
rect 66616 13223 66662 13269
rect 66720 13223 66766 13269
rect 66824 13223 66870 13269
rect 66928 13223 66974 13269
rect 67032 13223 67078 13269
rect 67136 13223 67182 13269
rect 67240 13223 67286 13269
rect 67344 13223 67390 13269
rect 67448 13223 67494 13269
rect 67552 13223 67598 13269
rect 67656 13223 67702 13269
rect 67760 13223 67806 13269
rect 67864 13223 67910 13269
rect 67968 13223 68014 13269
rect 68072 13223 68118 13269
rect 68176 13223 68222 13269
rect 68280 13223 68326 13269
rect 68384 13223 68430 13269
rect 68488 13223 68534 13269
rect 68592 13223 68638 13269
rect 68696 13223 68742 13269
rect 68800 13223 68846 13269
rect 68904 13223 68950 13269
rect 69008 13223 69054 13269
rect 69112 13223 69158 13269
rect 69216 13223 69262 13269
rect 69320 13223 69366 13269
rect 69424 13223 69470 13269
rect 69528 13223 69574 13269
rect 69632 13223 69678 13269
rect 69736 13223 69782 13269
rect 69840 13223 69886 13269
rect 69944 13223 69990 13269
rect 70048 13223 70094 13269
rect 70152 13223 70198 13269
rect 70256 13223 70302 13269
rect 70360 13223 70406 13269
rect 70464 13223 70510 13269
rect 70568 13223 70614 13269
rect 70672 13223 70718 13269
rect 70776 13223 70822 13269
rect 70880 13223 70926 13269
rect 45088 13119 45134 13165
rect 45192 13119 45238 13165
rect 45296 13119 45342 13165
rect 45400 13119 45446 13165
rect 45504 13119 45550 13165
rect 45608 13119 45654 13165
rect 45712 13119 45758 13165
rect 45816 13119 45862 13165
rect 45920 13119 45966 13165
rect 46024 13119 46070 13165
rect 46128 13119 46174 13165
rect 46232 13119 46278 13165
rect 46336 13119 46382 13165
rect 46440 13119 46486 13165
rect 46544 13119 46590 13165
rect 46648 13119 46694 13165
rect 46752 13119 46798 13165
rect 46856 13119 46902 13165
rect 46960 13119 47006 13165
rect 47064 13119 47110 13165
rect 47168 13119 47214 13165
rect 47272 13119 47318 13165
rect 47376 13119 47422 13165
rect 47480 13119 47526 13165
rect 47584 13119 47630 13165
rect 47688 13119 47734 13165
rect 47792 13119 47838 13165
rect 47896 13119 47942 13165
rect 48000 13119 48046 13165
rect 48104 13119 48150 13165
rect 48208 13119 48254 13165
rect 48312 13119 48358 13165
rect 48416 13119 48462 13165
rect 48520 13119 48566 13165
rect 48624 13119 48670 13165
rect 48728 13119 48774 13165
rect 48832 13119 48878 13165
rect 48936 13119 48982 13165
rect 49040 13119 49086 13165
rect 49144 13119 49190 13165
rect 49248 13119 49294 13165
rect 49352 13119 49398 13165
rect 49456 13119 49502 13165
rect 49560 13119 49606 13165
rect 49664 13119 49710 13165
rect 49768 13119 49814 13165
rect 49872 13119 49918 13165
rect 49976 13119 50022 13165
rect 50080 13119 50126 13165
rect 50184 13119 50230 13165
rect 50288 13119 50334 13165
rect 50392 13119 50438 13165
rect 50496 13119 50542 13165
rect 50600 13119 50646 13165
rect 50704 13119 50750 13165
rect 50808 13119 50854 13165
rect 50912 13119 50958 13165
rect 51016 13119 51062 13165
rect 51120 13119 51166 13165
rect 51224 13119 51270 13165
rect 51328 13119 51374 13165
rect 51432 13119 51478 13165
rect 51536 13119 51582 13165
rect 51640 13119 51686 13165
rect 51744 13119 51790 13165
rect 51848 13119 51894 13165
rect 51952 13119 51998 13165
rect 52056 13119 52102 13165
rect 52160 13119 52206 13165
rect 52264 13119 52310 13165
rect 52368 13119 52414 13165
rect 52472 13119 52518 13165
rect 52576 13119 52622 13165
rect 52680 13119 52726 13165
rect 52784 13119 52830 13165
rect 52888 13119 52934 13165
rect 52992 13119 53038 13165
rect 53096 13119 53142 13165
rect 53200 13119 53246 13165
rect 53304 13119 53350 13165
rect 53408 13119 53454 13165
rect 53512 13119 53558 13165
rect 53616 13119 53662 13165
rect 53720 13119 53766 13165
rect 53824 13119 53870 13165
rect 53928 13119 53974 13165
rect 54032 13119 54078 13165
rect 54136 13119 54182 13165
rect 54240 13119 54286 13165
rect 54344 13119 54390 13165
rect 54448 13119 54494 13165
rect 54552 13119 54598 13165
rect 54656 13119 54702 13165
rect 54760 13119 54806 13165
rect 54864 13119 54910 13165
rect 54968 13119 55014 13165
rect 55072 13119 55118 13165
rect 55176 13119 55222 13165
rect 55280 13119 55326 13165
rect 55384 13119 55430 13165
rect 55488 13119 55534 13165
rect 55592 13119 55638 13165
rect 55696 13119 55742 13165
rect 55800 13119 55846 13165
rect 55904 13119 55950 13165
rect 56008 13119 56054 13165
rect 56112 13119 56158 13165
rect 56216 13119 56262 13165
rect 56320 13119 56366 13165
rect 56424 13119 56470 13165
rect 56528 13119 56574 13165
rect 56632 13119 56678 13165
rect 56736 13119 56782 13165
rect 56840 13119 56886 13165
rect 56944 13119 56990 13165
rect 57048 13119 57094 13165
rect 57152 13119 57198 13165
rect 57256 13119 57302 13165
rect 57360 13119 57406 13165
rect 57464 13119 57510 13165
rect 57568 13119 57614 13165
rect 57672 13119 57718 13165
rect 57776 13119 57822 13165
rect 57880 13119 57926 13165
rect 57984 13119 58030 13165
rect 58088 13119 58134 13165
rect 58192 13119 58238 13165
rect 58296 13119 58342 13165
rect 58400 13119 58446 13165
rect 58504 13119 58550 13165
rect 58608 13119 58654 13165
rect 58712 13119 58758 13165
rect 58816 13119 58862 13165
rect 58920 13119 58966 13165
rect 59024 13119 59070 13165
rect 59128 13119 59174 13165
rect 59232 13119 59278 13165
rect 59336 13119 59382 13165
rect 59440 13119 59486 13165
rect 59544 13119 59590 13165
rect 59648 13119 59694 13165
rect 59752 13119 59798 13165
rect 59856 13119 59902 13165
rect 59960 13119 60006 13165
rect 60064 13119 60110 13165
rect 60168 13119 60214 13165
rect 60272 13119 60318 13165
rect 60376 13119 60422 13165
rect 60480 13119 60526 13165
rect 60584 13119 60630 13165
rect 60688 13119 60734 13165
rect 60792 13119 60838 13165
rect 60896 13119 60942 13165
rect 61000 13119 61046 13165
rect 61104 13119 61150 13165
rect 61208 13119 61254 13165
rect 61312 13119 61358 13165
rect 61416 13119 61462 13165
rect 61520 13119 61566 13165
rect 61624 13119 61670 13165
rect 61728 13119 61774 13165
rect 61832 13119 61878 13165
rect 61936 13119 61982 13165
rect 62040 13119 62086 13165
rect 62144 13119 62190 13165
rect 62248 13119 62294 13165
rect 62352 13119 62398 13165
rect 62456 13119 62502 13165
rect 62560 13119 62606 13165
rect 62664 13119 62710 13165
rect 62768 13119 62814 13165
rect 62872 13119 62918 13165
rect 62976 13119 63022 13165
rect 63080 13119 63126 13165
rect 63184 13119 63230 13165
rect 63288 13119 63334 13165
rect 63392 13119 63438 13165
rect 63496 13119 63542 13165
rect 63600 13119 63646 13165
rect 63704 13119 63750 13165
rect 63808 13119 63854 13165
rect 63912 13119 63958 13165
rect 64016 13119 64062 13165
rect 64120 13119 64166 13165
rect 64224 13119 64270 13165
rect 64328 13119 64374 13165
rect 64432 13119 64478 13165
rect 64536 13119 64582 13165
rect 64640 13119 64686 13165
rect 64744 13119 64790 13165
rect 64848 13119 64894 13165
rect 64952 13119 64998 13165
rect 65056 13119 65102 13165
rect 65160 13119 65206 13165
rect 65264 13119 65310 13165
rect 65368 13119 65414 13165
rect 65472 13119 65518 13165
rect 65576 13119 65622 13165
rect 65680 13119 65726 13165
rect 65784 13119 65830 13165
rect 65888 13119 65934 13165
rect 65992 13119 66038 13165
rect 66096 13119 66142 13165
rect 66200 13119 66246 13165
rect 66304 13119 66350 13165
rect 66408 13119 66454 13165
rect 66512 13119 66558 13165
rect 66616 13119 66662 13165
rect 66720 13119 66766 13165
rect 66824 13119 66870 13165
rect 66928 13119 66974 13165
rect 67032 13119 67078 13165
rect 67136 13119 67182 13165
rect 67240 13119 67286 13165
rect 67344 13119 67390 13165
rect 67448 13119 67494 13165
rect 67552 13119 67598 13165
rect 67656 13119 67702 13165
rect 67760 13119 67806 13165
rect 67864 13119 67910 13165
rect 67968 13119 68014 13165
rect 68072 13119 68118 13165
rect 68176 13119 68222 13165
rect 68280 13119 68326 13165
rect 68384 13119 68430 13165
rect 68488 13119 68534 13165
rect 68592 13119 68638 13165
rect 68696 13119 68742 13165
rect 68800 13119 68846 13165
rect 68904 13119 68950 13165
rect 69008 13119 69054 13165
rect 69112 13119 69158 13165
rect 69216 13119 69262 13165
rect 69320 13119 69366 13165
rect 69424 13119 69470 13165
rect 69528 13119 69574 13165
rect 69632 13119 69678 13165
rect 69736 13119 69782 13165
rect 69840 13119 69886 13165
rect 69944 13119 69990 13165
rect 70048 13119 70094 13165
rect 70152 13119 70198 13165
rect 70256 13119 70302 13165
rect 70360 13119 70406 13165
rect 70464 13119 70510 13165
rect 70568 13119 70614 13165
rect 70672 13119 70718 13165
rect 70776 13119 70822 13165
rect 70880 13119 70926 13165
<< metal1 >>
rect 13108 70975 69957 71000
rect 13108 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69957 70975
rect 13108 70871 69957 70929
rect 13108 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69957 70871
rect 13108 70814 69957 70825
rect 13108 70767 13280 70814
rect 13108 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13280 70767
rect 13108 70663 13280 70721
rect 13108 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13280 70663
rect 13108 70559 13280 70617
rect 13108 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13280 70559
rect 13108 70455 13280 70513
rect 13108 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13280 70455
rect 13108 70351 13280 70409
rect 13108 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13280 70351
rect 13108 70247 13280 70305
rect 13108 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13280 70247
rect 13108 70143 13280 70201
rect 13108 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13280 70143
rect 13108 70039 13280 70097
rect 13108 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13280 70039
rect 13108 69935 13280 69993
rect 13108 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13280 69935
rect 13108 69831 13280 69889
rect 13108 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13280 69831
rect 69785 70720 69957 70814
rect 69785 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69957 70720
rect 69785 70616 69957 70674
rect 69785 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69957 70616
rect 69785 70512 69957 70570
rect 69785 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69957 70512
rect 69785 70408 69957 70466
rect 69785 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69957 70408
rect 69785 70304 69957 70362
rect 69785 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69957 70304
rect 69785 70200 69957 70258
rect 69785 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69957 70200
rect 69785 70096 69957 70154
rect 69785 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69957 70096
rect 69785 69957 69957 70050
rect 69785 69946 71000 69957
rect 69785 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69785 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69785 69842 71000 69862
rect 69785 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69785 69785 70824 69796
rect 13108 69727 13280 69785
rect 13108 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13280 69727
rect 13108 69623 13280 69681
rect 13108 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13280 69623
rect 13108 69519 13280 69577
rect 13108 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13280 69519
rect 13108 69415 13280 69473
rect 13108 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13280 69415
rect 13108 69311 13280 69369
rect 13108 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13280 69311
rect 13108 69207 13280 69265
rect 13108 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13280 69207
rect 13108 69103 13280 69161
rect 13108 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13280 69103
rect 13108 68999 13280 69057
rect 13108 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13280 68999
rect 13108 68895 13280 68953
rect 13108 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13280 68895
rect 13108 68791 13280 68849
rect 13108 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13280 68791
rect 13108 68687 13280 68745
rect 13108 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13280 68687
rect 13108 68583 13280 68641
rect 13108 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13280 68583
rect 13108 68479 13280 68537
rect 13108 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13280 68479
rect 13108 68375 13280 68433
rect 13108 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13280 68375
rect 13108 68271 13280 68329
rect 13108 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13280 68271
rect 13108 68167 13280 68225
rect 13108 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13280 68167
rect 13108 68063 13280 68121
rect 13108 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13280 68063
rect 13108 67959 13280 68017
rect 13108 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13280 67959
rect 13108 67855 13280 67913
rect 13108 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13280 67855
rect 13108 67751 13280 67809
rect 13108 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13280 67751
rect 13108 67647 13280 67705
rect 13108 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13280 67647
rect 13108 67543 13280 67601
rect 13108 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13280 67543
rect 13108 67439 13280 67497
rect 13108 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13280 67439
rect 13108 67335 13280 67393
rect 13108 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13280 67335
rect 13108 67231 13280 67289
rect 13108 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13280 67231
rect 13108 67127 13280 67185
rect 13108 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13280 67127
rect 13108 67023 13280 67081
rect 13108 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13280 67023
rect 13108 66919 13280 66977
rect 13108 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13280 66919
rect 13108 66815 13280 66873
rect 13108 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13280 66815
rect 13108 66711 13280 66769
rect 13108 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13280 66711
rect 13108 66607 13280 66665
rect 13108 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13280 66607
rect 13108 66503 13280 66561
rect 13108 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13280 66503
rect 13108 66399 13280 66457
rect 13108 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13280 66399
rect 13108 66295 13280 66353
rect 13108 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13280 66295
rect 13108 66191 13280 66249
rect 13108 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13280 66191
rect 13108 66087 13280 66145
rect 13108 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13280 66087
rect 13108 65983 13280 66041
rect 13108 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13280 65983
rect 13108 65879 13280 65937
rect 13108 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13280 65879
rect 13108 65775 13280 65833
rect 13108 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13280 65775
rect 13108 65671 13280 65729
rect 13108 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13280 65671
rect 13108 65567 13280 65625
rect 13108 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13280 65567
rect 13108 65463 13280 65521
rect 13108 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13280 65463
rect 13108 65359 13280 65417
rect 13108 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13280 65359
rect 13108 65255 13280 65313
rect 13108 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13280 65255
rect 13108 65151 13280 65209
rect 13108 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13280 65151
rect 13108 65047 13280 65105
rect 13108 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13280 65047
rect 13108 64943 13280 65001
rect 13108 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13280 64943
rect 13108 64839 13280 64897
rect 13108 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13280 64839
rect 13108 64735 13280 64793
rect 13108 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13280 64735
rect 13108 64631 13280 64689
rect 13108 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13280 64631
rect 13108 64527 13280 64585
rect 13108 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13280 64527
rect 13108 64423 13280 64481
rect 13108 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13280 64423
rect 13108 64319 13280 64377
rect 13108 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13280 64319
rect 13108 64215 13280 64273
rect 13108 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13280 64215
rect 13108 64111 13280 64169
rect 13108 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13280 64111
rect 13108 64007 13280 64065
rect 13108 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13280 64007
rect 13108 63903 13280 63961
rect 13108 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13280 63903
rect 13108 63799 13280 63857
rect 13108 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13280 63799
rect 13108 63695 13280 63753
rect 13108 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13280 63695
rect 13108 63591 13280 63649
rect 13108 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13280 63591
rect 13108 63487 13280 63545
rect 13108 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13280 63487
rect 13108 63383 13280 63441
rect 13108 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13280 63383
rect 13108 63279 13280 63337
rect 13108 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13280 63279
rect 13108 63175 13280 63233
rect 13108 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13280 63175
rect 13108 63071 13280 63129
rect 13108 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13280 63071
rect 13108 62967 13280 63025
rect 13108 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13280 62967
rect 13108 62863 13280 62921
rect 13108 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13280 62863
rect 13108 62759 13280 62817
rect 13108 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13280 62759
rect 13108 62655 13280 62713
rect 13108 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13280 62655
rect 13108 62551 13280 62609
rect 13108 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13280 62551
rect 13108 62447 13280 62505
rect 13108 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13280 62447
rect 13108 62343 13280 62401
rect 13108 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13280 62343
rect 13108 62239 13280 62297
rect 13108 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13280 62239
rect 13108 62135 13280 62193
rect 13108 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13280 62135
rect 13108 62031 13280 62089
rect 13108 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13280 62031
rect 13108 61927 13280 61985
rect 13108 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13280 61927
rect 13108 61823 13280 61881
rect 13108 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13280 61823
rect 13108 61719 13280 61777
rect 13108 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13280 61719
rect 13108 61615 13280 61673
rect 13108 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13280 61615
rect 13108 61511 13280 61569
rect 13108 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13280 61511
rect 13108 61407 13280 61465
rect 13108 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13280 61407
rect 13108 61303 13280 61361
rect 13108 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13280 61303
rect 13108 61199 13280 61257
rect 13108 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13280 61199
rect 13108 61095 13280 61153
rect 13108 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13280 61095
rect 13108 60991 13280 61049
rect 13108 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13280 60991
rect 13108 60887 13280 60945
rect 13108 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13280 60887
rect 13108 60783 13280 60841
rect 13108 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13280 60783
rect 13108 60679 13280 60737
rect 13108 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13280 60679
rect 13108 60575 13280 60633
rect 13108 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13280 60575
rect 13108 60471 13280 60529
rect 13108 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13280 60471
rect 13108 60367 13280 60425
rect 13108 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13280 60367
rect 13108 60263 13280 60321
rect 13108 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13280 60263
rect 13108 60159 13280 60217
rect 13108 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13280 60159
rect 13108 60055 13280 60113
rect 13108 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13280 60055
rect 13108 59951 13280 60009
rect 13108 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13280 59951
rect 13108 59847 13280 59905
rect 13108 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13280 59847
rect 13108 59743 13280 59801
rect 13108 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13280 59743
rect 13108 59639 13280 59697
rect 13108 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13280 59639
rect 13108 59535 13280 59593
rect 13108 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13280 59535
rect 13108 59431 13280 59489
rect 13108 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13280 59431
rect 13108 59327 13280 59385
rect 13108 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13280 59327
rect 13108 59223 13280 59281
rect 13108 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13280 59223
rect 13108 59119 13280 59177
rect 13108 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13280 59119
rect 13108 59015 13280 59073
rect 13108 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13280 59015
rect 13108 58911 13280 58969
rect 13108 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13280 58911
rect 13108 58807 13280 58865
rect 13108 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13280 58807
rect 13108 58703 13280 58761
rect 13108 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13280 58703
rect 13108 58599 13280 58657
rect 13108 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13280 58599
rect 13108 58495 13280 58553
rect 13108 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13280 58495
rect 13108 58391 13280 58449
rect 13108 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13280 58391
rect 13108 58287 13280 58345
rect 13108 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13280 58287
rect 13108 58183 13280 58241
rect 13108 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13280 58183
rect 13108 58079 13280 58137
rect 13108 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13280 58079
rect 13108 57975 13280 58033
rect 13108 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13280 57975
rect 13108 57871 13280 57929
rect 13108 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13280 57871
rect 13108 57767 13280 57825
rect 13108 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13280 57767
rect 13108 57663 13280 57721
rect 13108 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13280 57663
rect 13108 57559 13280 57617
rect 13108 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13280 57559
rect 13108 57455 13280 57513
rect 13108 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13280 57455
rect 13108 57351 13280 57409
rect 13108 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13280 57351
rect 13108 57247 13280 57305
rect 13108 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13280 57247
rect 13108 57143 13280 57201
rect 13108 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13280 57143
rect 13108 57039 13280 57097
rect 13108 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13280 57039
rect 13108 56935 13280 56993
rect 13108 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13280 56935
rect 13108 56831 13280 56889
rect 13108 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13280 56831
rect 13108 56727 13280 56785
rect 13108 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13280 56727
rect 13108 56623 13280 56681
rect 13108 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13280 56623
rect 13108 56519 13280 56577
rect 13108 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13280 56519
rect 13108 56415 13280 56473
rect 13108 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13280 56415
rect 13108 56311 13280 56369
rect 13108 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13280 56311
rect 13108 56207 13280 56265
rect 13108 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13280 56207
rect 13108 56103 13280 56161
rect 13108 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13280 56103
rect 13108 55999 13280 56057
rect 13108 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13280 55999
rect 13108 55895 13280 55953
rect 13108 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13280 55895
rect 13108 55791 13280 55849
rect 13108 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13280 55791
rect 13108 55687 13280 55745
rect 13108 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13280 55687
rect 13108 55583 13280 55641
rect 13108 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13280 55583
rect 13108 55479 13280 55537
rect 13108 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13280 55479
rect 13108 55375 13280 55433
rect 13108 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13280 55375
rect 13108 55271 13280 55329
rect 13108 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13280 55271
rect 13108 55167 13280 55225
rect 13108 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13280 55167
rect 13108 55063 13280 55121
rect 13108 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13280 55063
rect 13108 54959 13280 55017
rect 13108 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13280 54959
rect 13108 54855 13280 54913
rect 13108 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13280 54855
rect 13108 54751 13280 54809
rect 13108 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13280 54751
rect 13108 54647 13280 54705
rect 13108 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13280 54647
rect 13108 54543 13280 54601
rect 13108 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13280 54543
rect 13108 54439 13280 54497
rect 13108 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13280 54439
rect 13108 54335 13280 54393
rect 13108 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13280 54335
rect 13108 54231 13280 54289
rect 13108 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13280 54231
rect 13108 54127 13280 54185
rect 13108 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13280 54127
rect 13108 54023 13280 54081
rect 13108 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13280 54023
rect 13108 53919 13280 53977
rect 13108 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13280 53919
rect 13108 53815 13280 53873
rect 13108 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13280 53815
rect 13108 53711 13280 53769
rect 13108 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13280 53711
rect 13108 53607 13280 53665
rect 13108 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13280 53607
rect 13108 53503 13280 53561
rect 13108 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13280 53503
rect 13108 53399 13280 53457
rect 13108 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13280 53399
rect 13108 53295 13280 53353
rect 13108 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13280 53295
rect 13108 53191 13280 53249
rect 13108 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13280 53191
rect 13108 53087 13280 53145
rect 13108 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13280 53087
rect 13108 52983 13280 53041
rect 13108 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13280 52983
rect 13108 52879 13280 52937
rect 13108 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13280 52879
rect 13108 52775 13280 52833
rect 13108 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13280 52775
rect 13108 52671 13280 52729
rect 13108 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13280 52671
rect 13108 52567 13280 52625
rect 13108 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13280 52567
rect 13108 52463 13280 52521
rect 13108 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13280 52463
rect 13108 52359 13280 52417
rect 13108 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13280 52359
rect 13108 52255 13280 52313
rect 13108 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13280 52255
rect 13108 52151 13280 52209
rect 13108 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13280 52151
rect 13108 52047 13280 52105
rect 13108 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13280 52047
rect 13108 51943 13280 52001
rect 13108 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13280 51943
rect 13108 51839 13280 51897
rect 13108 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13280 51839
rect 13108 51735 13280 51793
rect 13108 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13280 51735
rect 13108 51631 13280 51689
rect 13108 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13280 51631
rect 13108 51527 13280 51585
rect 13108 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13280 51527
rect 13108 51423 13280 51481
rect 13108 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13280 51423
rect 13108 51319 13280 51377
rect 13108 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13280 51319
rect 13108 51215 13280 51273
rect 13108 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13280 51215
rect 13108 51111 13280 51169
rect 13108 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13280 51111
rect 13108 51007 13280 51065
rect 13108 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13280 51007
rect 13108 50903 13280 50961
rect 13108 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13280 50903
rect 13108 50799 13280 50857
rect 13108 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13280 50799
rect 13108 50695 13280 50753
rect 13108 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13280 50695
rect 13108 50591 13280 50649
rect 13108 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13280 50591
rect 13108 50487 13280 50545
rect 13108 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13280 50487
rect 13108 50383 13280 50441
rect 13108 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13280 50383
rect 13108 50279 13280 50337
rect 13108 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13280 50279
rect 13108 50175 13280 50233
rect 13108 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13280 50175
rect 13108 50071 13280 50129
rect 13108 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13280 50071
rect 13108 49967 13280 50025
rect 13108 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13280 49967
rect 13108 49863 13280 49921
rect 13108 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13280 49863
rect 13108 49759 13280 49817
rect 13108 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13280 49759
rect 13108 49655 13280 49713
rect 13108 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13280 49655
rect 13108 49551 13280 49609
rect 13108 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13280 49551
rect 13108 49447 13280 49505
rect 13108 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13280 49447
rect 13108 49343 13280 49401
rect 13108 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13280 49343
rect 13108 49239 13280 49297
rect 13108 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13280 49239
rect 13108 49135 13280 49193
rect 13108 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13280 49135
rect 13108 49031 13280 49089
rect 13108 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13280 49031
rect 13108 48927 13280 48985
rect 13108 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13280 48927
rect 13108 48823 13280 48881
rect 13108 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13280 48823
rect 13108 48719 13280 48777
rect 13108 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13280 48719
rect 13108 48615 13280 48673
rect 13108 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13280 48615
rect 13108 48511 13280 48569
rect 13108 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13280 48511
rect 13108 48407 13280 48465
rect 13108 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13280 48407
rect 13108 48303 13280 48361
rect 13108 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13280 48303
rect 13108 48199 13280 48257
rect 13108 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13280 48199
rect 13108 48095 13280 48153
rect 13108 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13280 48095
rect 13108 47991 13280 48049
rect 13108 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13280 47991
rect 13108 47887 13280 47945
rect 13108 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13280 47887
rect 13108 47783 13280 47841
rect 13108 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13280 47783
rect 13108 47679 13280 47737
rect 13108 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13280 47679
rect 13108 47575 13280 47633
rect 13108 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13280 47575
rect 13108 47471 13280 47529
rect 13108 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13280 47471
rect 13108 47367 13280 47425
rect 13108 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13280 47367
rect 13108 47263 13280 47321
rect 13108 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13280 47263
rect 13108 47159 13280 47217
rect 13108 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13280 47159
rect 13108 47055 13280 47113
rect 13108 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13280 47055
rect 13108 46951 13280 47009
rect 13108 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13280 46951
rect 13108 46847 13280 46905
rect 13108 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13280 46847
rect 13108 46743 13280 46801
rect 13108 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13280 46743
rect 13108 46639 13280 46697
rect 13108 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13280 46639
rect 13108 46535 13280 46593
rect 13108 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13280 46535
rect 13108 46431 13280 46489
rect 13108 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13280 46431
rect 13108 46327 13280 46385
rect 13108 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13280 46327
rect 13108 46223 13280 46281
rect 13108 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13280 46223
rect 13108 46119 13280 46177
rect 13108 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13280 46119
rect 13108 46015 13280 46073
rect 13108 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13280 46015
rect 13108 45911 13280 45969
rect 13108 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13280 45911
rect 13108 45807 13280 45865
rect 13108 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13280 45807
rect 13108 45703 13280 45761
rect 13108 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13280 45703
rect 13108 45599 13280 45657
rect 13108 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13280 45599
rect 13108 45495 13280 45553
rect 13108 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13280 45495
rect 13108 45391 13280 45449
rect 13108 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13280 45391
rect 13108 45287 13280 45345
rect 13108 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13280 45287
rect 13108 45183 13280 45241
rect 13108 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13280 45183
rect 13108 45079 13280 45137
rect 13108 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13280 45079
rect 13108 44848 13280 45033
rect 70813 69758 70824 69785
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70813 69700 71000 69758
rect 70813 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70813 69596 71000 69654
rect 70813 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70813 69492 71000 69550
rect 70813 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70813 69388 71000 69446
rect 70813 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70813 69284 71000 69342
rect 70813 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70813 69180 71000 69238
rect 70813 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70813 69076 71000 69134
rect 70813 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70813 68972 71000 69030
rect 70813 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70813 68868 71000 68926
rect 70813 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70813 68764 71000 68822
rect 70813 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70813 68660 71000 68718
rect 70813 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70813 68556 71000 68614
rect 70813 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70813 68452 71000 68510
rect 70813 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70813 68348 71000 68406
rect 70813 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70813 68244 71000 68302
rect 70813 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70813 68140 71000 68198
rect 70813 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70813 68036 71000 68094
rect 70813 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70813 67932 71000 67990
rect 70813 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70813 67828 71000 67886
rect 70813 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70813 67724 71000 67782
rect 70813 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70813 67620 71000 67678
rect 70813 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70813 67516 71000 67574
rect 70813 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70813 67412 71000 67470
rect 70813 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70813 67308 71000 67366
rect 70813 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70813 67204 71000 67262
rect 70813 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70813 67100 71000 67158
rect 70813 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70813 66996 71000 67054
rect 70813 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70813 66892 71000 66950
rect 70813 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70813 66788 71000 66846
rect 70813 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70813 66684 71000 66742
rect 70813 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70813 66580 71000 66638
rect 70813 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70813 66476 71000 66534
rect 70813 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70813 66372 71000 66430
rect 70813 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70813 66268 71000 66326
rect 70813 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70813 66164 71000 66222
rect 70813 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70813 66060 71000 66118
rect 70813 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70813 65956 71000 66014
rect 70813 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70813 65852 71000 65910
rect 70813 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70813 65748 71000 65806
rect 70813 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70813 65644 71000 65702
rect 70813 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70813 65540 71000 65598
rect 70813 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70813 65436 71000 65494
rect 70813 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70813 65332 71000 65390
rect 70813 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70813 65228 71000 65286
rect 70813 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70813 65124 71000 65182
rect 70813 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70813 65020 71000 65078
rect 70813 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70813 64916 71000 64974
rect 70813 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70813 64812 71000 64870
rect 70813 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70813 64708 71000 64766
rect 70813 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70813 64604 71000 64662
rect 70813 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70813 64500 71000 64558
rect 70813 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70813 64396 71000 64454
rect 70813 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70813 64292 71000 64350
rect 70813 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70813 64188 71000 64246
rect 70813 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70813 64084 71000 64142
rect 70813 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70813 63980 71000 64038
rect 70813 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70813 63876 71000 63934
rect 70813 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70813 63772 71000 63830
rect 70813 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70813 63668 71000 63726
rect 70813 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70813 63564 71000 63622
rect 70813 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70813 63460 71000 63518
rect 70813 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70813 63356 71000 63414
rect 70813 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70813 63252 71000 63310
rect 70813 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70813 63148 71000 63206
rect 70813 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70813 63044 71000 63102
rect 70813 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70813 62940 71000 62998
rect 70813 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70813 62836 71000 62894
rect 70813 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70813 62732 71000 62790
rect 70813 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70813 62628 71000 62686
rect 70813 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70813 62524 71000 62582
rect 70813 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70813 62420 71000 62478
rect 70813 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70813 62316 71000 62374
rect 70813 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70813 62212 71000 62270
rect 70813 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70813 62108 71000 62166
rect 70813 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70813 62004 71000 62062
rect 70813 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70813 61900 71000 61958
rect 70813 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70813 61796 71000 61854
rect 70813 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70813 61692 71000 61750
rect 70813 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70813 61588 71000 61646
rect 70813 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70813 61484 71000 61542
rect 70813 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70813 61380 71000 61438
rect 70813 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70813 61276 71000 61334
rect 70813 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70813 61172 71000 61230
rect 70813 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70813 61068 71000 61126
rect 70813 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70813 60964 71000 61022
rect 70813 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70813 60860 71000 60918
rect 70813 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70813 60756 71000 60814
rect 70813 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70813 60652 71000 60710
rect 70813 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70813 60548 71000 60606
rect 70813 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70813 60444 71000 60502
rect 70813 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70813 60340 71000 60398
rect 70813 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70813 60236 71000 60294
rect 70813 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70813 60132 71000 60190
rect 70813 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70813 60028 71000 60086
rect 70813 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70813 59924 71000 59982
rect 70813 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70813 59820 71000 59878
rect 70813 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70813 59716 71000 59774
rect 70813 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70813 59612 71000 59670
rect 70813 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70813 59508 71000 59566
rect 70813 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70813 59404 71000 59462
rect 70813 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70813 59300 71000 59358
rect 70813 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70813 59196 71000 59254
rect 70813 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70813 59092 71000 59150
rect 70813 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70813 58988 71000 59046
rect 70813 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70813 58884 71000 58942
rect 70813 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70813 58780 71000 58838
rect 70813 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70813 58676 71000 58734
rect 70813 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70813 58572 71000 58630
rect 70813 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70813 58468 71000 58526
rect 70813 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70813 58364 71000 58422
rect 70813 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70813 58260 71000 58318
rect 70813 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70813 58156 71000 58214
rect 70813 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70813 58052 71000 58110
rect 70813 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70813 57948 71000 58006
rect 70813 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70813 57844 71000 57902
rect 70813 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70813 57740 71000 57798
rect 70813 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70813 57636 71000 57694
rect 70813 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70813 57532 71000 57590
rect 70813 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70813 57428 71000 57486
rect 70813 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70813 57324 71000 57382
rect 70813 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70813 57220 71000 57278
rect 70813 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70813 57116 71000 57174
rect 70813 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70813 57012 71000 57070
rect 70813 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70813 56908 71000 56966
rect 70813 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70813 56804 71000 56862
rect 70813 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70813 56700 71000 56758
rect 70813 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70813 56596 71000 56654
rect 70813 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70813 56492 71000 56550
rect 70813 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70813 56388 71000 56446
rect 70813 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70813 56284 71000 56342
rect 70813 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70813 56180 71000 56238
rect 70813 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70813 56076 71000 56134
rect 70813 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70813 55972 71000 56030
rect 70813 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70813 55868 71000 55926
rect 70813 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70813 55764 71000 55822
rect 70813 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70813 55660 71000 55718
rect 70813 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70813 55556 71000 55614
rect 70813 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70813 55452 71000 55510
rect 70813 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70813 55348 71000 55406
rect 70813 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70813 55244 71000 55302
rect 70813 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70813 55140 71000 55198
rect 70813 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70813 55036 71000 55094
rect 70813 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70813 54932 71000 54990
rect 70813 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70813 54828 71000 54886
rect 70813 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70813 54724 71000 54782
rect 70813 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70813 54620 71000 54678
rect 70813 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70813 54516 71000 54574
rect 70813 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70813 54412 71000 54470
rect 70813 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70813 54308 71000 54366
rect 70813 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70813 54204 71000 54262
rect 70813 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70813 54100 71000 54158
rect 70813 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70813 53996 71000 54054
rect 70813 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70813 53892 71000 53950
rect 70813 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70813 53788 71000 53846
rect 70813 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70813 53684 71000 53742
rect 70813 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70813 53580 71000 53638
rect 70813 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70813 53476 71000 53534
rect 70813 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70813 53372 71000 53430
rect 70813 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70813 53268 71000 53326
rect 70813 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70813 53164 71000 53222
rect 70813 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70813 53060 71000 53118
rect 70813 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70813 52956 71000 53014
rect 70813 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70813 52852 71000 52910
rect 70813 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70813 52748 71000 52806
rect 70813 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70813 52644 71000 52702
rect 70813 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70813 52540 71000 52598
rect 70813 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70813 52436 71000 52494
rect 70813 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70813 52332 71000 52390
rect 70813 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70813 52228 71000 52286
rect 70813 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70813 52124 71000 52182
rect 70813 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70813 52020 71000 52078
rect 70813 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70813 51916 71000 51974
rect 70813 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70813 51812 71000 51870
rect 70813 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70813 51708 71000 51766
rect 70813 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70813 51604 71000 51662
rect 70813 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70813 51500 71000 51558
rect 70813 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70813 51396 71000 51454
rect 70813 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70813 51292 71000 51350
rect 70813 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70813 51188 71000 51246
rect 70813 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70813 51084 71000 51142
rect 70813 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70813 50980 71000 51038
rect 70813 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70813 50876 71000 50934
rect 70813 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70813 50772 71000 50830
rect 70813 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70813 50668 71000 50726
rect 70813 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70813 50564 71000 50622
rect 70813 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70813 50460 71000 50518
rect 70813 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70813 50356 71000 50414
rect 70813 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70813 50252 71000 50310
rect 70813 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70813 50148 71000 50206
rect 70813 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70813 50044 71000 50102
rect 70813 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70813 49940 71000 49998
rect 70813 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70813 49836 71000 49894
rect 70813 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70813 49732 71000 49790
rect 70813 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70813 49628 71000 49686
rect 70813 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70813 49524 71000 49582
rect 70813 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70813 49420 71000 49478
rect 70813 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70813 49316 71000 49374
rect 70813 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70813 49212 71000 49270
rect 70813 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70813 49108 71000 49166
rect 70813 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70813 49004 71000 49062
rect 70813 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70813 48900 71000 48958
rect 70813 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70813 48796 71000 48854
rect 70813 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70813 48692 71000 48750
rect 70813 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70813 48588 71000 48646
rect 70813 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70813 48484 71000 48542
rect 70813 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70813 48380 71000 48438
rect 70813 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70813 48276 71000 48334
rect 70813 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70813 48172 71000 48230
rect 70813 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70813 48068 71000 48126
rect 70813 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70813 47964 71000 48022
rect 70813 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70813 47860 71000 47918
rect 70813 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70813 47756 71000 47814
rect 70813 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70813 47652 71000 47710
rect 70813 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70813 47548 71000 47606
rect 70813 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70813 47444 71000 47502
rect 70813 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70813 47340 71000 47398
rect 70813 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70813 47236 71000 47294
rect 70813 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70813 47132 71000 47190
rect 70813 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70813 47028 71000 47086
rect 70813 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70813 46924 71000 46982
rect 70813 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70813 46820 71000 46878
rect 70813 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70813 46716 71000 46774
rect 70813 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70813 46612 71000 46670
rect 70813 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70813 46508 71000 46566
rect 70813 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70813 46404 71000 46462
rect 70813 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70813 46300 71000 46358
rect 70813 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70813 46196 71000 46254
rect 70813 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70813 46092 71000 46150
rect 70813 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70813 45988 71000 46046
rect 70813 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70813 45884 71000 45942
rect 70813 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70813 45780 71000 45838
rect 70813 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70813 45676 71000 45734
rect 70813 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70813 45572 71000 45630
rect 70813 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70813 45468 71000 45526
rect 70813 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70813 45364 71000 45422
rect 70813 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70813 45260 71000 45318
rect 70813 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70813 45156 71000 45214
rect 70813 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70813 45052 71000 45110
rect 70813 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70813 44948 71000 45006
tri 13108 44703 13253 44848 ne
rect 13253 44828 13280 44848
tri 13280 44828 13372 44920 sw
rect 70813 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 70813 44844 71000 44902
rect 13253 44824 13372 44828
rect 13253 44778 13254 44824
rect 13300 44778 13372 44824
rect 13253 44703 13372 44778
tri 13372 44703 13497 44828 sw
rect 70813 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
rect 70813 44740 71000 44798
tri 13253 44571 13385 44703 ne
rect 13385 44692 13497 44703
rect 13385 44646 13386 44692
rect 13432 44646 13497 44692
rect 13385 44584 13497 44646
tri 13497 44584 13616 44703 sw
rect 70813 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
rect 70813 44636 71000 44694
rect 70813 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
rect 13385 44571 13616 44584
tri 13385 44439 13517 44571 ne
rect 13517 44560 13616 44571
rect 13517 44514 13518 44560
rect 13564 44514 13616 44560
rect 13517 44439 13616 44514
tri 13616 44439 13761 44584 sw
rect 70813 44532 71000 44590
rect 70813 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
tri 13517 44307 13649 44439 ne
rect 13649 44428 13761 44439
rect 13649 44382 13650 44428
rect 13696 44382 13761 44428
rect 13649 44340 13761 44382
tri 13761 44340 13860 44439 sw
rect 70813 44428 71000 44486
rect 70813 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
rect 13649 44307 13860 44340
tri 13649 44175 13781 44307 ne
rect 13781 44296 13860 44307
rect 13781 44250 13782 44296
rect 13828 44250 13860 44296
rect 13781 44175 13860 44250
tri 13860 44175 14025 44340 sw
rect 70813 44324 71000 44382
rect 70813 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
rect 70813 44220 71000 44278
tri 13781 44043 13913 44175 ne
rect 13913 44164 14025 44175
rect 13913 44118 13914 44164
rect 13960 44118 14025 44164
rect 13913 44096 14025 44118
tri 14025 44096 14104 44175 sw
rect 70813 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
rect 70813 44116 71000 44174
rect 13913 44043 14104 44096
tri 13913 43911 14045 44043 ne
rect 14045 44032 14104 44043
rect 14045 43986 14046 44032
rect 14092 43986 14104 44032
rect 14045 43911 14104 43986
tri 14104 43911 14289 44096 sw
rect 70813 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
rect 70813 44012 71000 44070
rect 70813 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
tri 14045 43779 14177 43911 ne
rect 14177 43900 14289 43911
rect 14177 43854 14178 43900
rect 14224 43854 14289 43900
rect 14177 43779 14289 43854
tri 14289 43779 14421 43911 sw
rect 70813 43908 71000 43966
rect 70813 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
rect 70813 43804 71000 43862
tri 14177 43647 14309 43779 ne
rect 14309 43768 14421 43779
rect 14309 43722 14310 43768
rect 14356 43722 14421 43768
rect 14309 43647 14421 43722
tri 14421 43647 14553 43779 sw
rect 70813 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 70813 43700 71000 43758
rect 70813 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
tri 14309 43515 14441 43647 ne
rect 14441 43636 14553 43647
rect 14441 43590 14442 43636
rect 14488 43590 14553 43636
rect 14441 43515 14553 43590
tri 14553 43515 14685 43647 sw
rect 70813 43596 71000 43654
rect 70813 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
tri 14441 43383 14573 43515 ne
rect 14573 43504 14685 43515
rect 14573 43458 14574 43504
rect 14620 43458 14685 43504
rect 14573 43383 14685 43458
tri 14685 43383 14817 43515 sw
rect 70813 43492 71000 43550
rect 70813 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
rect 70813 43388 71000 43446
tri 14573 43251 14705 43383 ne
rect 14705 43372 14817 43383
rect 14705 43326 14706 43372
rect 14752 43326 14817 43372
rect 14705 43251 14817 43326
tri 14817 43251 14949 43383 sw
rect 70813 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
rect 70813 43284 71000 43342
tri 14705 43119 14837 43251 ne
rect 14837 43240 14949 43251
rect 14837 43194 14838 43240
rect 14884 43194 14949 43240
rect 14837 43120 14949 43194
tri 14949 43120 15080 43251 sw
rect 70813 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 70813 43180 71000 43238
rect 70813 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
rect 14837 43119 15080 43120
tri 14837 42987 14969 43119 ne
rect 14969 43108 15080 43119
rect 14969 43062 14970 43108
rect 15016 43062 15080 43108
rect 14969 42987 15080 43062
tri 15080 42987 15213 43120 sw
rect 70813 43076 71000 43134
rect 70813 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
tri 14969 42855 15101 42987 ne
rect 15101 42976 15213 42987
rect 15101 42930 15102 42976
rect 15148 42930 15213 42976
rect 15101 42876 15213 42930
tri 15213 42876 15324 42987 sw
rect 70813 42972 71000 43030
rect 70813 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
rect 15101 42855 15324 42876
tri 15101 42723 15233 42855 ne
rect 15233 42844 15324 42855
rect 15233 42798 15234 42844
rect 15280 42798 15324 42844
rect 15233 42723 15324 42798
tri 15324 42723 15477 42876 sw
rect 70813 42868 71000 42926
rect 70813 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
rect 70813 42764 71000 42822
tri 15233 42591 15365 42723 ne
rect 15365 42712 15477 42723
rect 15365 42666 15366 42712
rect 15412 42666 15477 42712
rect 15365 42632 15477 42666
tri 15477 42632 15568 42723 sw
rect 70813 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
rect 70813 42660 71000 42718
rect 15365 42591 15568 42632
tri 15365 42459 15497 42591 ne
rect 15497 42580 15568 42591
rect 15497 42534 15498 42580
rect 15544 42534 15568 42580
rect 15497 42459 15568 42534
tri 15568 42459 15741 42632 sw
rect 70813 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
rect 70813 42556 71000 42614
rect 70813 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
tri 15497 42327 15629 42459 ne
rect 15629 42448 15741 42459
rect 15629 42402 15630 42448
rect 15676 42402 15741 42448
rect 15629 42327 15741 42402
tri 15741 42327 15873 42459 sw
rect 70813 42452 71000 42510
rect 70813 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
rect 70813 42348 71000 42406
tri 15629 42195 15761 42327 ne
rect 15761 42316 15873 42327
rect 15761 42270 15762 42316
rect 15808 42270 15873 42316
rect 15761 42195 15873 42270
tri 15873 42195 16005 42327 sw
rect 70813 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 70813 42244 71000 42302
rect 70813 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
tri 15761 42063 15893 42195 ne
rect 15893 42184 16005 42195
rect 15893 42138 15894 42184
rect 15940 42138 16005 42184
rect 15893 42063 16005 42138
tri 16005 42063 16137 42195 sw
rect 70813 42140 71000 42198
rect 70813 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
tri 15893 41931 16025 42063 ne
rect 16025 42052 16137 42063
rect 16025 42006 16026 42052
rect 16072 42006 16137 42052
rect 16025 41931 16137 42006
tri 16137 41931 16269 42063 sw
rect 70813 42036 71000 42094
rect 70813 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
rect 70813 41932 71000 41990
tri 16025 41799 16157 41931 ne
rect 16157 41920 16269 41931
rect 16157 41874 16158 41920
rect 16204 41874 16269 41920
rect 16157 41799 16269 41874
tri 16269 41799 16401 41931 sw
rect 70813 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
rect 70813 41828 71000 41886
tri 16157 41667 16289 41799 ne
rect 16289 41788 16401 41799
rect 16289 41742 16290 41788
rect 16336 41742 16401 41788
rect 16289 41667 16401 41742
tri 16289 41599 16357 41667 ne
rect 16357 41656 16401 41667
tri 16401 41656 16544 41799 sw
rect 70813 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 70813 41724 71000 41782
rect 70813 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
rect 16357 41610 16422 41656
rect 16468 41610 16544 41656
rect 16357 41599 16544 41610
tri 16357 41412 16544 41599 ne
tri 16544 41535 16665 41656 sw
rect 70813 41620 71000 41678
rect 70813 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
rect 16544 41524 16665 41535
rect 16544 41478 16554 41524
rect 16600 41478 16665 41524
rect 16544 41412 16665 41478
tri 16665 41412 16788 41535 sw
rect 70813 41516 71000 41574
rect 70813 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
rect 70813 41412 71000 41470
tri 16544 41271 16685 41412 ne
rect 16685 41392 16788 41412
rect 16685 41346 16686 41392
rect 16732 41346 16788 41392
rect 16685 41271 16788 41346
tri 16788 41271 16929 41412 sw
rect 70813 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
rect 70813 41308 71000 41366
tri 16685 41139 16817 41271 ne
rect 16817 41260 16929 41271
rect 16817 41214 16818 41260
rect 16864 41214 16929 41260
rect 16817 41168 16929 41214
tri 16929 41168 17032 41271 sw
rect 70813 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
rect 70813 41204 71000 41262
rect 16817 41139 17032 41168
tri 16817 41007 16949 41139 ne
rect 16949 41128 17032 41139
rect 16949 41082 16950 41128
rect 16996 41082 17032 41128
rect 16949 41007 17032 41082
tri 17032 41007 17193 41168 sw
rect 70813 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
rect 70813 41100 71000 41158
rect 70813 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
tri 16949 40875 17081 41007 ne
rect 17081 40996 17193 41007
rect 17081 40950 17082 40996
rect 17128 40950 17193 40996
rect 17081 40924 17193 40950
tri 17193 40924 17276 41007 sw
rect 70813 40996 71000 41054
rect 70813 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
rect 17081 40875 17276 40924
tri 17081 40743 17213 40875 ne
rect 17213 40864 17276 40875
rect 17213 40818 17214 40864
rect 17260 40818 17276 40864
rect 17213 40743 17276 40818
tri 17276 40743 17457 40924 sw
rect 70813 40892 71000 40950
rect 70813 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 70813 40788 71000 40846
tri 17213 40611 17345 40743 ne
rect 17345 40732 17457 40743
rect 17345 40686 17346 40732
rect 17392 40686 17457 40732
rect 17345 40611 17457 40686
tri 17457 40611 17589 40743 sw
rect 70813 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
rect 70813 40684 71000 40742
rect 70813 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
tri 17345 40479 17477 40611 ne
rect 17477 40600 17589 40611
rect 17477 40554 17478 40600
rect 17524 40554 17589 40600
rect 17477 40479 17589 40554
tri 17589 40479 17721 40611 sw
rect 70813 40580 71000 40638
rect 70813 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
tri 17477 40347 17609 40479 ne
rect 17609 40468 17721 40479
rect 17609 40422 17610 40468
rect 17656 40422 17721 40468
rect 17609 40347 17721 40422
tri 17721 40347 17853 40479 sw
rect 70813 40476 71000 40534
rect 70813 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
rect 70813 40372 71000 40430
tri 17609 40215 17741 40347 ne
rect 17741 40336 17853 40347
rect 17741 40290 17742 40336
rect 17788 40290 17853 40336
rect 17741 40215 17853 40290
tri 17853 40215 17985 40347 sw
rect 70813 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 70813 40268 71000 40326
rect 70813 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
tri 17741 40083 17873 40215 ne
rect 17873 40204 17985 40215
rect 17873 40158 17874 40204
rect 17920 40158 17985 40204
rect 17873 40083 17985 40158
tri 17985 40083 18117 40215 sw
rect 70813 40164 71000 40222
rect 70813 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
tri 17873 39951 18005 40083 ne
rect 18005 40072 18117 40083
rect 18005 40026 18006 40072
rect 18052 40026 18117 40072
rect 18005 39951 18117 40026
tri 18005 39883 18073 39951 ne
rect 18073 39948 18117 39951
tri 18117 39948 18252 40083 sw
rect 70813 40060 71000 40118
rect 70813 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
rect 70813 39956 71000 40014
rect 18073 39940 18252 39948
rect 18073 39894 18138 39940
rect 18184 39894 18252 39940
rect 18073 39883 18252 39894
tri 18073 39704 18252 39883 ne
tri 18252 39819 18381 39948 sw
rect 70813 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
rect 70813 39852 71000 39910
rect 18252 39808 18381 39819
rect 18252 39762 18270 39808
rect 18316 39762 18381 39808
rect 18252 39704 18381 39762
tri 18381 39704 18496 39819 sw
rect 70813 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 70813 39748 71000 39806
tri 18252 39555 18401 39704 ne
rect 18401 39676 18496 39704
rect 18401 39630 18402 39676
rect 18448 39630 18496 39676
rect 18401 39555 18496 39630
tri 18496 39555 18645 39704 sw
rect 70813 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
rect 70813 39644 71000 39702
rect 70813 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
tri 18401 39423 18533 39555 ne
rect 18533 39544 18645 39555
rect 18533 39498 18534 39544
rect 18580 39498 18645 39544
rect 18533 39460 18645 39498
tri 18645 39460 18740 39555 sw
rect 70813 39540 71000 39598
rect 70813 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
rect 18533 39423 18740 39460
tri 18533 39291 18665 39423 ne
rect 18665 39412 18740 39423
rect 18665 39366 18666 39412
rect 18712 39366 18740 39412
rect 18665 39291 18740 39366
tri 18740 39291 18909 39460 sw
rect 70813 39436 71000 39494
rect 70813 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
rect 70813 39332 71000 39390
tri 18665 39159 18797 39291 ne
rect 18797 39280 18909 39291
rect 18797 39234 18798 39280
rect 18844 39234 18909 39280
rect 18797 39159 18909 39234
tri 18909 39159 19041 39291 sw
rect 70813 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
rect 70813 39228 71000 39286
rect 70813 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
tri 18797 39027 18929 39159 ne
rect 18929 39148 19041 39159
rect 18929 39102 18930 39148
rect 18976 39102 19041 39148
rect 18929 39027 19041 39102
tri 19041 39027 19173 39159 sw
rect 70813 39124 71000 39182
rect 70813 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
tri 18929 38895 19061 39027 ne
rect 19061 39016 19173 39027
rect 19061 38970 19062 39016
rect 19108 38970 19173 39016
rect 19061 38895 19173 38970
tri 19173 38895 19305 39027 sw
rect 70813 39020 71000 39078
rect 70813 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
rect 70813 38916 71000 38974
tri 19061 38763 19193 38895 ne
rect 19193 38884 19305 38895
rect 19193 38838 19194 38884
rect 19240 38838 19305 38884
rect 19193 38763 19305 38838
tri 19305 38763 19437 38895 sw
rect 70813 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 70813 38812 71000 38870
rect 70813 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
tri 19193 38631 19325 38763 ne
rect 19325 38752 19437 38763
rect 19325 38706 19326 38752
rect 19372 38706 19437 38752
rect 19325 38631 19437 38706
tri 19437 38631 19569 38763 sw
rect 70813 38708 71000 38766
rect 70813 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
tri 19325 38499 19457 38631 ne
rect 19457 38620 19569 38631
rect 19457 38574 19458 38620
rect 19504 38574 19569 38620
rect 19457 38499 19569 38574
tri 19569 38499 19701 38631 sw
rect 70813 38604 71000 38662
rect 70813 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
rect 70813 38500 71000 38558
tri 19457 38367 19589 38499 ne
rect 19589 38488 19701 38499
rect 19589 38442 19590 38488
rect 19636 38442 19701 38488
rect 19589 38367 19701 38442
tri 19701 38367 19833 38499 sw
rect 70813 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 70813 38396 71000 38454
tri 19589 38235 19721 38367 ne
rect 19721 38356 19833 38367
rect 19721 38310 19722 38356
rect 19768 38310 19833 38356
rect 19721 38240 19833 38310
tri 19833 38240 19960 38367 sw
rect 70813 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
rect 70813 38292 71000 38350
rect 70813 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
rect 19721 38235 19960 38240
tri 19721 38103 19853 38235 ne
rect 19853 38224 19960 38235
rect 19853 38178 19854 38224
rect 19900 38178 19960 38224
rect 19853 38103 19960 38178
tri 19960 38103 20097 38240 sw
rect 70813 38188 71000 38246
rect 70813 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
tri 19853 37971 19985 38103 ne
rect 19985 38092 20097 38103
rect 19985 38046 19986 38092
rect 20032 38046 20097 38092
rect 19985 37996 20097 38046
tri 20097 37996 20204 38103 sw
rect 70813 38084 71000 38142
rect 70813 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
rect 19985 37971 20204 37996
tri 19985 37839 20117 37971 ne
rect 20117 37960 20204 37971
rect 20117 37914 20118 37960
rect 20164 37914 20204 37960
rect 20117 37839 20204 37914
tri 20204 37839 20361 37996 sw
rect 70813 37980 71000 38038
rect 70813 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
rect 70813 37876 71000 37934
tri 20117 37707 20249 37839 ne
rect 20249 37828 20361 37839
rect 20249 37782 20250 37828
rect 20296 37782 20361 37828
rect 20249 37752 20361 37782
tri 20361 37752 20448 37839 sw
rect 70813 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
rect 70813 37772 71000 37830
rect 20249 37707 20448 37752
tri 20249 37575 20381 37707 ne
rect 20381 37696 20448 37707
rect 20381 37650 20382 37696
rect 20428 37650 20448 37696
rect 20381 37575 20448 37650
tri 20448 37575 20625 37752 sw
rect 70813 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
rect 70813 37668 71000 37726
rect 70813 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
tri 20381 37443 20513 37575 ne
rect 20513 37564 20625 37575
rect 20513 37518 20514 37564
rect 20560 37518 20625 37564
rect 20513 37443 20625 37518
tri 20625 37443 20757 37575 sw
rect 70813 37564 71000 37622
rect 70813 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
rect 70813 37460 71000 37518
tri 20513 37311 20645 37443 ne
rect 20645 37432 20757 37443
rect 20645 37386 20646 37432
rect 20692 37386 20757 37432
rect 20645 37311 20757 37386
tri 20757 37311 20889 37443 sw
rect 70813 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
rect 70813 37356 71000 37414
tri 20645 37179 20777 37311 ne
rect 20777 37300 20889 37311
rect 20777 37254 20778 37300
rect 20824 37254 20889 37300
rect 20777 37179 20889 37254
tri 20889 37179 21021 37311 sw
rect 70813 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
rect 70813 37252 71000 37310
rect 70813 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
tri 20777 37047 20909 37179 ne
rect 20909 37168 21021 37179
rect 20909 37122 20910 37168
rect 20956 37122 21021 37168
rect 20909 37047 21021 37122
tri 21021 37047 21153 37179 sw
rect 70813 37148 71000 37206
rect 70813 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
tri 20909 36915 21041 37047 ne
rect 21041 37036 21153 37047
rect 21041 36990 21042 37036
rect 21088 36990 21153 37036
rect 21041 36915 21153 36990
tri 21153 36915 21285 37047 sw
rect 70813 37044 71000 37102
rect 70813 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
rect 70813 36940 71000 36998
tri 21041 36783 21173 36915 ne
rect 21173 36904 21285 36915
rect 21173 36858 21174 36904
rect 21220 36858 21285 36904
rect 21173 36783 21285 36858
tri 21173 36715 21241 36783 ne
rect 21241 36776 21285 36783
tri 21285 36776 21424 36915 sw
rect 70813 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
rect 70813 36836 71000 36894
rect 70813 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
rect 21241 36772 21424 36776
rect 21241 36726 21306 36772
rect 21352 36726 21424 36772
rect 21241 36715 21424 36726
tri 21241 36532 21424 36715 ne
tri 21424 36651 21549 36776 sw
rect 70813 36732 71000 36790
rect 70813 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
rect 21424 36640 21549 36651
rect 21424 36594 21438 36640
rect 21484 36594 21549 36640
rect 21424 36532 21549 36594
tri 21549 36532 21668 36651 sw
rect 70813 36628 71000 36686
rect 70813 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
tri 21424 36387 21569 36532 ne
rect 21569 36508 21668 36532
rect 21569 36462 21570 36508
rect 21616 36462 21668 36508
rect 21569 36387 21668 36462
tri 21668 36387 21813 36532 sw
rect 70813 36524 71000 36582
rect 70813 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
rect 70813 36420 71000 36478
tri 21569 36255 21701 36387 ne
rect 21701 36376 21813 36387
rect 21701 36330 21702 36376
rect 21748 36330 21813 36376
rect 21701 36288 21813 36330
tri 21813 36288 21912 36387 sw
rect 70813 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 70813 36316 71000 36374
rect 21701 36255 21912 36288
tri 21701 36123 21833 36255 ne
rect 21833 36244 21912 36255
rect 21833 36198 21834 36244
rect 21880 36198 21912 36244
rect 21833 36123 21912 36198
tri 21912 36123 22077 36288 sw
rect 70813 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
rect 70813 36212 71000 36270
rect 70813 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
tri 21833 35991 21965 36123 ne
rect 21965 36112 22077 36123
rect 21965 36066 21966 36112
rect 22012 36066 22077 36112
rect 21965 36044 22077 36066
tri 22077 36044 22156 36123 sw
rect 70813 36108 71000 36166
rect 70813 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
rect 21965 35991 22156 36044
tri 21965 35859 22097 35991 ne
rect 22097 35980 22156 35991
rect 22097 35934 22098 35980
rect 22144 35934 22156 35980
rect 22097 35859 22156 35934
tri 22156 35859 22341 36044 sw
rect 70813 36004 71000 36062
rect 70813 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 70813 35900 71000 35958
tri 22097 35727 22229 35859 ne
rect 22229 35848 22341 35859
rect 22229 35802 22230 35848
rect 22276 35802 22341 35848
rect 22229 35727 22341 35802
tri 22341 35727 22473 35859 sw
rect 70813 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
rect 70813 35796 71000 35854
rect 70813 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
tri 22229 35595 22361 35727 ne
rect 22361 35716 22473 35727
rect 22361 35670 22362 35716
rect 22408 35670 22473 35716
rect 22361 35595 22473 35670
tri 22473 35595 22605 35727 sw
rect 70813 35692 71000 35750
rect 70813 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
tri 22361 35463 22493 35595 ne
rect 22493 35584 22605 35595
rect 22493 35538 22494 35584
rect 22540 35538 22605 35584
rect 22493 35463 22605 35538
tri 22605 35463 22737 35595 sw
rect 70813 35588 71000 35646
rect 70813 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
rect 70813 35484 71000 35542
tri 22493 35331 22625 35463 ne
rect 22625 35452 22737 35463
rect 22625 35406 22626 35452
rect 22672 35406 22737 35452
rect 22625 35331 22737 35406
tri 22737 35331 22869 35463 sw
rect 70813 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 70813 35380 71000 35438
rect 70813 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
tri 22625 35199 22757 35331 ne
rect 22757 35320 22869 35331
rect 22757 35274 22758 35320
rect 22804 35274 22869 35320
rect 22757 35199 22869 35274
tri 22869 35199 23001 35331 sw
rect 70813 35276 71000 35334
rect 70813 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
tri 22757 35067 22889 35199 ne
rect 22889 35188 23001 35199
rect 22889 35142 22890 35188
rect 22936 35142 23001 35188
rect 22889 35068 23001 35142
tri 23001 35068 23132 35199 sw
rect 70813 35172 71000 35230
rect 70813 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
rect 70813 35068 71000 35126
rect 22889 35067 23132 35068
tri 22889 34935 23021 35067 ne
rect 23021 35056 23132 35067
rect 23021 35010 23022 35056
rect 23068 35010 23132 35056
rect 23021 34935 23132 35010
tri 23132 34935 23265 35068 sw
rect 70813 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
rect 70813 34964 71000 35022
tri 23021 34803 23153 34935 ne
rect 23153 34924 23265 34935
rect 23153 34878 23154 34924
rect 23200 34878 23265 34924
rect 23153 34824 23265 34878
tri 23265 34824 23376 34935 sw
rect 70813 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 70813 34860 71000 34918
rect 23153 34803 23376 34824
tri 23153 34671 23285 34803 ne
rect 23285 34792 23376 34803
rect 23285 34746 23286 34792
rect 23332 34746 23376 34792
rect 23285 34671 23376 34746
tri 23376 34671 23529 34824 sw
rect 70813 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
rect 70813 34756 71000 34814
rect 70813 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
tri 23285 34539 23417 34671 ne
rect 23417 34660 23529 34671
rect 23417 34614 23418 34660
rect 23464 34614 23529 34660
rect 23417 34580 23529 34614
tri 23529 34580 23620 34671 sw
rect 70813 34652 71000 34710
rect 70813 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
rect 23417 34539 23620 34580
tri 23417 34407 23549 34539 ne
rect 23549 34528 23620 34539
rect 23549 34482 23550 34528
rect 23596 34482 23620 34528
rect 23549 34407 23620 34482
tri 23620 34407 23793 34580 sw
rect 70813 34548 71000 34606
rect 70813 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
rect 70813 34444 71000 34502
tri 23549 34275 23681 34407 ne
rect 23681 34396 23793 34407
rect 23681 34350 23682 34396
rect 23728 34350 23793 34396
rect 23681 34275 23793 34350
tri 23793 34275 23925 34407 sw
rect 70813 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
rect 70813 34340 71000 34398
rect 70813 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
tri 23681 34143 23813 34275 ne
rect 23813 34264 23925 34275
rect 23813 34218 23814 34264
rect 23860 34218 23925 34264
rect 23813 34143 23925 34218
tri 23925 34143 24057 34275 sw
rect 70813 34236 71000 34294
rect 70813 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
tri 23813 34011 23945 34143 ne
rect 23945 34132 24057 34143
rect 23945 34086 23946 34132
rect 23992 34086 24057 34132
rect 23945 34011 24057 34086
tri 24057 34011 24189 34143 sw
rect 70813 34132 71000 34190
rect 70813 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
rect 70813 34028 71000 34086
tri 23945 33879 24077 34011 ne
rect 24077 34000 24189 34011
rect 24077 33954 24078 34000
rect 24124 33954 24189 34000
rect 24077 33879 24189 33954
tri 24189 33879 24321 34011 sw
rect 70813 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 70813 33924 71000 33982
tri 24077 33747 24209 33879 ne
rect 24209 33868 24321 33879
rect 24209 33822 24210 33868
rect 24256 33822 24321 33868
rect 24209 33747 24321 33822
tri 24321 33747 24453 33879 sw
rect 70813 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
rect 70813 33820 71000 33878
rect 70813 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
tri 24209 33615 24341 33747 ne
rect 24341 33736 24453 33747
rect 24341 33690 24342 33736
rect 24388 33690 24453 33736
rect 24341 33615 24453 33690
tri 24341 33547 24409 33615 ne
rect 24409 33604 24453 33615
tri 24453 33604 24596 33747 sw
rect 70813 33716 71000 33774
rect 70813 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
rect 70813 33612 71000 33670
rect 24409 33558 24474 33604
rect 24520 33558 24596 33604
rect 24409 33547 24596 33558
tri 24409 33360 24596 33547 ne
tri 24596 33483 24717 33604 sw
rect 70813 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
rect 70813 33508 71000 33566
rect 24596 33472 24717 33483
rect 24596 33426 24606 33472
rect 24652 33426 24717 33472
rect 24596 33360 24717 33426
tri 24717 33360 24840 33483 sw
rect 70813 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 70813 33404 71000 33462
tri 24596 33219 24737 33360 ne
rect 24737 33340 24840 33360
rect 24737 33294 24738 33340
rect 24784 33294 24840 33340
rect 24737 33219 24840 33294
tri 24840 33219 24981 33360 sw
rect 70813 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
rect 70813 33300 71000 33358
rect 70813 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
tri 24737 33087 24869 33219 ne
rect 24869 33208 24981 33219
rect 24869 33162 24870 33208
rect 24916 33162 24981 33208
rect 24869 33116 24981 33162
tri 24981 33116 25084 33219 sw
rect 70813 33196 71000 33254
rect 70813 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
rect 24869 33087 25084 33116
tri 24869 32955 25001 33087 ne
rect 25001 33076 25084 33087
rect 25001 33030 25002 33076
rect 25048 33030 25084 33076
rect 25001 32955 25084 33030
tri 25084 32955 25245 33116 sw
rect 70813 33092 71000 33150
rect 70813 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
rect 70813 32988 71000 33046
tri 25001 32823 25133 32955 ne
rect 25133 32944 25245 32955
rect 25133 32898 25134 32944
rect 25180 32898 25245 32944
rect 25133 32872 25245 32898
tri 25245 32872 25328 32955 sw
rect 70813 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 70813 32884 71000 32942
rect 25133 32823 25328 32872
tri 25133 32691 25265 32823 ne
rect 25265 32812 25328 32823
rect 25265 32766 25266 32812
rect 25312 32766 25328 32812
rect 25265 32691 25328 32766
tri 25328 32691 25509 32872 sw
rect 70813 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
rect 70813 32780 71000 32838
rect 70813 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
tri 25265 32559 25397 32691 ne
rect 25397 32680 25509 32691
rect 25397 32634 25398 32680
rect 25444 32634 25509 32680
rect 25397 32559 25509 32634
tri 25509 32559 25641 32691 sw
rect 70813 32676 71000 32734
rect 70813 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
rect 70813 32572 71000 32630
tri 25397 32427 25529 32559 ne
rect 25529 32548 25641 32559
rect 25529 32502 25530 32548
rect 25576 32502 25641 32548
rect 25529 32427 25641 32502
tri 25641 32427 25773 32559 sw
rect 70813 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
rect 70813 32468 71000 32526
tri 25529 32295 25661 32427 ne
rect 25661 32416 25773 32427
rect 25661 32370 25662 32416
rect 25708 32370 25773 32416
rect 25661 32295 25773 32370
tri 25773 32295 25905 32427 sw
rect 70813 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
rect 70813 32364 71000 32422
rect 70813 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
tri 25661 32163 25793 32295 ne
rect 25793 32284 25905 32295
rect 25793 32238 25794 32284
rect 25840 32238 25905 32284
rect 25793 32163 25905 32238
tri 25905 32163 26037 32295 sw
rect 70813 32260 71000 32318
rect 70813 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
tri 25793 32031 25925 32163 ne
rect 25925 32152 26037 32163
rect 25925 32106 25926 32152
rect 25972 32106 26037 32152
rect 25925 32031 26037 32106
tri 26037 32031 26169 32163 sw
rect 70813 32156 71000 32214
rect 70813 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
rect 70813 32052 71000 32110
tri 25925 31899 26057 32031 ne
rect 26057 32020 26169 32031
rect 26057 31974 26058 32020
rect 26104 31974 26169 32020
rect 26057 31899 26169 31974
tri 26057 31831 26125 31899 ne
rect 26125 31896 26169 31899
tri 26169 31896 26304 32031 sw
rect 70813 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 70813 31948 71000 32006
rect 70813 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
rect 26125 31888 26304 31896
rect 26125 31842 26190 31888
rect 26236 31842 26304 31888
rect 26125 31831 26304 31842
tri 26125 31652 26304 31831 ne
tri 26304 31767 26433 31896 sw
rect 70813 31844 71000 31902
rect 70813 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
rect 26304 31756 26433 31767
rect 26304 31710 26322 31756
rect 26368 31710 26433 31756
rect 26304 31652 26433 31710
tri 26433 31652 26548 31767 sw
rect 70813 31740 71000 31798
rect 70813 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
tri 26304 31503 26453 31652 ne
rect 26453 31624 26548 31652
rect 26453 31578 26454 31624
rect 26500 31578 26548 31624
rect 26453 31503 26548 31578
tri 26548 31503 26697 31652 sw
rect 70813 31636 71000 31694
rect 70813 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
rect 70813 31532 71000 31590
tri 26453 31371 26585 31503 ne
rect 26585 31492 26697 31503
rect 26585 31446 26586 31492
rect 26632 31446 26697 31492
rect 26585 31408 26697 31446
tri 26697 31408 26792 31503 sw
rect 70813 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 70813 31428 71000 31486
rect 26585 31371 26792 31408
tri 26585 31239 26717 31371 ne
rect 26717 31360 26792 31371
rect 26717 31314 26718 31360
rect 26764 31314 26792 31360
rect 26717 31239 26792 31314
tri 26792 31239 26961 31408 sw
rect 70813 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
rect 70813 31324 71000 31382
rect 70813 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
tri 26717 31107 26849 31239 ne
rect 26849 31228 26961 31239
rect 26849 31182 26850 31228
rect 26896 31182 26961 31228
rect 26849 31107 26961 31182
tri 26961 31107 27093 31239 sw
rect 70813 31220 71000 31278
rect 70813 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
rect 70813 31116 71000 31174
tri 26849 30975 26981 31107 ne
rect 26981 31096 27093 31107
rect 26981 31050 26982 31096
rect 27028 31050 27093 31096
rect 26981 30975 27093 31050
tri 27093 30975 27225 31107 sw
rect 70813 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
rect 70813 31012 71000 31070
tri 26981 30843 27113 30975 ne
rect 27113 30964 27225 30975
rect 27113 30918 27114 30964
rect 27160 30918 27225 30964
rect 27113 30843 27225 30918
tri 27225 30843 27357 30975 sw
rect 70813 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
rect 70813 30908 71000 30966
rect 70813 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
tri 27113 30711 27245 30843 ne
rect 27245 30832 27357 30843
rect 27245 30786 27246 30832
rect 27292 30786 27357 30832
rect 27245 30711 27357 30786
tri 27357 30711 27489 30843 sw
rect 70813 30804 71000 30862
rect 70813 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
tri 27245 30579 27377 30711 ne
rect 27377 30700 27489 30711
rect 27377 30654 27378 30700
rect 27424 30654 27489 30700
rect 27377 30579 27489 30654
tri 27489 30579 27621 30711 sw
rect 70813 30700 71000 30758
rect 70813 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
rect 70813 30596 71000 30654
tri 27377 30447 27509 30579 ne
rect 27509 30568 27621 30579
rect 27509 30522 27510 30568
rect 27556 30522 27621 30568
rect 27509 30447 27621 30522
tri 27621 30447 27753 30579 sw
rect 70813 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 70813 30492 71000 30550
tri 27509 30315 27641 30447 ne
rect 27641 30436 27753 30447
rect 27641 30390 27642 30436
rect 27688 30390 27753 30436
rect 27641 30315 27753 30390
tri 27753 30315 27885 30447 sw
rect 70813 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
rect 70813 30388 71000 30446
rect 70813 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
tri 27641 30183 27773 30315 ne
rect 27773 30304 27885 30315
rect 27773 30258 27774 30304
rect 27820 30258 27885 30304
rect 27773 30188 27885 30258
tri 27885 30188 28012 30315 sw
rect 70813 30284 71000 30342
rect 70813 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
rect 27773 30183 28012 30188
tri 27773 30051 27905 30183 ne
rect 27905 30172 28012 30183
rect 27905 30126 27906 30172
rect 27952 30126 28012 30172
rect 27905 30051 28012 30126
tri 28012 30051 28149 30188 sw
rect 70813 30180 71000 30238
rect 70813 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
rect 70813 30076 71000 30134
tri 27905 29919 28037 30051 ne
rect 28037 30040 28149 30051
rect 28037 29994 28038 30040
rect 28084 29994 28149 30040
rect 28037 29944 28149 29994
tri 28149 29944 28256 30051 sw
rect 70813 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 70813 29972 71000 30030
rect 28037 29919 28256 29944
tri 28037 29787 28169 29919 ne
rect 28169 29908 28256 29919
rect 28169 29862 28170 29908
rect 28216 29862 28256 29908
rect 28169 29787 28256 29862
tri 28256 29787 28413 29944 sw
rect 70813 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
rect 70813 29868 71000 29926
rect 70813 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
tri 28169 29655 28301 29787 ne
rect 28301 29776 28413 29787
rect 28301 29730 28302 29776
rect 28348 29730 28413 29776
rect 28301 29700 28413 29730
tri 28413 29700 28500 29787 sw
rect 70813 29764 71000 29822
rect 70813 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
rect 28301 29655 28500 29700
tri 28301 29523 28433 29655 ne
rect 28433 29644 28500 29655
rect 28433 29598 28434 29644
rect 28480 29598 28500 29644
rect 28433 29523 28500 29598
tri 28500 29523 28677 29700 sw
rect 70813 29660 71000 29718
rect 70813 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
rect 70813 29556 71000 29614
tri 28433 29391 28565 29523 ne
rect 28565 29512 28677 29523
rect 28565 29466 28566 29512
rect 28612 29466 28677 29512
rect 28565 29391 28677 29466
tri 28677 29391 28809 29523 sw
rect 70813 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 70813 29452 71000 29510
rect 70813 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
tri 28565 29259 28697 29391 ne
rect 28697 29380 28809 29391
rect 28697 29334 28698 29380
rect 28744 29334 28809 29380
rect 28697 29259 28809 29334
tri 28809 29259 28941 29391 sw
rect 70813 29348 71000 29406
rect 70813 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
tri 28697 29127 28829 29259 ne
rect 28829 29248 28941 29259
rect 28829 29202 28830 29248
rect 28876 29202 28941 29248
rect 28829 29127 28941 29202
tri 28941 29127 29073 29259 sw
rect 70813 29244 71000 29302
rect 70813 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
rect 70813 29140 71000 29198
tri 28829 28995 28961 29127 ne
rect 28961 29116 29073 29127
rect 28961 29070 28962 29116
rect 29008 29070 29073 29116
rect 28961 28995 29073 29070
tri 29073 28995 29205 29127 sw
rect 70813 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
rect 70813 29036 71000 29094
tri 28961 28863 29093 28995 ne
rect 29093 28984 29205 28995
rect 29093 28938 29094 28984
rect 29140 28938 29205 28984
rect 29093 28863 29205 28938
tri 29205 28863 29337 28995 sw
rect 70813 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
rect 70813 28932 71000 28990
rect 70813 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
tri 29093 28731 29225 28863 ne
rect 29225 28852 29337 28863
rect 29225 28806 29226 28852
rect 29272 28806 29337 28852
rect 29225 28731 29337 28806
tri 29225 28663 29293 28731 ne
rect 29293 28724 29337 28731
tri 29337 28724 29476 28863 sw
rect 70813 28828 71000 28886
rect 70813 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
rect 70813 28724 71000 28782
rect 29293 28720 29476 28724
rect 29293 28674 29358 28720
rect 29404 28674 29476 28720
rect 29293 28663 29476 28674
tri 29293 28480 29476 28663 ne
tri 29476 28599 29601 28724 sw
rect 70813 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
rect 70813 28620 71000 28678
rect 29476 28588 29601 28599
rect 29476 28542 29490 28588
rect 29536 28542 29601 28588
rect 29476 28480 29601 28542
tri 29601 28480 29720 28599 sw
rect 70813 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 70813 28516 71000 28574
tri 29476 28335 29621 28480 ne
rect 29621 28456 29720 28480
rect 29621 28410 29622 28456
rect 29668 28410 29720 28456
rect 29621 28335 29720 28410
tri 29720 28335 29865 28480 sw
rect 70813 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
rect 70813 28412 71000 28470
rect 70813 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
tri 29621 28203 29753 28335 ne
rect 29753 28324 29865 28335
rect 29753 28278 29754 28324
rect 29800 28278 29865 28324
rect 29753 28236 29865 28278
tri 29865 28236 29964 28335 sw
rect 70813 28308 71000 28366
rect 70813 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
rect 29753 28203 29964 28236
tri 29753 28071 29885 28203 ne
rect 29885 28192 29964 28203
rect 29885 28146 29886 28192
rect 29932 28146 29964 28192
rect 29885 28071 29964 28146
tri 29964 28071 30129 28236 sw
rect 70813 28204 71000 28262
rect 70813 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
rect 70813 28100 71000 28158
tri 29885 27939 30017 28071 ne
rect 30017 28060 30129 28071
rect 30017 28014 30018 28060
rect 30064 28014 30129 28060
rect 30017 27992 30129 28014
tri 30129 27992 30208 28071 sw
rect 70813 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 70813 27996 71000 28054
rect 30017 27939 30208 27992
tri 30017 27807 30149 27939 ne
rect 30149 27928 30208 27939
rect 30149 27882 30150 27928
rect 30196 27882 30208 27928
rect 30149 27807 30208 27882
tri 30208 27807 30393 27992 sw
rect 70813 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
rect 70813 27892 71000 27950
rect 70813 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
tri 30149 27675 30281 27807 ne
rect 30281 27796 30393 27807
rect 30281 27750 30282 27796
rect 30328 27750 30393 27796
rect 30281 27675 30393 27750
tri 30393 27675 30525 27807 sw
rect 70813 27788 71000 27846
rect 70813 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
rect 70813 27684 71000 27742
tri 30281 27543 30413 27675 ne
rect 30413 27664 30525 27675
rect 30413 27618 30414 27664
rect 30460 27618 30525 27664
rect 30413 27543 30525 27618
tri 30525 27543 30657 27675 sw
rect 70813 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 70813 27580 71000 27638
tri 30413 27411 30545 27543 ne
rect 30545 27532 30657 27543
rect 30545 27486 30546 27532
rect 30592 27486 30657 27532
rect 30545 27411 30657 27486
tri 30657 27411 30789 27543 sw
rect 70813 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
rect 70813 27476 71000 27534
rect 70813 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
tri 30545 27279 30677 27411 ne
rect 30677 27400 30789 27411
rect 30677 27354 30678 27400
rect 30724 27354 30789 27400
rect 30677 27279 30789 27354
tri 30789 27279 30921 27411 sw
rect 70813 27372 71000 27430
rect 70813 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
tri 30677 27147 30809 27279 ne
rect 30809 27268 30921 27279
rect 30809 27222 30810 27268
rect 30856 27222 30921 27268
rect 30809 27147 30921 27222
tri 30921 27147 31053 27279 sw
rect 70813 27268 71000 27326
rect 70813 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
rect 70813 27164 71000 27222
tri 30809 27015 30941 27147 ne
rect 30941 27136 31053 27147
rect 30941 27090 30942 27136
rect 30988 27090 31053 27136
rect 30941 27016 31053 27090
tri 31053 27016 31184 27147 sw
rect 70813 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
rect 70813 27060 71000 27118
rect 30941 27015 31184 27016
tri 30941 26883 31073 27015 ne
rect 31073 27004 31184 27015
rect 31073 26958 31074 27004
rect 31120 26958 31184 27004
rect 31073 26883 31184 26958
tri 31184 26883 31317 27016 sw
rect 70813 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
rect 70813 26956 71000 27014
rect 70813 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
tri 31073 26751 31205 26883 ne
rect 31205 26872 31317 26883
rect 31205 26826 31206 26872
rect 31252 26826 31317 26872
rect 31205 26772 31317 26826
tri 31317 26772 31428 26883 sw
rect 70813 26852 71000 26910
rect 70813 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
rect 31205 26751 31428 26772
tri 31205 26619 31337 26751 ne
rect 31337 26740 31428 26751
rect 31337 26694 31338 26740
rect 31384 26694 31428 26740
rect 31337 26619 31428 26694
tri 31428 26619 31581 26772 sw
rect 70813 26748 71000 26806
rect 70813 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
rect 70813 26644 71000 26702
tri 31337 26487 31469 26619 ne
rect 31469 26608 31581 26619
rect 31469 26562 31470 26608
rect 31516 26562 31581 26608
rect 31469 26528 31581 26562
tri 31581 26528 31672 26619 sw
rect 70813 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
rect 70813 26540 71000 26598
rect 31469 26487 31672 26528
tri 31469 26355 31601 26487 ne
rect 31601 26476 31672 26487
rect 31601 26430 31602 26476
rect 31648 26430 31672 26476
rect 31601 26355 31672 26430
tri 31672 26355 31845 26528 sw
rect 70813 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
rect 70813 26436 71000 26494
rect 70813 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
tri 31601 26223 31733 26355 ne
rect 31733 26344 31845 26355
rect 31733 26298 31734 26344
rect 31780 26298 31845 26344
rect 31733 26223 31845 26298
tri 31845 26223 31977 26355 sw
rect 70813 26332 71000 26390
rect 70813 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
rect 70813 26228 71000 26286
tri 31733 26091 31865 26223 ne
rect 31865 26212 31977 26223
rect 31865 26166 31866 26212
rect 31912 26166 31977 26212
rect 31865 26091 31977 26166
tri 31977 26091 32109 26223 sw
rect 70813 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
rect 70813 26124 71000 26182
tri 31865 25959 31997 26091 ne
rect 31997 26080 32109 26091
rect 31997 26034 31998 26080
rect 32044 26034 32109 26080
rect 31997 25959 32109 26034
tri 32109 25959 32241 26091 sw
rect 70813 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 70813 26020 71000 26078
rect 70813 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
tri 31997 25827 32129 25959 ne
rect 32129 25948 32241 25959
rect 32129 25902 32130 25948
rect 32176 25902 32241 25948
rect 32129 25827 32241 25902
tri 32241 25827 32373 25959 sw
rect 70813 25916 71000 25974
rect 70813 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
tri 32129 25695 32261 25827 ne
rect 32261 25816 32373 25827
rect 32261 25770 32262 25816
rect 32308 25770 32373 25816
rect 32261 25695 32373 25770
tri 32373 25695 32505 25827 sw
rect 70813 25812 71000 25870
rect 70813 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
rect 70813 25708 71000 25766
tri 32261 25563 32393 25695 ne
rect 32393 25684 32505 25695
rect 32393 25638 32394 25684
rect 32440 25638 32505 25684
rect 32393 25563 32505 25638
tri 32393 25495 32461 25563 ne
rect 32461 25552 32505 25563
tri 32505 25552 32648 25695 sw
rect 70813 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 70813 25604 71000 25662
rect 70813 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
rect 32461 25506 32526 25552
rect 32572 25506 32648 25552
rect 32461 25495 32648 25506
tri 32461 25308 32648 25495 ne
tri 32648 25431 32769 25552 sw
rect 70813 25500 71000 25558
rect 70813 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
rect 32648 25420 32769 25431
rect 32648 25374 32658 25420
rect 32704 25374 32769 25420
rect 32648 25308 32769 25374
tri 32769 25308 32892 25431 sw
rect 70813 25396 71000 25454
rect 70813 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
tri 32648 25167 32789 25308 ne
rect 32789 25288 32892 25308
rect 32789 25242 32790 25288
rect 32836 25242 32892 25288
rect 32789 25167 32892 25242
tri 32892 25167 33033 25308 sw
rect 70813 25292 71000 25350
rect 70813 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
rect 70813 25188 71000 25246
tri 32789 25035 32921 25167 ne
rect 32921 25156 33033 25167
rect 32921 25110 32922 25156
rect 32968 25110 33033 25156
rect 32921 25064 33033 25110
tri 33033 25064 33136 25167 sw
rect 70813 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
rect 70813 25084 71000 25142
rect 32921 25035 33136 25064
tri 32921 24903 33053 25035 ne
rect 33053 25024 33136 25035
rect 33053 24978 33054 25024
rect 33100 24978 33136 25024
rect 33053 24903 33136 24978
tri 33136 24903 33297 25064 sw
rect 70813 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
rect 70813 24980 71000 25038
rect 70813 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
tri 33053 24771 33185 24903 ne
rect 33185 24892 33297 24903
rect 33185 24846 33186 24892
rect 33232 24846 33297 24892
rect 33185 24820 33297 24846
tri 33297 24820 33380 24903 sw
rect 70813 24876 71000 24934
rect 70813 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
rect 33185 24771 33380 24820
tri 33185 24639 33317 24771 ne
rect 33317 24760 33380 24771
rect 33317 24714 33318 24760
rect 33364 24714 33380 24760
rect 33317 24639 33380 24714
tri 33380 24639 33561 24820 sw
rect 70813 24772 71000 24830
rect 70813 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
rect 70813 24668 71000 24726
tri 33317 24507 33449 24639 ne
rect 33449 24628 33561 24639
rect 33449 24582 33450 24628
rect 33496 24582 33561 24628
rect 33449 24507 33561 24582
tri 33561 24507 33693 24639 sw
rect 70813 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 70813 24564 71000 24622
rect 70813 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
tri 33449 24375 33581 24507 ne
rect 33581 24496 33693 24507
rect 33581 24450 33582 24496
rect 33628 24450 33693 24496
rect 33581 24375 33693 24450
tri 33693 24375 33825 24507 sw
rect 70813 24460 71000 24518
rect 70813 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
tri 33581 24243 33713 24375 ne
rect 33713 24364 33825 24375
rect 33713 24318 33714 24364
rect 33760 24318 33825 24364
rect 33713 24243 33825 24318
tri 33825 24243 33957 24375 sw
rect 70813 24356 71000 24414
rect 70813 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
rect 70813 24252 71000 24310
tri 33713 24111 33845 24243 ne
rect 33845 24232 33957 24243
rect 33845 24186 33846 24232
rect 33892 24186 33957 24232
rect 33845 24111 33957 24186
tri 33957 24111 34089 24243 sw
rect 70813 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
rect 70813 24148 71000 24206
tri 33845 23979 33977 24111 ne
rect 33977 24100 34089 24111
rect 33977 24054 33978 24100
rect 34024 24054 34089 24100
rect 33977 23979 34089 24054
tri 34089 23979 34221 24111 sw
rect 70813 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
rect 70813 24044 71000 24102
rect 70813 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
tri 33977 23847 34109 23979 ne
rect 34109 23968 34221 23979
rect 34109 23922 34110 23968
rect 34156 23922 34221 23968
rect 34109 23847 34221 23922
tri 34109 23779 34177 23847 ne
rect 34177 23844 34221 23847
tri 34221 23844 34356 23979 sw
rect 70813 23940 71000 23998
rect 70813 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
rect 34177 23836 34356 23844
rect 34177 23790 34242 23836
rect 34288 23790 34356 23836
rect 34177 23779 34356 23790
tri 34177 23600 34356 23779 ne
tri 34356 23715 34485 23844 sw
rect 70813 23836 71000 23894
rect 70813 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
rect 70813 23732 71000 23790
rect 34356 23704 34485 23715
rect 34356 23658 34374 23704
rect 34420 23658 34485 23704
rect 34356 23600 34485 23658
tri 34485 23600 34600 23715 sw
rect 70813 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 70813 23628 71000 23686
tri 34356 23451 34505 23600 ne
rect 34505 23572 34600 23600
rect 34505 23526 34506 23572
rect 34552 23526 34600 23572
rect 34505 23451 34600 23526
tri 34600 23451 34749 23600 sw
rect 70813 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
rect 70813 23524 71000 23582
rect 70813 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
tri 34505 23319 34637 23451 ne
rect 34637 23440 34749 23451
rect 34637 23394 34638 23440
rect 34684 23394 34749 23440
rect 34637 23356 34749 23394
tri 34749 23356 34844 23451 sw
rect 70813 23420 71000 23478
rect 70813 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
rect 34637 23319 34844 23356
tri 34637 23187 34769 23319 ne
rect 34769 23308 34844 23319
rect 34769 23262 34770 23308
rect 34816 23262 34844 23308
rect 34769 23187 34844 23262
tri 34844 23187 35013 23356 sw
rect 70813 23316 71000 23374
rect 70813 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
rect 70813 23212 71000 23270
tri 34769 23055 34901 23187 ne
rect 34901 23176 35013 23187
rect 34901 23130 34902 23176
rect 34948 23130 35013 23176
rect 34901 23055 35013 23130
tri 35013 23055 35145 23187 sw
rect 70813 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
rect 70813 23108 71000 23166
rect 70813 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
tri 34901 22923 35033 23055 ne
rect 35033 23044 35145 23055
rect 35033 22998 35034 23044
rect 35080 22998 35145 23044
rect 35033 22923 35145 22998
tri 35145 22923 35277 23055 sw
rect 70813 23004 71000 23062
rect 70813 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
tri 35033 22791 35165 22923 ne
rect 35165 22912 35277 22923
rect 35165 22866 35166 22912
rect 35212 22866 35277 22912
rect 35165 22791 35277 22866
tri 35277 22791 35409 22923 sw
rect 70813 22900 71000 22958
rect 70813 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
rect 70813 22796 71000 22854
tri 35165 22659 35297 22791 ne
rect 35297 22780 35409 22791
rect 35297 22734 35298 22780
rect 35344 22734 35409 22780
rect 35297 22659 35409 22734
tri 35409 22659 35541 22791 sw
rect 70813 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
rect 70813 22692 71000 22750
tri 35297 22527 35429 22659 ne
rect 35429 22648 35541 22659
rect 35429 22602 35430 22648
rect 35476 22602 35541 22648
rect 35429 22527 35541 22602
tri 35541 22527 35673 22659 sw
rect 70813 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 70813 22588 71000 22646
rect 70813 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
tri 35429 22395 35561 22527 ne
rect 35561 22516 35673 22527
rect 35561 22470 35562 22516
rect 35608 22470 35673 22516
rect 35561 22395 35673 22470
tri 35673 22395 35805 22527 sw
rect 70813 22484 71000 22542
rect 70813 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
tri 35561 22263 35693 22395 ne
rect 35693 22384 35805 22395
rect 35693 22338 35694 22384
rect 35740 22338 35805 22384
rect 35693 22263 35805 22338
tri 35805 22263 35937 22395 sw
rect 70813 22380 71000 22438
rect 70813 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
rect 70813 22276 71000 22334
tri 35693 22131 35825 22263 ne
rect 35825 22252 35937 22263
rect 35825 22206 35826 22252
rect 35872 22206 35937 22252
rect 35825 22136 35937 22206
tri 35937 22136 36064 22263 sw
rect 70813 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 70813 22172 71000 22230
rect 35825 22131 36064 22136
tri 35825 21999 35957 22131 ne
rect 35957 22120 36064 22131
rect 35957 22074 35958 22120
rect 36004 22074 36064 22120
rect 35957 21999 36064 22074
tri 36064 21999 36201 22136 sw
rect 70813 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
rect 70813 22068 71000 22126
rect 70813 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
tri 35957 21867 36089 21999 ne
rect 36089 21988 36201 21999
rect 36089 21942 36090 21988
rect 36136 21942 36201 21988
rect 36089 21892 36201 21942
tri 36201 21892 36308 21999 sw
rect 70813 21964 71000 22022
rect 70813 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
rect 36089 21867 36308 21892
tri 36089 21735 36221 21867 ne
rect 36221 21856 36308 21867
rect 36221 21810 36222 21856
rect 36268 21810 36308 21856
rect 36221 21735 36308 21810
tri 36308 21735 36465 21892 sw
rect 70813 21860 71000 21918
rect 70813 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
rect 70813 21756 71000 21814
tri 36221 21603 36353 21735 ne
rect 36353 21724 36465 21735
rect 36353 21678 36354 21724
rect 36400 21678 36465 21724
rect 36353 21648 36465 21678
tri 36465 21648 36552 21735 sw
rect 70813 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
rect 70813 21652 71000 21710
rect 36353 21603 36552 21648
tri 36353 21471 36485 21603 ne
rect 36485 21592 36552 21603
rect 36485 21546 36486 21592
rect 36532 21546 36552 21592
rect 36485 21471 36552 21546
tri 36552 21471 36729 21648 sw
rect 70813 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
rect 70813 21548 71000 21606
rect 70813 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
tri 36485 21339 36617 21471 ne
rect 36617 21460 36729 21471
rect 36617 21414 36618 21460
rect 36664 21414 36729 21460
rect 36617 21339 36729 21414
tri 36729 21339 36861 21471 sw
rect 70813 21444 71000 21502
rect 70813 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
rect 70813 21340 71000 21398
tri 36617 21207 36749 21339 ne
rect 36749 21328 36861 21339
rect 36749 21282 36750 21328
rect 36796 21282 36861 21328
rect 36749 21207 36861 21282
tri 36861 21207 36993 21339 sw
rect 70813 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 70813 21236 71000 21294
tri 36749 21075 36881 21207 ne
rect 36881 21196 36993 21207
rect 36881 21150 36882 21196
rect 36928 21150 36993 21196
rect 36881 21075 36993 21150
tri 36993 21075 37125 21207 sw
rect 70813 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 70813 21132 71000 21190
rect 70813 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
tri 36881 20943 37013 21075 ne
rect 37013 21064 37125 21075
rect 37013 21018 37014 21064
rect 37060 21018 37125 21064
rect 37013 20943 37125 21018
tri 37125 20943 37257 21075 sw
rect 70813 21028 71000 21086
rect 70813 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
tri 37013 20811 37145 20943 ne
rect 37145 20932 37257 20943
rect 37145 20886 37146 20932
rect 37192 20886 37257 20932
rect 37145 20811 37257 20886
tri 37257 20811 37389 20943 sw
rect 70813 20924 71000 20982
rect 70813 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
rect 70813 20820 71000 20878
tri 37145 20679 37277 20811 ne
rect 37277 20800 37389 20811
rect 37277 20754 37278 20800
rect 37324 20754 37389 20800
rect 37277 20679 37389 20754
tri 37277 20611 37345 20679 ne
rect 37345 20672 37389 20679
tri 37389 20672 37528 20811 sw
rect 70813 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
rect 70813 20716 71000 20774
rect 37345 20668 37528 20672
rect 37345 20622 37410 20668
rect 37456 20622 37528 20668
rect 37345 20611 37528 20622
tri 37345 20428 37528 20611 ne
tri 37528 20547 37653 20672 sw
rect 70813 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
rect 70813 20612 71000 20670
rect 70813 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
rect 37528 20536 37653 20547
rect 37528 20490 37542 20536
rect 37588 20490 37653 20536
rect 37528 20428 37653 20490
tri 37653 20428 37772 20547 sw
rect 70813 20508 71000 20566
rect 70813 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
tri 37528 20283 37673 20428 ne
rect 37673 20404 37772 20428
rect 37673 20358 37674 20404
rect 37720 20358 37772 20404
rect 37673 20283 37772 20358
tri 37772 20283 37917 20428 sw
rect 70813 20404 71000 20462
rect 70813 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
rect 70813 20300 71000 20358
tri 37673 20151 37805 20283 ne
rect 37805 20272 37917 20283
rect 37805 20226 37806 20272
rect 37852 20226 37917 20272
rect 37805 20184 37917 20226
tri 37917 20184 38016 20283 sw
rect 70813 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 70813 20196 71000 20254
rect 37805 20151 38016 20184
tri 37805 20019 37937 20151 ne
rect 37937 20140 38016 20151
rect 37937 20094 37938 20140
rect 37984 20094 38016 20140
rect 37937 20019 38016 20094
tri 38016 20019 38181 20184 sw
rect 70813 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
rect 70813 20092 71000 20150
rect 70813 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
tri 37937 19887 38069 20019 ne
rect 38069 20008 38181 20019
rect 38069 19962 38070 20008
rect 38116 19962 38181 20008
rect 38069 19940 38181 19962
tri 38181 19940 38260 20019 sw
rect 70813 19988 71000 20046
rect 70813 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
rect 38069 19887 38260 19940
tri 38069 19755 38201 19887 ne
rect 38201 19876 38260 19887
rect 38201 19830 38202 19876
rect 38248 19830 38260 19876
rect 38201 19755 38260 19830
tri 38260 19755 38445 19940 sw
rect 70813 19884 71000 19942
rect 70813 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
rect 70813 19780 71000 19838
tri 38201 19623 38333 19755 ne
rect 38333 19744 38445 19755
rect 38333 19698 38334 19744
rect 38380 19698 38445 19744
rect 38333 19623 38445 19698
tri 38445 19623 38577 19755 sw
rect 70813 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
rect 70813 19676 71000 19734
rect 70813 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
tri 38333 19491 38465 19623 ne
rect 38465 19612 38577 19623
rect 38465 19566 38466 19612
rect 38512 19566 38577 19612
rect 38465 19491 38577 19566
tri 38577 19491 38709 19623 sw
rect 70813 19572 71000 19630
rect 70813 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
tri 38465 19359 38597 19491 ne
rect 38597 19480 38709 19491
rect 38597 19434 38598 19480
rect 38644 19434 38709 19480
rect 38597 19359 38709 19434
tri 38709 19359 38841 19491 sw
rect 70813 19468 71000 19526
rect 70813 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
rect 70813 19364 71000 19422
tri 38597 19227 38729 19359 ne
rect 38729 19348 38841 19359
rect 38729 19302 38730 19348
rect 38776 19302 38841 19348
rect 38729 19227 38841 19302
tri 38841 19227 38973 19359 sw
rect 70813 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
rect 70813 19260 71000 19318
tri 38729 19095 38861 19227 ne
rect 38861 19216 38973 19227
rect 38861 19170 38862 19216
rect 38908 19170 38973 19216
rect 38861 19095 38973 19170
tri 38973 19095 39105 19227 sw
rect 70813 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 70813 19156 71000 19214
rect 70813 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
tri 38861 18963 38993 19095 ne
rect 38993 19084 39105 19095
rect 38993 19038 38994 19084
rect 39040 19038 39105 19084
rect 38993 18964 39105 19038
tri 39105 18964 39236 19095 sw
rect 70813 19052 71000 19110
rect 70813 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
rect 38993 18963 39236 18964
tri 38993 18831 39125 18963 ne
rect 39125 18952 39236 18963
rect 39125 18906 39126 18952
rect 39172 18906 39236 18952
rect 39125 18831 39236 18906
tri 39236 18831 39369 18964 sw
rect 70813 18948 71000 19006
rect 70813 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
rect 70813 18844 71000 18902
tri 39125 18699 39257 18831 ne
rect 39257 18820 39369 18831
rect 39257 18774 39258 18820
rect 39304 18774 39369 18820
rect 39257 18720 39369 18774
tri 39369 18720 39480 18831 sw
rect 70813 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 70813 18740 71000 18798
rect 39257 18699 39480 18720
tri 39257 18567 39389 18699 ne
rect 39389 18688 39480 18699
rect 39389 18642 39390 18688
rect 39436 18642 39480 18688
rect 39389 18567 39480 18642
tri 39480 18567 39633 18720 sw
rect 70813 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
rect 70813 18636 71000 18694
rect 70813 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
tri 39389 18435 39521 18567 ne
rect 39521 18556 39633 18567
rect 39521 18510 39522 18556
rect 39568 18510 39633 18556
rect 39521 18476 39633 18510
tri 39633 18476 39724 18567 sw
rect 70813 18532 71000 18590
rect 70813 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
rect 39521 18435 39724 18476
tri 39521 18303 39653 18435 ne
rect 39653 18424 39724 18435
rect 39653 18378 39654 18424
rect 39700 18378 39724 18424
rect 39653 18303 39724 18378
tri 39724 18303 39897 18476 sw
rect 70813 18428 71000 18486
rect 70813 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
rect 70813 18324 71000 18382
tri 39653 18171 39785 18303 ne
rect 39785 18292 39897 18303
rect 39785 18246 39786 18292
rect 39832 18246 39897 18292
rect 39785 18171 39897 18246
tri 39897 18171 40029 18303 sw
rect 70813 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
rect 70813 18220 71000 18278
rect 70813 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
tri 39785 18039 39917 18171 ne
rect 39917 18160 40029 18171
rect 39917 18114 39918 18160
rect 39964 18114 40029 18160
rect 39917 18039 40029 18114
tri 40029 18039 40161 18171 sw
rect 70813 18116 71000 18174
rect 70813 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
tri 39917 17907 40049 18039 ne
rect 40049 18028 40161 18039
rect 40049 17982 40050 18028
rect 40096 17982 40161 18028
rect 40049 17907 40161 17982
tri 40161 17907 40293 18039 sw
rect 70813 18012 71000 18070
rect 70813 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
rect 70813 17908 71000 17966
tri 40049 17775 40181 17907 ne
rect 40181 17896 40293 17907
rect 40181 17850 40182 17896
rect 40228 17850 40293 17896
rect 40181 17775 40293 17850
tri 40293 17775 40425 17907 sw
rect 70813 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
rect 70813 17804 71000 17862
tri 40181 17643 40313 17775 ne
rect 40313 17764 40425 17775
rect 40313 17718 40314 17764
rect 40360 17718 40425 17764
rect 40313 17643 40425 17718
tri 40425 17643 40557 17775 sw
rect 70813 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 70813 17700 71000 17758
rect 70813 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
tri 40313 17511 40445 17643 ne
rect 40445 17632 40557 17643
rect 40445 17586 40446 17632
rect 40492 17586 40557 17632
rect 40445 17511 40557 17586
tri 40445 17443 40513 17511 ne
rect 40513 17500 40557 17511
tri 40557 17500 40700 17643 sw
rect 70813 17596 71000 17654
rect 70813 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
rect 40513 17454 40578 17500
rect 40624 17454 40700 17500
rect 40513 17443 40700 17454
tri 40513 17256 40700 17443 ne
tri 40700 17379 40821 17500 sw
rect 70813 17492 71000 17550
rect 70813 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
rect 70813 17388 71000 17446
rect 40700 17368 40821 17379
rect 40700 17322 40710 17368
rect 40756 17322 40821 17368
rect 40700 17256 40821 17322
tri 40821 17256 40944 17379 sw
rect 70813 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 70813 17284 71000 17342
tri 40700 17115 40841 17256 ne
rect 40841 17236 40944 17256
rect 40841 17190 40842 17236
rect 40888 17190 40944 17236
rect 40841 17115 40944 17190
tri 40944 17115 41085 17256 sw
rect 70813 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
rect 70813 17180 71000 17238
rect 70813 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
tri 40841 16983 40973 17115 ne
rect 40973 17104 41085 17115
rect 40973 17058 40974 17104
rect 41020 17058 41085 17104
rect 40973 17012 41085 17058
tri 41085 17012 41188 17115 sw
rect 70813 17076 71000 17134
rect 70813 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
rect 40973 16983 41188 17012
tri 40973 16851 41105 16983 ne
rect 41105 16972 41188 16983
rect 41105 16926 41106 16972
rect 41152 16926 41188 16972
rect 41105 16851 41188 16926
tri 41188 16851 41349 17012 sw
rect 70813 16972 71000 17030
rect 70813 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
rect 70813 16868 71000 16926
tri 41105 16719 41237 16851 ne
rect 41237 16840 41349 16851
rect 41237 16794 41238 16840
rect 41284 16794 41349 16840
rect 41237 16768 41349 16794
tri 41349 16768 41432 16851 sw
rect 70813 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 41237 16719 41432 16768
tri 41237 16587 41369 16719 ne
rect 41369 16708 41432 16719
rect 41369 16662 41370 16708
rect 41416 16662 41432 16708
rect 41369 16587 41432 16662
tri 41432 16587 41613 16768 sw
rect 70813 16764 71000 16822
rect 70813 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
rect 70813 16660 71000 16718
rect 70813 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
tri 41369 16455 41501 16587 ne
rect 41501 16576 41613 16587
rect 41501 16530 41502 16576
rect 41548 16530 41613 16576
rect 41501 16455 41613 16530
tri 41613 16455 41745 16587 sw
rect 70813 16556 71000 16614
rect 70813 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
tri 41501 16323 41633 16455 ne
rect 41633 16444 41745 16455
rect 41633 16398 41634 16444
rect 41680 16398 41745 16444
rect 41633 16323 41745 16398
tri 41745 16323 41877 16455 sw
rect 70813 16452 71000 16510
rect 70813 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
rect 70813 16348 71000 16406
tri 41633 16191 41765 16323 ne
rect 41765 16312 41877 16323
rect 41765 16266 41766 16312
rect 41812 16266 41877 16312
rect 41765 16191 41877 16266
tri 41877 16191 42009 16323 sw
rect 70813 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 70813 16244 71000 16302
rect 70813 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
tri 41765 16059 41897 16191 ne
rect 41897 16180 42009 16191
rect 41897 16134 41898 16180
rect 41944 16134 42009 16180
rect 41897 16059 42009 16134
tri 42009 16059 42141 16191 sw
rect 70813 16140 71000 16198
rect 70813 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
tri 41897 15927 42029 16059 ne
rect 42029 16048 42141 16059
rect 42029 16002 42030 16048
rect 42076 16002 42141 16048
rect 42029 15927 42141 16002
tri 42141 15927 42273 16059 sw
rect 70813 16036 71000 16094
rect 70813 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
rect 70813 15932 71000 15990
tri 42029 15795 42161 15927 ne
rect 42161 15916 42273 15927
rect 42161 15870 42162 15916
rect 42208 15870 42273 15916
rect 42161 15795 42273 15870
tri 42161 15727 42229 15795 ne
rect 42229 15792 42273 15795
tri 42273 15792 42408 15927 sw
rect 70813 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
rect 70813 15828 71000 15886
rect 42229 15784 42408 15792
rect 42229 15738 42294 15784
rect 42340 15738 42408 15784
rect 42229 15727 42408 15738
tri 42229 15548 42408 15727 ne
tri 42408 15663 42537 15792 sw
rect 70813 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 70813 15724 71000 15782
rect 70813 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
rect 42408 15652 42537 15663
rect 42408 15606 42426 15652
rect 42472 15606 42537 15652
rect 42408 15548 42537 15606
tri 42537 15548 42652 15663 sw
rect 70813 15620 71000 15678
rect 70813 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
tri 42408 15399 42557 15548 ne
rect 42557 15520 42652 15548
rect 42557 15474 42558 15520
rect 42604 15474 42652 15520
rect 42557 15399 42652 15474
tri 42652 15399 42801 15548 sw
rect 70813 15516 71000 15574
rect 70813 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
rect 70813 15412 71000 15470
tri 42557 15267 42689 15399 ne
rect 42689 15388 42801 15399
rect 42689 15342 42690 15388
rect 42736 15342 42801 15388
rect 42689 15304 42801 15342
tri 42801 15304 42896 15399 sw
rect 70813 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 70813 15308 71000 15366
rect 42689 15267 42896 15304
tri 42689 15135 42821 15267 ne
rect 42821 15256 42896 15267
rect 42821 15210 42822 15256
rect 42868 15210 42896 15256
rect 42821 15135 42896 15210
tri 42896 15135 43065 15304 sw
rect 70813 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
rect 70813 15204 71000 15262
rect 70813 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
tri 42821 15003 42953 15135 ne
rect 42953 15124 43065 15135
rect 42953 15078 42954 15124
rect 43000 15078 43065 15124
rect 42953 15003 43065 15078
tri 43065 15003 43197 15135 sw
rect 70813 15100 71000 15158
rect 70813 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
tri 42953 14871 43085 15003 ne
rect 43085 14992 43197 15003
rect 43085 14946 43086 14992
rect 43132 14946 43197 14992
rect 43085 14871 43197 14946
tri 43197 14871 43329 15003 sw
rect 70813 14996 71000 15054
rect 70813 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
rect 70813 14892 71000 14950
tri 43085 14739 43217 14871 ne
rect 43217 14860 43329 14871
rect 43217 14814 43218 14860
rect 43264 14814 43329 14860
rect 43217 14739 43329 14814
tri 43329 14739 43461 14871 sw
rect 70813 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
rect 70813 14788 71000 14846
rect 70813 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
tri 43217 14607 43349 14739 ne
rect 43349 14728 43461 14739
rect 43349 14682 43350 14728
rect 43396 14682 43461 14728
rect 43349 14607 43461 14682
tri 43461 14607 43593 14739 sw
rect 70813 14684 71000 14742
rect 70813 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
tri 43349 14475 43481 14607 ne
rect 43481 14596 43593 14607
rect 43481 14550 43482 14596
rect 43528 14550 43593 14596
rect 43481 14475 43593 14550
tri 43593 14475 43725 14607 sw
rect 70813 14580 71000 14638
rect 70813 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
rect 70813 14476 71000 14534
tri 43481 14343 43613 14475 ne
rect 43613 14464 43725 14475
rect 43613 14418 43614 14464
rect 43660 14418 43725 14464
rect 43613 14343 43725 14418
tri 43725 14343 43857 14475 sw
rect 70813 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
rect 70813 14372 71000 14430
tri 43613 14211 43745 14343 ne
rect 43745 14332 43857 14343
rect 43745 14286 43746 14332
rect 43792 14286 43857 14332
rect 43745 14211 43857 14286
tri 43857 14211 43989 14343 sw
rect 70813 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 70813 14268 71000 14326
rect 70813 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
tri 43745 14079 43877 14211 ne
rect 43877 14200 43989 14211
rect 43877 14154 43878 14200
rect 43924 14154 43989 14200
rect 43877 14084 43989 14154
tri 43989 14084 44116 14211 sw
rect 70813 14164 71000 14222
rect 70813 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
rect 43877 14079 44116 14084
tri 43877 13947 44009 14079 ne
rect 44009 14068 44116 14079
rect 44009 14022 44010 14068
rect 44056 14022 44116 14068
rect 44009 13947 44116 14022
tri 44116 13947 44253 14084 sw
rect 70813 14060 71000 14118
rect 70813 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
rect 70813 13956 71000 14014
tri 44009 13815 44141 13947 ne
rect 44141 13936 44253 13947
rect 44141 13890 44142 13936
rect 44188 13890 44253 13936
rect 44141 13840 44253 13890
tri 44253 13840 44360 13947 sw
rect 70813 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
rect 70813 13852 71000 13910
rect 44141 13815 44360 13840
tri 44141 13683 44273 13815 ne
rect 44273 13804 44360 13815
rect 44273 13758 44274 13804
rect 44320 13758 44360 13804
rect 44273 13683 44360 13758
tri 44360 13683 44517 13840 sw
rect 70813 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
rect 70813 13748 71000 13806
rect 70813 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
tri 44273 13551 44405 13683 ne
rect 44405 13672 44517 13683
rect 44405 13626 44406 13672
rect 44452 13626 44517 13672
rect 44405 13596 44517 13626
tri 44517 13596 44604 13683 sw
rect 70813 13644 71000 13702
rect 70813 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
rect 44405 13551 44604 13596
tri 44405 13419 44537 13551 ne
rect 44537 13540 44604 13551
rect 44537 13494 44538 13540
rect 44584 13494 44604 13540
rect 44537 13419 44604 13494
tri 44604 13419 44781 13596 sw
rect 70813 13540 71000 13598
rect 70813 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
rect 70813 13436 71000 13494
tri 44537 13351 44605 13419 ne
rect 44605 13408 44781 13419
rect 44605 13362 44670 13408
rect 44716 13362 44781 13408
rect 44605 13352 44781 13362
tri 44781 13352 44848 13419 sw
rect 70813 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 44605 13351 44848 13352
tri 44605 13108 44848 13351 ne
tri 44848 13280 44920 13352 sw
rect 70813 13280 71000 13390
rect 44848 13269 71000 13280
rect 44848 13256 45088 13269
rect 44848 13210 44850 13256
rect 44896 13223 45088 13256
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 44896 13210 71000 13223
rect 44848 13165 71000 13210
rect 44848 13119 45088 13165
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
rect 44848 13108 71000 13119
<< metal2 >>
rect 70584 68116 70702 68200
rect 70584 66916 70613 68116
rect 70669 66916 70702 68116
rect 70584 60120 70702 66916
rect 70584 58920 70613 60120
rect 70669 58920 70702 60120
rect 70584 56910 70702 58920
rect 70584 55710 70613 56910
rect 70669 55710 70702 56910
rect 70584 55302 70702 55710
rect 70584 54102 70613 55302
rect 70669 54102 70702 55302
rect 70584 53722 70702 54102
rect 70584 52522 70613 53722
rect 70669 52522 70702 53722
rect 70584 45739 70702 52522
rect 70584 42875 70613 45739
rect 70669 42875 70702 45739
rect 70584 42497 70702 42875
rect 70584 41297 70613 42497
rect 70669 41297 70702 42497
rect 70584 39332 70702 41297
rect 70584 36468 70613 39332
rect 70669 36468 70702 39332
rect 70584 36132 70702 36468
rect 70584 33268 70613 36132
rect 70669 33268 70702 36132
rect 70584 32920 70702 33268
rect 70584 30056 70613 32920
rect 70669 30056 70702 32920
rect 70584 29752 70702 30056
rect 70584 26888 70613 29752
rect 70669 26888 70702 29752
rect 70584 24906 70702 26888
rect 70584 23706 70613 24906
rect 70669 23706 70702 24906
rect 70584 23599 70702 23706
<< via2 >>
rect 70613 66916 70669 68116
rect 70613 58920 70669 60120
rect 70613 55710 70669 56910
rect 70613 54102 70669 55302
rect 70613 52522 70669 53722
rect 70613 42875 70669 45739
rect 70613 41297 70669 42497
rect 70613 36468 70669 39332
rect 70613 33268 70669 36132
rect 70613 30056 70669 32920
rect 70613 26888 70669 29752
rect 70613 23706 70669 24906
<< metal3 >>
rect 14000 47020 17000 71000
rect 17200 48366 20200 71000
rect 20400 49677 23400 71000
rect 23600 50451 25000 71000
rect 25200 51120 26600 71000
rect 26800 52360 29800 71000
rect 30000 53704 33000 71000
rect 33200 55027 36200 71000
rect 36400 56372 39400 71000
rect 39600 57138 41000 71000
rect 41200 57810 42600 71000
rect 42800 59039 45800 71000
rect 46000 60425 49000 71000
rect 49200 61175 50600 71000
rect 50800 61839 52200 71000
rect 52400 62507 53800 71000
rect 54000 63320 55400 71000
rect 55600 63836 57000 71000
rect 57200 64540 58600 71000
rect 58800 65166 60200 71000
rect 60400 65831 61800 71000
rect 62000 66494 63400 71000
rect 63600 67166 65000 71000
rect 65200 67829 66600 71000
rect 66800 68493 68200 71000
rect 68400 69678 69678 71000
rect 68400 68769 71000 69678
tri 68200 68493 68400 68693 sw
tri 68400 68493 68676 68769 ne
rect 68676 68493 71000 68769
rect 66800 68400 68400 68493
tri 68400 68400 68493 68493 sw
tri 68676 68400 68769 68493 ne
rect 68769 68400 71000 68493
rect 66800 68200 68493 68400
tri 68493 68200 68693 68400 sw
rect 66800 68116 71000 68200
rect 66800 68113 70613 68116
tri 66800 68029 66884 68113 ne
rect 66884 68029 70613 68113
tri 66600 67829 66800 68029 sw
tri 66884 67829 67084 68029 ne
rect 67084 67829 70613 68029
rect 65200 67545 66800 67829
tri 66800 67545 67084 67829 sw
tri 67084 67545 67368 67829 ne
rect 67368 67545 70613 67829
rect 65200 67449 67084 67545
tri 65200 67366 65283 67449 ne
rect 65283 67368 67084 67449
tri 67084 67368 67261 67545 sw
tri 67368 67368 67545 67545 ne
rect 67545 67368 70613 67545
rect 65283 67366 67261 67368
tri 65000 67166 65200 67366 sw
tri 65283 67166 65483 67366 ne
rect 65483 67166 67261 67366
rect 63600 66883 65200 67166
tri 65200 66883 65483 67166 sw
tri 65483 66883 65766 67166 ne
rect 65766 67084 67261 67166
tri 67261 67084 67545 67368 sw
tri 67545 67084 67829 67368 ne
rect 67829 67084 70613 67368
rect 65766 66883 67545 67084
rect 63600 66786 65483 66883
tri 63600 66694 63692 66786 ne
rect 63692 66694 65483 66786
tri 63400 66494 63600 66694 sw
tri 63692 66494 63892 66694 ne
rect 63892 66600 65483 66694
tri 65483 66600 65766 66883 sw
tri 65766 66600 66049 66883 ne
rect 66049 66800 67545 66883
tri 67545 66800 67829 67084 sw
tri 67829 66800 68113 67084 ne
rect 68113 66916 70613 67084
rect 70669 66916 71000 68116
rect 68113 66800 71000 66916
rect 66049 66600 67829 66800
tri 67829 66600 68029 66800 sw
rect 63892 66494 65766 66600
rect 62000 66202 63600 66494
tri 63600 66202 63892 66494 sw
tri 63892 66202 64184 66494 ne
rect 64184 66332 65766 66494
tri 65766 66332 66034 66600 sw
tri 66049 66332 66317 66600 ne
rect 66317 66332 71000 66600
rect 64184 66202 66034 66332
rect 62000 66114 63892 66202
tri 62000 66031 62083 66114 ne
rect 62083 66031 63892 66114
tri 61800 65831 62000 66031 sw
tri 62083 65831 62283 66031 ne
rect 62283 65964 63892 66031
tri 63892 65964 64130 66202 sw
tri 64184 65964 64422 66202 ne
rect 64422 66049 66034 66202
tri 66034 66049 66317 66332 sw
tri 66317 66049 66600 66332 ne
rect 66600 66049 71000 66332
rect 64422 65964 66317 66049
rect 62283 65831 64130 65964
rect 60400 65663 62000 65831
tri 62000 65663 62168 65831 sw
tri 62283 65663 62451 65831 ne
rect 62451 65672 64130 65831
tri 64130 65672 64422 65964 sw
tri 64422 65672 64714 65964 ne
rect 64714 65766 66317 65964
tri 66317 65766 66600 66049 sw
tri 66600 65766 66883 66049 ne
rect 66883 65766 71000 66049
rect 64714 65672 66600 65766
rect 62451 65663 64422 65672
rect 60400 65451 62168 65663
tri 60400 65366 60485 65451 ne
rect 60485 65380 62168 65451
tri 62168 65380 62451 65663 sw
tri 62451 65380 62734 65663 ne
rect 62734 65380 64422 65663
tri 64422 65380 64714 65672 sw
tri 64714 65380 65006 65672 ne
rect 65006 65483 66600 65672
tri 66600 65483 66883 65766 sw
tri 66883 65483 67166 65766 ne
rect 67166 65483 71000 65766
rect 65006 65380 66883 65483
rect 60485 65366 62451 65380
tri 60200 65166 60400 65366 sw
tri 60485 65166 60685 65366 ne
rect 60685 65166 62451 65366
rect 58800 64881 60400 65166
tri 60400 64881 60685 65166 sw
tri 60685 64881 60970 65166 ne
rect 60970 65097 62451 65166
tri 62451 65097 62734 65380 sw
tri 62734 65097 63017 65380 ne
rect 63017 65292 64714 65380
tri 64714 65292 64802 65380 sw
tri 65006 65292 65094 65380 ne
rect 65094 65292 66883 65380
rect 63017 65097 64802 65292
rect 60970 64997 62734 65097
tri 62734 64997 62834 65097 sw
tri 63017 64997 63117 65097 ne
rect 63117 65000 64802 65097
tri 64802 65000 65094 65292 sw
tri 65094 65000 65386 65292 ne
rect 65386 65200 66883 65292
tri 66883 65200 67166 65483 sw
tri 67166 65200 67449 65483 ne
rect 67449 65200 71000 65483
rect 65386 65000 67166 65200
tri 67166 65000 67366 65200 sw
rect 63117 64997 65094 65000
rect 60970 64881 62834 64997
rect 58800 64786 60685 64881
tri 58800 64699 58887 64786 ne
rect 58887 64730 60685 64786
tri 60685 64730 60836 64881 sw
tri 60970 64730 61121 64881 ne
rect 61121 64730 62834 64881
rect 58887 64699 60836 64730
tri 58600 64540 58759 64699 sw
tri 58887 64540 59046 64699 ne
rect 59046 64540 60836 64699
rect 57200 64499 58759 64540
tri 58759 64499 58800 64540 sw
tri 59046 64499 59087 64540 ne
rect 59087 64499 60836 64540
rect 57200 64447 58800 64499
tri 58800 64447 58852 64499 sw
tri 59087 64447 59139 64499 ne
rect 59139 64447 60836 64499
rect 57200 64160 58852 64447
tri 58852 64160 59139 64447 sw
tri 59139 64160 59426 64447 ne
rect 59426 64445 60836 64447
tri 60836 64445 61121 64730 sw
tri 61121 64445 61406 64730 ne
rect 61406 64714 62834 64730
tri 62834 64714 63117 64997 sw
tri 63117 64714 63400 64997 ne
rect 63400 64714 65094 64997
rect 61406 64445 63117 64714
rect 59426 64160 61121 64445
tri 61121 64160 61406 64445 sw
tri 61406 64160 61691 64445 ne
rect 61691 64431 63117 64445
tri 63117 64431 63400 64714 sw
tri 63400 64431 63683 64714 ne
rect 63683 64708 65094 64714
tri 65094 64708 65386 65000 sw
tri 65386 64708 65678 65000 ne
rect 65678 64708 71000 65000
rect 63683 64431 65386 64708
rect 61691 64160 63400 64431
rect 57200 64119 59139 64160
tri 57200 64036 57283 64119 ne
rect 57283 64036 59139 64119
tri 57000 63836 57200 64036 sw
tri 57283 63836 57483 64036 ne
rect 57483 63873 59139 64036
tri 59139 63873 59426 64160 sw
tri 59426 63873 59713 64160 ne
rect 59713 64065 61406 64160
tri 61406 64065 61501 64160 sw
tri 61691 64065 61786 64160 ne
rect 61786 64148 63400 64160
tri 63400 64148 63683 64431 sw
tri 63683 64148 63966 64431 ne
rect 63966 64416 65386 64431
tri 65386 64416 65678 64708 sw
tri 65678 64416 65970 64708 ne
rect 65970 64416 71000 64708
rect 63966 64184 65678 64416
tri 65678 64184 65910 64416 sw
tri 65970 64184 66202 64416 ne
rect 66202 64184 71000 64416
rect 63966 64148 65910 64184
rect 61786 64065 63683 64148
rect 59713 63873 61501 64065
rect 57483 63836 59426 63873
rect 55600 63553 57200 63836
tri 57200 63553 57483 63836 sw
tri 57483 63553 57766 63836 ne
rect 57766 63673 59426 63836
tri 59426 63673 59626 63873 sw
tri 59713 63673 59913 63873 ne
rect 59913 63780 61501 63873
tri 61501 63780 61786 64065 sw
tri 61786 63780 62071 64065 ne
rect 62071 63966 63683 64065
tri 63683 63966 63865 64148 sw
tri 63966 63966 64148 64148 ne
rect 64148 63966 65910 64148
rect 62071 63780 63865 63966
rect 59913 63673 61786 63780
rect 57766 63553 59626 63673
rect 55600 63506 57483 63553
tri 57483 63506 57530 63553 sw
tri 57766 63506 57813 63553 ne
rect 57813 63506 59626 63553
rect 55600 63456 57530 63506
tri 55600 63373 55683 63456 ne
rect 55683 63373 57530 63456
tri 55400 63320 55453 63373 sw
tri 55683 63320 55736 63373 ne
rect 55736 63320 57530 63373
rect 54000 63173 55453 63320
tri 55453 63173 55600 63320 sw
tri 55736 63173 55883 63320 ne
rect 55883 63223 57530 63320
tri 57530 63223 57813 63506 sw
tri 57813 63223 58096 63506 ne
rect 58096 63386 59626 63506
tri 59626 63386 59913 63673 sw
tri 59913 63386 60200 63673 ne
rect 60200 63495 61786 63673
tri 61786 63495 62071 63780 sw
tri 62071 63495 62356 63780 ne
rect 62356 63683 63865 63780
tri 63865 63683 64148 63966 sw
tri 64148 63683 64431 63966 ne
rect 64431 63892 65910 63966
tri 65910 63892 66202 64184 sw
tri 66202 63892 66494 64184 ne
rect 66494 63892 71000 64184
rect 64431 63683 66202 63892
rect 62356 63495 64148 63683
rect 60200 63386 62071 63495
rect 58096 63223 59913 63386
rect 55883 63173 57813 63223
rect 54000 62940 55600 63173
tri 55600 62940 55833 63173 sw
tri 55883 62940 56116 63173 ne
rect 56116 62940 57813 63173
tri 57813 62940 58096 63223 sw
tri 58096 62940 58379 63223 ne
rect 58379 63099 59913 63223
tri 59913 63099 60200 63386 sw
tri 60200 63099 60487 63386 ne
rect 60487 63210 62071 63386
tri 62071 63210 62356 63495 sw
tri 62356 63210 62641 63495 ne
rect 62641 63400 64148 63495
tri 64148 63400 64431 63683 sw
tri 64431 63400 64714 63683 ne
rect 64714 63600 66202 63683
tri 66202 63600 66494 63892 sw
tri 66494 63600 66786 63892 ne
rect 66786 63600 71000 63892
rect 64714 63400 66494 63600
tri 66494 63400 66694 63600 sw
rect 62641 63210 64431 63400
rect 60487 63099 62356 63210
rect 58379 62940 60200 63099
rect 54000 62793 55833 62940
tri 54000 62707 54086 62793 ne
rect 54086 62707 55833 62793
tri 53800 62507 54000 62707 sw
tri 54086 62507 54286 62707 ne
rect 54286 62657 55833 62707
tri 55833 62657 56116 62940 sw
tri 56116 62657 56399 62940 ne
rect 56399 62843 58096 62940
tri 58096 62843 58193 62940 sw
tri 58379 62843 58476 62940 ne
rect 58476 62843 60200 62940
rect 56399 62657 58193 62843
rect 54286 62622 56116 62657
tri 56116 62622 56151 62657 sw
tri 56399 62622 56434 62657 ne
rect 56434 62622 58193 62657
rect 54286 62507 56151 62622
rect 52400 62221 54000 62507
tri 54000 62221 54286 62507 sw
tri 54286 62221 54572 62507 ne
rect 54572 62339 56151 62507
tri 56151 62339 56434 62622 sw
tri 56434 62339 56717 62622 ne
rect 56717 62560 58193 62622
tri 58193 62560 58476 62843 sw
tri 58476 62560 58759 62843 ne
rect 58759 62812 60200 62843
tri 60200 62812 60487 63099 sw
tri 60487 62812 60774 63099 ne
rect 60774 62925 62356 63099
tri 62356 62925 62641 63210 sw
tri 62641 62925 62926 63210 ne
rect 62926 63117 64431 63210
tri 64431 63117 64714 63400 sw
tri 64714 63117 64997 63400 ne
rect 64997 63117 71000 63400
rect 62926 62925 64714 63117
rect 60774 62812 62641 62925
rect 58759 62754 60487 62812
tri 60487 62754 60545 62812 sw
tri 60774 62754 60832 62812 ne
rect 60832 62754 62641 62812
rect 58759 62560 60545 62754
rect 56717 62339 58476 62560
rect 54572 62221 56434 62339
rect 52400 62127 54286 62221
tri 52400 62039 52488 62127 ne
rect 52488 62039 54286 62127
tri 52200 61839 52400 62039 sw
tri 52488 61839 52688 62039 ne
rect 52688 62006 54286 62039
tri 54286 62006 54501 62221 sw
tri 54572 62006 54787 62221 ne
rect 54787 62056 56434 62221
tri 56434 62056 56717 62339 sw
tri 56717 62056 57000 62339 ne
rect 57000 62277 58476 62339
tri 58476 62277 58759 62560 sw
tri 58759 62277 59042 62560 ne
rect 59042 62467 60545 62560
tri 60545 62467 60832 62754 sw
tri 60832 62467 61119 62754 ne
rect 61119 62750 62641 62754
tri 62641 62750 62816 62925 sw
tri 62926 62750 63101 62925 ne
rect 63101 62834 64714 62925
tri 64714 62834 64997 63117 sw
tri 64997 62834 65280 63117 ne
rect 65280 62834 71000 63117
rect 63101 62750 64997 62834
rect 61119 62467 62816 62750
rect 59042 62277 60832 62467
rect 57000 62056 58759 62277
rect 54787 62006 56717 62056
rect 52688 61839 54501 62006
rect 50800 61720 52400 61839
tri 52400 61720 52519 61839 sw
tri 52688 61720 52807 61839 ne
rect 52807 61720 54501 61839
tri 54501 61720 54787 62006 sw
tri 54787 61720 55073 62006 ne
rect 55073 61773 56717 62006
tri 56717 61773 57000 62056 sw
tri 57000 61773 57283 62056 ne
rect 57283 61994 58759 62056
tri 58759 61994 59042 62277 sw
tri 59042 61994 59325 62277 ne
rect 59325 62180 60832 62277
tri 60832 62180 61119 62467 sw
tri 61119 62180 61406 62467 ne
rect 61406 62465 62816 62467
tri 62816 62465 63101 62750 sw
tri 63101 62465 63386 62750 ne
rect 63386 62566 64997 62750
tri 64997 62566 65265 62834 sw
tri 65280 62566 65548 62834 ne
rect 65548 62566 71000 62834
rect 63386 62465 65265 62566
rect 61406 62180 63101 62465
tri 63101 62180 63386 62465 sw
tri 63386 62180 63671 62465 ne
rect 63671 62283 65265 62465
tri 65265 62283 65548 62566 sw
tri 65548 62283 65831 62566 ne
rect 65831 62283 71000 62566
rect 63671 62180 65548 62283
rect 59325 61994 61119 62180
rect 57283 61773 59042 61994
rect 55073 61720 57000 61773
rect 50800 61459 52519 61720
tri 50800 61375 50884 61459 ne
rect 50884 61432 52519 61459
tri 52519 61432 52807 61720 sw
tri 52807 61432 53095 61720 ne
rect 53095 61626 54787 61720
tri 54787 61626 54881 61720 sw
tri 55073 61626 55167 61720 ne
rect 55167 61626 57000 61720
rect 53095 61432 54881 61626
rect 50884 61375 52807 61432
tri 50600 61175 50800 61375 sw
tri 50884 61175 51084 61375 ne
rect 51084 61303 52807 61375
tri 52807 61303 52936 61432 sw
tri 53095 61303 53224 61432 ne
rect 53224 61340 54881 61432
tri 54881 61340 55167 61626 sw
tri 55167 61340 55453 61626 ne
rect 55453 61490 57000 61626
tri 57000 61490 57283 61773 sw
tri 57283 61490 57566 61773 ne
rect 57566 61711 59042 61773
tri 59042 61711 59325 61994 sw
tri 59325 61711 59608 61994 ne
rect 59608 61893 61119 61994
tri 61119 61893 61406 62180 sw
tri 61406 61893 61693 62180 ne
rect 61693 62085 63386 62180
tri 63386 62085 63481 62180 sw
tri 63671 62085 63766 62180 ne
rect 63766 62085 65548 62180
rect 61693 61893 63481 62085
rect 59608 61711 61406 61893
rect 57566 61526 59325 61711
tri 59325 61526 59510 61711 sw
tri 59608 61526 59793 61711 ne
rect 59793 61606 61406 61711
tri 61406 61606 61693 61893 sw
tri 61693 61606 61980 61893 ne
rect 61980 61800 63481 61893
tri 63481 61800 63766 62085 sw
tri 63766 61800 64051 62085 ne
rect 64051 62000 65548 62085
tri 65548 62000 65831 62283 sw
tri 65831 62000 66114 62283 ne
rect 66114 62000 71000 62283
rect 64051 61800 65831 62000
tri 65831 61800 66031 62000 sw
rect 61980 61606 63766 61800
rect 59793 61526 61693 61606
rect 57566 61490 59510 61526
rect 55453 61340 57283 61490
rect 53224 61303 55167 61340
rect 51084 61175 52936 61303
rect 49200 60891 50800 61175
tri 50800 60891 51084 61175 sw
tri 51084 60891 51368 61175 ne
rect 51368 61015 52936 61175
tri 52936 61015 53224 61303 sw
tri 53224 61015 53512 61303 ne
rect 53512 61054 55167 61303
tri 55167 61054 55453 61340 sw
tri 55453 61054 55739 61340 ne
rect 55739 61243 57283 61340
tri 57283 61243 57530 61490 sw
tri 57566 61243 57813 61490 ne
rect 57813 61243 59510 61490
tri 59510 61243 59793 61526 sw
tri 59793 61243 60076 61526 ne
rect 60076 61319 61693 61526
tri 61693 61319 61980 61606 sw
tri 61980 61319 62267 61606 ne
rect 62267 61515 63766 61606
tri 63766 61515 64051 61800 sw
tri 64051 61515 64336 61800 ne
rect 64336 61515 71000 61800
rect 62267 61319 64051 61515
rect 60076 61243 61980 61319
rect 55739 61054 57530 61243
rect 53512 61015 55453 61054
rect 51368 60891 53224 61015
rect 49200 60795 51084 60891
tri 49200 60710 49285 60795 ne
rect 49285 60784 51084 60795
tri 51084 60784 51191 60891 sw
tri 51368 60784 51475 60891 ne
rect 51475 60784 53224 60891
rect 49285 60710 51191 60784
tri 49000 60425 49285 60710 sw
tri 49285 60425 49570 60710 ne
rect 49570 60500 51191 60710
tri 51191 60500 51475 60784 sw
tri 51475 60500 51759 60784 ne
rect 51759 60727 53224 60784
tri 53224 60727 53512 61015 sw
tri 53512 60727 53800 61015 ne
rect 53800 60768 55453 61015
tri 55453 60768 55739 61054 sw
tri 55739 60768 56025 61054 ne
rect 56025 60960 57530 61054
tri 57530 60960 57813 61243 sw
tri 57813 60960 58096 61243 ne
rect 58096 60960 59793 61243
tri 59793 60960 60076 61243 sw
tri 60076 60960 60359 61243 ne
rect 60359 61154 61980 61243
tri 61980 61154 62145 61319 sw
tri 62267 61154 62432 61319 ne
rect 62432 61230 64051 61319
tri 64051 61230 64336 61515 sw
tri 64336 61230 64621 61515 ne
rect 64621 61230 71000 61515
rect 62432 61154 64336 61230
rect 60359 60960 62145 61154
rect 56025 60768 57813 60960
rect 53800 60727 55739 60768
rect 51759 60500 53512 60727
rect 49570 60425 51475 60500
rect 46000 60140 49285 60425
tri 49285 60140 49570 60425 sw
tri 49570 60140 49855 60425 ne
rect 49855 60404 51475 60425
tri 51475 60404 51571 60500 sw
tri 51759 60404 51855 60500 ne
rect 51855 60439 53512 60500
tri 53512 60439 53800 60727 sw
tri 53800 60439 54088 60727 ne
rect 54088 60482 55739 60727
tri 55739 60482 56025 60768 sw
tri 56025 60482 56311 60768 ne
rect 56311 60677 57813 60768
tri 57813 60677 58096 60960 sw
tri 58096 60677 58379 60960 ne
rect 58379 60863 60076 60960
tri 60076 60863 60173 60960 sw
tri 60359 60863 60456 60960 ne
rect 60456 60867 62145 60960
tri 62145 60867 62432 61154 sw
tri 62432 60867 62719 61154 ne
rect 62719 60970 64336 61154
tri 64336 60970 64596 61230 sw
tri 64621 60970 64881 61230 ne
rect 64881 60970 71000 61230
rect 62719 60867 64596 60970
rect 60456 60863 62432 60867
rect 58379 60677 60173 60863
rect 56311 60482 58096 60677
rect 54088 60439 56025 60482
rect 51855 60404 53800 60439
rect 49855 60140 51571 60404
rect 46000 59965 49570 60140
tri 49570 59965 49745 60140 sw
tri 49855 59965 50030 60140 ne
rect 50030 60120 51571 60140
tri 51571 60120 51855 60404 sw
tri 51855 60120 52139 60404 ne
rect 52139 60151 53800 60404
tri 53800 60151 54088 60439 sw
tri 54088 60151 54376 60439 ne
rect 54376 60312 56025 60439
tri 56025 60312 56195 60482 sw
tri 56311 60312 56481 60482 ne
rect 56481 60394 58096 60482
tri 58096 60394 58379 60677 sw
tri 58379 60394 58662 60677 ne
rect 58662 60580 60173 60677
tri 60173 60580 60456 60863 sw
tri 60456 60580 60739 60863 ne
rect 60739 60580 62432 60863
tri 62432 60580 62719 60867 sw
tri 62719 60580 63006 60867 ne
rect 63006 60685 64596 60867
tri 64596 60685 64881 60970 sw
tri 64881 60685 65166 60970 ne
rect 65166 60685 71000 60970
rect 63006 60580 64881 60685
rect 58662 60394 60456 60580
rect 56481 60312 58379 60394
rect 54376 60151 56195 60312
rect 52139 60120 54088 60151
rect 50030 60059 51855 60120
tri 51855 60059 51916 60120 sw
tri 52139 60059 52200 60120 ne
rect 52200 60059 54088 60120
rect 50030 59965 51916 60059
rect 46000 59680 49745 59965
tri 49745 59680 50030 59965 sw
tri 50030 59680 50315 59965 ne
rect 50315 59775 51916 59965
tri 51916 59775 52200 60059 sw
tri 52200 59775 52484 60059 ne
rect 52484 60028 54088 60059
tri 54088 60028 54211 60151 sw
tri 54376 60028 54499 60151 ne
rect 54499 60028 56195 60151
rect 52484 59775 54211 60028
rect 50315 59680 52200 59775
rect 46000 59461 50030 59680
tri 46000 59350 46111 59461 ne
rect 46111 59395 50030 59461
tri 50030 59395 50315 59680 sw
tri 50315 59395 50600 59680 ne
rect 50600 59491 52200 59680
tri 52200 59491 52484 59775 sw
tri 52484 59491 52768 59775 ne
rect 52768 59740 54211 59775
tri 54211 59740 54499 60028 sw
tri 54499 59740 54787 60028 ne
rect 54787 60026 56195 60028
tri 56195 60026 56481 60312 sw
tri 56481 60026 56767 60312 ne
rect 56767 60111 58379 60312
tri 58379 60111 58662 60394 sw
tri 58662 60111 58945 60394 ne
rect 58945 60297 60456 60394
tri 60456 60297 60739 60580 sw
tri 60739 60297 61022 60580 ne
rect 61022 60487 62719 60580
tri 62719 60487 62812 60580 sw
tri 63006 60487 63099 60580 ne
rect 63099 60487 64881 60580
rect 61022 60297 62812 60487
rect 58945 60111 60739 60297
rect 56767 60026 58662 60111
rect 54787 59740 56481 60026
tri 56481 59740 56767 60026 sw
tri 56767 59740 57053 60026 ne
rect 57053 59926 58662 60026
tri 58662 59926 58847 60111 sw
tri 58945 59926 59130 60111 ne
rect 59130 60014 60739 60111
tri 60739 60014 61022 60297 sw
tri 61022 60014 61305 60297 ne
rect 61305 60200 62812 60297
tri 62812 60200 63099 60487 sw
tri 63099 60200 63386 60487 ne
rect 63386 60400 64881 60487
tri 64881 60400 65166 60685 sw
tri 65166 60400 65451 60685 ne
rect 65451 60400 71000 60685
rect 63386 60200 65166 60400
tri 65166 60200 65366 60400 sw
rect 61305 60014 63099 60200
rect 59130 59926 61022 60014
rect 57053 59740 58847 59926
rect 52768 59491 54499 59740
rect 50600 59395 52484 59491
rect 46111 59350 50315 59395
tri 45800 59039 46111 59350 sw
tri 46111 59039 46422 59350 ne
rect 46422 59110 50315 59350
tri 50315 59110 50600 59395 sw
tri 50600 59110 50885 59395 ne
rect 50885 59207 52484 59395
tri 52484 59207 52768 59491 sw
tri 52768 59207 53052 59491 ne
rect 53052 59452 54499 59491
tri 54499 59452 54787 59740 sw
tri 54787 59452 55075 59740 ne
rect 55075 59646 56767 59740
tri 56767 59646 56861 59740 sw
tri 57053 59646 57147 59740 ne
rect 57147 59646 58847 59740
rect 55075 59452 56861 59646
rect 53052 59207 54787 59452
rect 50885 59110 52768 59207
rect 46422 59039 50600 59110
rect 42800 58728 46111 59039
tri 46111 58728 46422 59039 sw
tri 46422 58728 46733 59039 ne
rect 46733 59032 50600 59039
tri 50600 59032 50678 59110 sw
tri 50885 59032 50963 59110 ne
rect 50963 59088 52768 59110
tri 52768 59088 52887 59207 sw
tri 53052 59088 53171 59207 ne
rect 53171 59164 54787 59207
tri 54787 59164 55075 59452 sw
tri 55075 59164 55363 59452 ne
rect 55363 59360 56861 59452
tri 56861 59360 57147 59646 sw
tri 57147 59360 57433 59646 ne
rect 57433 59643 58847 59646
tri 58847 59643 59130 59926 sw
tri 59130 59643 59413 59926 ne
rect 59413 59731 61022 59926
tri 61022 59731 61305 60014 sw
tri 61305 59731 61588 60014 ne
rect 61588 59913 63099 60014
tri 63099 59913 63386 60200 sw
tri 63386 59913 63673 60200 ne
rect 63673 60120 71000 60200
rect 63673 59913 70613 60120
rect 61588 59731 63386 59913
rect 59413 59643 61305 59731
rect 57433 59360 59130 59643
tri 59130 59360 59413 59643 sw
tri 59413 59360 59696 59643 ne
rect 59696 59546 61305 59643
tri 61305 59546 61490 59731 sw
tri 61588 59546 61773 59731 ne
rect 61773 59626 63386 59731
tri 63386 59626 63673 59913 sw
tri 63673 59626 63960 59913 ne
rect 63960 59626 70613 59913
rect 61773 59546 63673 59626
rect 59696 59360 61490 59546
rect 55363 59164 57147 59360
rect 53171 59088 55075 59164
rect 50963 59032 52887 59088
rect 46733 58747 50678 59032
tri 50678 58747 50963 59032 sw
tri 50963 58747 51248 59032 ne
rect 51248 58804 52887 59032
tri 52887 58804 53171 59088 sw
tri 53171 58804 53455 59088 ne
rect 53455 58876 55075 59088
tri 55075 58876 55363 59164 sw
tri 55363 58876 55651 59164 ne
rect 55651 59074 57147 59164
tri 57147 59074 57433 59360 sw
tri 57433 59074 57719 59360 ne
rect 57719 59263 59413 59360
tri 59413 59263 59510 59360 sw
tri 59696 59263 59793 59360 ne
rect 59793 59263 61490 59360
tri 61490 59263 61773 59546 sw
tri 61773 59263 62056 59546 ne
rect 62056 59374 63673 59546
tri 63673 59374 63925 59626 sw
tri 63960 59374 64212 59626 ne
rect 64212 59374 70613 59626
rect 62056 59263 63925 59374
rect 57719 59074 59510 59263
rect 55651 58876 57433 59074
rect 53455 58804 55363 58876
rect 51248 58747 53171 58804
rect 46733 58728 50963 58747
rect 42800 58417 46422 58728
tri 46422 58417 46733 58728 sw
tri 46733 58417 47044 58728 ne
rect 47044 58462 50963 58728
tri 50963 58462 51248 58747 sw
tri 51248 58462 51533 58747 ne
rect 51533 58520 53171 58747
tri 53171 58520 53455 58804 sw
tri 53455 58520 53739 58804 ne
rect 53739 58716 55363 58804
tri 55363 58716 55523 58876 sw
tri 55651 58716 55811 58876 ne
rect 55811 58788 57433 58876
tri 57433 58788 57719 59074 sw
tri 57719 58788 58005 59074 ne
rect 58005 58980 59510 59074
tri 59510 58980 59793 59263 sw
tri 59793 58980 60076 59263 ne
rect 60076 58980 61773 59263
tri 61773 58980 62056 59263 sw
tri 62056 58980 62339 59263 ne
rect 62339 59087 63925 59263
tri 63925 59087 64212 59374 sw
tri 64212 59087 64499 59374 ne
rect 64499 59087 70613 59374
rect 62339 58980 64212 59087
rect 58005 58788 59793 58980
rect 55811 58716 57719 58788
rect 53739 58520 55523 58716
rect 51533 58462 53455 58520
rect 47044 58417 51248 58462
rect 42800 58106 46733 58417
tri 46733 58106 47044 58417 sw
tri 47044 58106 47355 58417 ne
rect 47355 58295 51248 58417
tri 51248 58295 51415 58462 sw
tri 51533 58295 51700 58462 ne
rect 51700 58424 53455 58462
tri 53455 58424 53551 58520 sw
tri 53739 58424 53835 58520 ne
rect 53835 58428 55523 58520
tri 55523 58428 55811 58716 sw
tri 55811 58428 56099 58716 ne
rect 56099 58502 57719 58716
tri 57719 58502 58005 58788 sw
tri 58005 58502 58291 58788 ne
rect 58291 58697 59793 58788
tri 59793 58697 60076 58980 sw
tri 60076 58697 60359 58980 ne
rect 60359 58883 62056 58980
tri 62056 58883 62153 58980 sw
tri 62339 58883 62436 58980 ne
rect 62436 58883 64212 58980
rect 60359 58697 62153 58883
rect 58291 58502 60076 58697
rect 56099 58428 58005 58502
rect 53835 58424 55811 58428
rect 51700 58295 53551 58424
rect 47355 58106 51415 58295
rect 42800 58097 47044 58106
tri 42600 57810 42800 58010 sw
tri 42800 57810 43087 58097 ne
rect 43087 57810 47044 58097
rect 41200 57523 42800 57810
tri 42800 57523 43087 57810 sw
tri 43087 57523 43374 57810 ne
rect 43374 57795 47044 57810
tri 47044 57795 47355 58106 sw
tri 47355 57795 47666 58106 ne
rect 47666 58010 51415 58106
tri 51415 58010 51700 58295 sw
tri 51700 58010 51985 58295 ne
rect 51985 58140 53551 58295
tri 53551 58140 53835 58424 sw
tri 53835 58140 54119 58424 ne
rect 54119 58140 55811 58424
tri 55811 58140 56099 58428 sw
tri 56099 58140 56387 58428 ne
rect 56387 58332 58005 58428
tri 58005 58332 58175 58502 sw
tri 58291 58332 58461 58502 ne
rect 58461 58414 60076 58502
tri 60076 58414 60359 58697 sw
tri 60359 58414 60642 58697 ne
rect 60642 58600 62153 58697
tri 62153 58600 62436 58883 sw
tri 62436 58600 62719 58883 ne
rect 62719 58800 64212 58883
tri 64212 58800 64499 59087 sw
tri 64499 58800 64786 59087 ne
rect 64786 58920 70613 59087
rect 70669 58920 71000 60120
rect 64786 58800 71000 58920
rect 62719 58600 64499 58800
tri 64499 58600 64699 58800 sw
rect 60642 58414 62436 58600
rect 58461 58332 60359 58414
rect 56387 58140 58175 58332
rect 51985 58010 53835 58140
rect 47666 57795 51700 58010
rect 43374 57704 47355 57795
tri 47355 57704 47446 57795 sw
tri 47666 57704 47757 57795 ne
rect 47757 57725 51700 57795
tri 51700 57725 51985 58010 sw
tri 51985 57725 52270 58010 ne
rect 52270 57856 53835 58010
tri 53835 57856 54119 58140 sw
tri 54119 57856 54403 58140 ne
rect 54403 58048 56099 58140
tri 56099 58048 56191 58140 sw
tri 56387 58048 56479 58140 ne
rect 56479 58048 58175 58140
rect 54403 57856 56191 58048
rect 52270 57725 54119 57856
rect 47757 57704 51985 57725
rect 43374 57523 47446 57704
rect 41200 57430 43087 57523
tri 41200 57338 41292 57430 ne
rect 41292 57338 43087 57430
tri 41000 57138 41200 57338 sw
tri 41292 57138 41492 57338 ne
rect 41492 57236 43087 57338
tri 43087 57236 43374 57523 sw
tri 43374 57236 43661 57523 ne
rect 43661 57393 47446 57523
tri 47446 57393 47757 57704 sw
tri 47757 57393 48068 57704 ne
rect 48068 57440 51985 57704
tri 51985 57440 52270 57725 sw
tri 52270 57440 52555 57725 ne
rect 52555 57572 54119 57725
tri 54119 57572 54403 57856 sw
tri 54403 57572 54687 57856 ne
rect 54687 57760 56191 57856
tri 56191 57760 56479 58048 sw
tri 56479 57760 56767 58048 ne
rect 56767 58046 58175 58048
tri 58175 58046 58461 58332 sw
tri 58461 58046 58747 58332 ne
rect 58747 58131 60359 58332
tri 60359 58131 60642 58414 sw
tri 60642 58131 60925 58414 ne
rect 60925 58317 62436 58414
tri 62436 58317 62719 58600 sw
tri 62719 58317 63002 58600 ne
rect 63002 58317 71000 58600
rect 60925 58131 62719 58317
rect 58747 58046 60642 58131
rect 56767 57760 58461 58046
tri 58461 57760 58747 58046 sw
tri 58747 57760 59033 58046 ne
rect 59033 57946 60642 58046
tri 60642 57946 60827 58131 sw
tri 60925 57946 61110 58131 ne
rect 61110 58034 62719 58131
tri 62719 58034 63002 58317 sw
tri 63002 58034 63285 58317 ne
rect 63285 58034 71000 58317
rect 61110 57946 63002 58034
rect 59033 57760 60827 57946
rect 54687 57572 56479 57760
rect 52555 57440 54403 57572
rect 48068 57393 52270 57440
rect 43661 57236 47757 57393
rect 41492 57138 43374 57236
rect 39600 57132 41200 57138
tri 41200 57132 41206 57138 sw
tri 41492 57132 41498 57138 ne
rect 41498 57132 43374 57138
rect 39600 56840 41206 57132
tri 41206 56840 41498 57132 sw
tri 41498 56840 41790 57132 ne
rect 41790 57034 43374 57132
tri 43374 57034 43576 57236 sw
tri 43661 57034 43863 57236 ne
rect 43863 57082 47757 57236
tri 47757 57082 48068 57393 sw
tri 48068 57082 48379 57393 ne
rect 48379 57155 52270 57393
tri 52270 57155 52555 57440 sw
tri 52555 57155 52840 57440 ne
rect 52840 57288 54403 57440
tri 54403 57288 54687 57572 sw
tri 54687 57288 54971 57572 ne
rect 54971 57472 56479 57572
tri 56479 57472 56767 57760 sw
tri 56767 57472 57055 57760 ne
rect 57055 57666 58747 57760
tri 58747 57666 58841 57760 sw
tri 59033 57666 59127 57760 ne
rect 59127 57666 60827 57760
rect 57055 57472 58841 57666
rect 54971 57288 56767 57472
rect 52840 57155 54687 57288
rect 48379 57110 52555 57155
tri 52555 57110 52600 57155 sw
tri 52840 57110 52885 57155 ne
rect 52885 57110 54687 57155
rect 48379 57082 52600 57110
rect 43863 57034 48068 57082
rect 41790 56840 43576 57034
rect 39600 56758 41498 56840
tri 39600 56665 39693 56758 ne
rect 39693 56752 41498 56758
tri 41498 56752 41586 56840 sw
tri 41790 56752 41878 56840 ne
rect 41878 56752 43576 56840
rect 39693 56665 41586 56752
tri 39400 56372 39693 56665 sw
tri 39693 56372 39986 56665 ne
rect 39986 56460 41586 56665
tri 41586 56460 41878 56752 sw
tri 41878 56460 42170 56752 ne
rect 42170 56747 43576 56752
tri 43576 56747 43863 57034 sw
tri 43863 56747 44150 57034 ne
rect 44150 56771 48068 57034
tri 48068 56771 48379 57082 sw
tri 48379 56771 48690 57082 ne
rect 48690 56825 52600 57082
tri 52600 56825 52885 57110 sw
tri 52885 56825 53170 57110 ne
rect 53170 57108 54687 57110
tri 54687 57108 54867 57288 sw
tri 54971 57108 55151 57288 ne
rect 55151 57184 56767 57288
tri 56767 57184 57055 57472 sw
tri 57055 57184 57343 57472 ne
rect 57343 57380 58841 57472
tri 58841 57380 59127 57666 sw
tri 59127 57380 59413 57666 ne
rect 59413 57663 60827 57666
tri 60827 57663 61110 57946 sw
tri 61110 57663 61393 57946 ne
rect 61393 57766 63002 57946
tri 63002 57766 63270 58034 sw
tri 63285 57766 63553 58034 ne
rect 63553 57766 71000 58034
rect 61393 57663 63270 57766
rect 59413 57380 61110 57663
tri 61110 57380 61393 57663 sw
tri 61393 57380 61676 57663 ne
rect 61676 57483 63270 57663
tri 63270 57483 63553 57766 sw
tri 63553 57483 63836 57766 ne
rect 63836 57483 71000 57766
rect 61676 57380 63553 57483
rect 57343 57184 59127 57380
rect 55151 57108 57055 57184
rect 53170 56825 54867 57108
rect 48690 56771 52885 56825
rect 44150 56747 48379 56771
rect 42170 56460 43863 56747
tri 43863 56460 44150 56747 sw
tri 44150 56460 44437 56747 ne
rect 44437 56460 48379 56747
tri 48379 56460 48690 56771 sw
tri 48690 56460 49001 56771 ne
rect 49001 56540 52885 56771
tri 52885 56540 53170 56825 sw
tri 53170 56540 53455 56825 ne
rect 53455 56824 54867 56825
tri 54867 56824 55151 57108 sw
tri 55151 56824 55435 57108 ne
rect 55435 56896 57055 57108
tri 57055 56896 57343 57184 sw
tri 57343 56896 57631 57184 ne
rect 57631 57094 59127 57184
tri 59127 57094 59413 57380 sw
tri 59413 57094 59699 57380 ne
rect 59699 57283 61393 57380
tri 61393 57283 61490 57380 sw
tri 61676 57283 61773 57380 ne
rect 61773 57283 63553 57380
rect 59699 57094 61490 57283
rect 57631 56896 59413 57094
rect 55435 56824 57343 56896
rect 53455 56540 55151 56824
tri 55151 56540 55435 56824 sw
tri 55435 56540 55719 56824 ne
rect 55719 56736 57343 56824
tri 57343 56736 57503 56896 sw
tri 57631 56736 57791 56896 ne
rect 57791 56808 59413 56896
tri 59413 56808 59699 57094 sw
tri 59699 56808 59985 57094 ne
rect 59985 57000 61490 57094
tri 61490 57000 61773 57283 sw
tri 61773 57000 62056 57283 ne
rect 62056 57200 63553 57283
tri 63553 57200 63836 57483 sw
tri 63836 57200 64119 57483 ne
rect 64119 57200 71000 57483
rect 62056 57000 63836 57200
tri 63836 57000 64036 57200 sw
rect 59985 56808 61773 57000
rect 57791 56736 59699 56808
rect 55719 56540 57503 56736
rect 49001 56460 53170 56540
tri 53170 56460 53250 56540 sw
tri 53455 56460 53535 56540 ne
rect 53535 56460 55435 56540
rect 39986 56372 41878 56460
rect 36400 56323 39693 56372
tri 39693 56323 39742 56372 sw
tri 39986 56323 40035 56372 ne
rect 40035 56323 41878 56372
rect 36400 56030 39742 56323
tri 39742 56030 40035 56323 sw
tri 40035 56030 40328 56323 ne
rect 40328 56322 41878 56323
tri 41878 56322 42016 56460 sw
tri 42170 56322 42308 56460 ne
rect 42308 56322 44150 56460
rect 40328 56030 42016 56322
tri 42016 56030 42308 56322 sw
tri 42308 56030 42600 56322 ne
rect 42600 56173 44150 56322
tri 44150 56173 44437 56460 sw
tri 44437 56173 44724 56460 ne
rect 44724 56173 48690 56460
rect 42600 56133 44437 56173
tri 44437 56133 44477 56173 sw
tri 44724 56133 44764 56173 ne
rect 44764 56149 48690 56173
tri 48690 56149 49001 56460 sw
tri 49001 56149 49312 56460 ne
rect 49312 56175 53250 56460
tri 53250 56175 53535 56460 sw
tri 53535 56175 53820 56460 ne
rect 53820 56444 55435 56460
tri 55435 56444 55531 56540 sw
tri 55719 56444 55815 56540 ne
rect 55815 56448 57503 56540
tri 57503 56448 57791 56736 sw
tri 57791 56448 58079 56736 ne
rect 58079 56522 59699 56736
tri 59699 56522 59985 56808 sw
tri 59985 56522 60271 56808 ne
rect 60271 56717 61773 56808
tri 61773 56717 62056 57000 sw
tri 62056 56717 62339 57000 ne
rect 62339 56910 71000 57000
rect 62339 56717 70613 56910
rect 60271 56522 62056 56717
rect 58079 56448 59985 56522
rect 55815 56444 57791 56448
rect 53820 56175 55531 56444
rect 49312 56160 53535 56175
tri 53535 56160 53550 56175 sw
tri 53820 56160 53835 56175 ne
rect 53835 56160 55531 56175
tri 55531 56160 55815 56444 sw
tri 55815 56160 56099 56444 ne
rect 56099 56160 57791 56444
tri 57791 56160 58079 56448 sw
tri 58079 56160 58367 56448 ne
rect 58367 56352 59985 56448
tri 59985 56352 60155 56522 sw
tri 60271 56352 60441 56522 ne
rect 60441 56434 62056 56522
tri 62056 56434 62339 56717 sw
tri 62339 56434 62622 56717 ne
rect 62622 56434 70613 56717
rect 60441 56352 62339 56434
rect 58367 56160 60155 56352
rect 49312 56149 53550 56160
rect 44764 56133 49001 56149
rect 42600 56030 44477 56133
rect 36400 55737 40035 56030
tri 40035 55737 40328 56030 sw
tri 40328 55737 40621 56030 ne
rect 40621 55738 42308 56030
tri 42308 55738 42600 56030 sw
tri 42600 55738 42892 56030 ne
rect 42892 55846 44477 56030
tri 44477 55846 44764 56133 sw
tri 44764 55846 45051 56133 ne
rect 45051 55870 49001 56133
tri 49001 55870 49280 56149 sw
tri 49312 55870 49591 56149 ne
rect 49591 55875 53550 56149
tri 53550 55875 53835 56160 sw
tri 53835 55875 54120 56160 ne
rect 54120 55876 55815 56160
tri 55815 55876 56099 56160 sw
tri 56099 55876 56383 56160 ne
rect 56383 56068 58079 56160
tri 58079 56068 58171 56160 sw
tri 58367 56068 58459 56160 ne
rect 58459 56068 60155 56160
rect 56383 55876 58171 56068
rect 54120 55875 56099 55876
rect 49591 55870 53835 55875
rect 45051 55846 49280 55870
rect 42892 55738 44764 55846
rect 40621 55737 42600 55738
rect 36400 55444 40328 55737
tri 40328 55444 40621 55737 sw
tri 40621 55444 40914 55737 ne
rect 40914 55446 42600 55737
tri 42600 55446 42892 55738 sw
tri 42892 55446 43184 55738 ne
rect 43184 55559 44764 55738
tri 44764 55559 45051 55846 sw
tri 45051 55559 45338 55846 ne
rect 45338 55559 49280 55846
tri 49280 55559 49591 55870 sw
tri 49591 55559 49902 55870 ne
rect 49902 55590 53835 55870
tri 53835 55590 54120 55875 sw
tri 54120 55590 54405 55875 ne
rect 54405 55592 56099 55875
tri 56099 55592 56383 55876 sw
tri 56383 55592 56667 55876 ne
rect 56667 55780 58171 55876
tri 58171 55780 58459 56068 sw
tri 58459 55780 58747 56068 ne
rect 58747 56066 60155 56068
tri 60155 56066 60441 56352 sw
tri 60441 56066 60727 56352 ne
rect 60727 56166 62339 56352
tri 62339 56166 62607 56434 sw
tri 62622 56166 62890 56434 ne
rect 62890 56166 70613 56434
rect 60727 56066 62607 56166
rect 58747 55780 60441 56066
tri 60441 55780 60727 56066 sw
tri 60727 55780 61013 56066 ne
rect 61013 55883 62607 56066
tri 62607 55883 62890 56166 sw
tri 62890 55883 63173 56166 ne
rect 63173 55883 70613 56166
rect 61013 55780 62890 55883
rect 56667 55592 58459 55780
rect 54405 55590 56383 55592
rect 49902 55559 54120 55590
rect 43184 55446 45051 55559
rect 40914 55444 42892 55446
tri 42892 55444 42894 55446 sw
tri 43184 55444 43186 55446 ne
rect 43186 55444 45051 55446
rect 36400 55421 40621 55444
tri 36400 55324 36497 55421 ne
rect 36497 55324 40621 55421
tri 36200 55027 36497 55324 sw
tri 36497 55027 36794 55324 ne
rect 36794 55153 40621 55324
tri 40621 55153 40912 55444 sw
tri 40914 55153 41205 55444 ne
rect 41205 55153 42894 55444
rect 36794 55027 40912 55153
rect 33200 54730 36497 55027
tri 36497 54730 36794 55027 sw
tri 36794 54730 37091 55027 ne
rect 37091 54860 40912 55027
tri 40912 54860 41205 55153 sw
tri 41205 54860 41498 55153 ne
rect 41498 55152 42894 55153
tri 42894 55152 43186 55444 sw
tri 43186 55152 43478 55444 ne
rect 43478 55272 45051 55444
tri 45051 55272 45338 55559 sw
tri 45338 55272 45625 55559 ne
rect 45625 55272 49591 55559
rect 43478 55152 45338 55272
rect 41498 54860 43186 55152
tri 43186 54860 43478 55152 sw
tri 43478 54860 43770 55152 ne
rect 43770 54985 45338 55152
tri 45338 54985 45625 55272 sw
tri 45625 54985 45912 55272 ne
rect 45912 55248 49591 55272
tri 49591 55248 49902 55559 sw
tri 49902 55248 50213 55559 ne
rect 50213 55353 54120 55559
tri 54120 55353 54357 55590 sw
tri 54405 55353 54642 55590 ne
rect 54642 55353 56383 55590
rect 50213 55248 54357 55353
rect 45912 54985 49902 55248
rect 43770 54860 45625 54985
rect 37091 54730 41205 54860
rect 33200 54674 36794 54730
tri 36794 54674 36850 54730 sw
tri 37091 54674 37147 54730 ne
rect 37147 54674 41205 54730
rect 33200 54377 36850 54674
tri 36850 54377 37147 54674 sw
tri 37147 54377 37444 54674 ne
rect 37444 54567 41205 54674
tri 41205 54567 41498 54860 sw
tri 41498 54567 41791 54860 ne
rect 41791 54772 43478 54860
tri 43478 54772 43566 54860 sw
tri 43770 54772 43858 54860 ne
rect 43858 54772 45625 54860
rect 41791 54567 43566 54772
rect 37444 54480 41498 54567
tri 41498 54480 41585 54567 sw
tri 41791 54480 41878 54567 ne
rect 41878 54480 43566 54567
tri 43566 54480 43858 54772 sw
tri 43858 54480 44150 54772 ne
rect 44150 54767 45625 54772
tri 45625 54767 45843 54985 sw
tri 45912 54767 46130 54985 ne
rect 46130 54937 49902 54985
tri 49902 54937 50213 55248 sw
tri 50213 54937 50524 55248 ne
rect 50524 55068 54357 55248
tri 54357 55068 54642 55353 sw
tri 54642 55068 54927 55353 ne
rect 54927 55308 56383 55353
tri 56383 55308 56667 55592 sw
tri 56667 55308 56951 55592 ne
rect 56951 55492 58459 55592
tri 58459 55492 58747 55780 sw
tri 58747 55492 59035 55780 ne
rect 59035 55686 60727 55780
tri 60727 55686 60821 55780 sw
tri 61013 55686 61107 55780 ne
rect 61107 55686 62890 55780
rect 59035 55492 60821 55686
rect 56951 55308 58747 55492
rect 54927 55128 56667 55308
tri 56667 55128 56847 55308 sw
tri 56951 55128 57131 55308 ne
rect 57131 55204 58747 55308
tri 58747 55204 59035 55492 sw
tri 59035 55204 59323 55492 ne
rect 59323 55400 60821 55492
tri 60821 55400 61107 55686 sw
tri 61107 55400 61393 55686 ne
rect 61393 55600 62890 55686
tri 62890 55600 63173 55883 sw
tri 63173 55600 63456 55883 ne
rect 63456 55710 70613 55883
rect 70669 55710 71000 56910
rect 63456 55600 71000 55710
rect 61393 55400 63173 55600
tri 63173 55400 63373 55600 sw
rect 59323 55204 61107 55400
rect 57131 55128 59035 55204
rect 54927 55068 56847 55128
rect 50524 54937 54642 55068
rect 46130 54767 50213 54937
rect 44150 54480 45843 54767
tri 45843 54480 46130 54767 sw
tri 46130 54480 46417 54767 ne
rect 46417 54626 50213 54767
tri 50213 54626 50524 54937 sw
tri 50524 54626 50835 54937 ne
rect 50835 54783 54642 54937
tri 54642 54783 54927 55068 sw
tri 54927 54783 55212 55068 ne
rect 55212 54844 56847 55068
tri 56847 54844 57131 55128 sw
tri 57131 54844 57415 55128 ne
rect 57415 54916 59035 55128
tri 59035 54916 59323 55204 sw
tri 59323 54916 59611 55204 ne
rect 59611 55114 61107 55204
tri 61107 55114 61393 55400 sw
tri 61393 55114 61679 55400 ne
rect 61679 55302 71000 55400
rect 61679 55114 70613 55302
rect 59611 54916 61393 55114
rect 57415 54844 59323 54916
rect 55212 54783 57131 54844
rect 50835 54626 54927 54783
rect 46417 54480 50524 54626
rect 37444 54377 41585 54480
rect 33200 54080 37147 54377
tri 37147 54080 37444 54377 sw
tri 37444 54080 37741 54377 ne
rect 37741 54187 41585 54377
tri 41585 54187 41878 54480 sw
tri 41878 54187 42171 54480 ne
rect 42171 54188 43858 54480
tri 43858 54188 44150 54480 sw
tri 44150 54188 44442 54480 ne
rect 44442 54193 46130 54480
tri 46130 54193 46417 54480 sw
tri 46417 54193 46704 54480 ne
rect 46704 54315 50524 54480
tri 50524 54315 50835 54626 sw
tri 50835 54315 51146 54626 ne
rect 51146 54498 54927 54626
tri 54927 54498 55212 54783 sw
tri 55212 54498 55497 54783 ne
rect 55497 54560 57131 54783
tri 57131 54560 57415 54844 sw
tri 57415 54560 57699 54844 ne
rect 57699 54756 59323 54844
tri 59323 54756 59483 54916 sw
tri 59611 54756 59771 54916 ne
rect 59771 54828 61393 54916
tri 61393 54828 61679 55114 sw
tri 61679 54828 61965 55114 ne
rect 61965 54828 70613 55114
rect 59771 54756 61679 54828
rect 57699 54560 59483 54756
rect 55497 54498 57415 54560
rect 51146 54315 55212 54498
rect 46704 54193 50835 54315
rect 44442 54188 46417 54193
rect 42171 54187 44150 54188
rect 37741 54080 41878 54187
tri 33200 53992 33288 54080 ne
rect 33288 53992 37444 54080
tri 33000 53704 33288 53992 sw
tri 33288 53704 33576 53992 ne
rect 33576 53783 37444 53992
tri 37444 53783 37741 54080 sw
tri 37741 53783 38038 54080 ne
rect 38038 53962 41878 54080
tri 41878 53962 42103 54187 sw
tri 42171 53962 42396 54187 ne
rect 42396 53962 44150 54187
rect 38038 53783 42103 53962
rect 33576 53704 37741 53783
rect 30000 53416 33288 53704
tri 33288 53416 33576 53704 sw
tri 33576 53416 33864 53704 ne
rect 33864 53486 37741 53704
tri 37741 53486 38038 53783 sw
tri 38038 53486 38335 53783 ne
rect 38335 53669 42103 53783
tri 42103 53669 42396 53962 sw
tri 42396 53669 42689 53962 ne
rect 42689 53896 44150 53962
tri 44150 53896 44442 54188 sw
tri 44442 53896 44734 54188 ne
rect 44734 53906 46417 54188
tri 46417 53906 46704 54193 sw
tri 46704 53906 46991 54193 ne
rect 46991 54004 50835 54193
tri 50835 54004 51146 54315 sw
tri 51146 54004 51457 54315 ne
rect 51457 54213 55212 54315
tri 55212 54213 55497 54498 sw
tri 55497 54213 55782 54498 ne
rect 55782 54464 57415 54498
tri 57415 54464 57511 54560 sw
tri 57699 54464 57795 54560 ne
rect 57795 54468 59483 54560
tri 59483 54468 59771 54756 sw
tri 59771 54468 60059 54756 ne
rect 60059 54572 61679 54756
tri 61679 54572 61935 54828 sw
tri 61965 54572 62221 54828 ne
rect 62221 54572 70613 54828
rect 60059 54468 61935 54572
rect 57795 54464 59771 54468
rect 55782 54213 57511 54464
rect 51457 54180 55497 54213
tri 55497 54180 55530 54213 sw
tri 55782 54180 55815 54213 ne
rect 55815 54180 57511 54213
tri 57511 54180 57795 54464 sw
tri 57795 54180 58079 54464 ne
rect 58079 54180 59771 54464
tri 59771 54180 60059 54468 sw
tri 60059 54180 60347 54468 ne
rect 60347 54286 61935 54468
tri 61935 54286 62221 54572 sw
tri 62221 54286 62507 54572 ne
rect 62507 54286 70613 54572
rect 60347 54180 62221 54286
rect 51457 54004 55530 54180
rect 46991 53906 51146 54004
rect 44734 53896 46704 53906
rect 42689 53669 44442 53896
rect 38335 53486 42396 53669
rect 33864 53416 38038 53486
rect 30000 53128 33576 53416
tri 33576 53128 33864 53416 sw
tri 33864 53128 34152 53416 ne
rect 34152 53189 38038 53416
tri 38038 53189 38335 53486 sw
tri 38335 53189 38632 53486 ne
rect 38632 53376 42396 53486
tri 42396 53376 42689 53669 sw
tri 42689 53376 42982 53669 ne
rect 42982 53604 44442 53669
tri 44442 53604 44734 53896 sw
tri 44734 53604 45026 53896 ne
rect 45026 53619 46704 53896
tri 46704 53619 46991 53906 sw
tri 46991 53619 47278 53906 ne
rect 47278 53744 51146 53906
tri 51146 53744 51406 54004 sw
tri 51457 53744 51717 54004 ne
rect 51717 53895 55530 54004
tri 55530 53895 55815 54180 sw
tri 55815 53895 56100 54180 ne
rect 56100 53896 57795 54180
tri 57795 53896 58079 54180 sw
tri 58079 53896 58363 54180 ne
rect 58363 54088 60059 54180
tri 60059 54088 60151 54180 sw
tri 60347 54088 60439 54180 ne
rect 60439 54088 62221 54180
rect 58363 53896 60151 54088
rect 56100 53895 58079 53896
rect 51717 53744 55815 53895
rect 47278 53619 51406 53744
rect 45026 53604 46991 53619
rect 42982 53464 44734 53604
tri 44734 53464 44874 53604 sw
tri 45026 53464 45166 53604 ne
rect 45166 53464 46991 53604
rect 42982 53376 44874 53464
rect 38632 53189 42689 53376
rect 34152 53128 38335 53189
rect 30000 52840 33864 53128
tri 33864 52840 34152 53128 sw
tri 34152 52840 34440 53128 ne
rect 34440 52892 38335 53128
tri 38335 52892 38632 53189 sw
tri 38632 52892 38929 53189 ne
rect 38929 53083 42689 53189
tri 42689 53083 42982 53376 sw
tri 42982 53083 43275 53376 ne
rect 43275 53172 44874 53376
tri 44874 53172 45166 53464 sw
tri 45166 53172 45458 53464 ne
rect 45458 53361 46991 53464
tri 46991 53361 47249 53619 sw
tri 47278 53361 47536 53619 ne
rect 47536 53433 51406 53619
tri 51406 53433 51717 53744 sw
tri 51717 53433 52028 53744 ne
rect 52028 53610 55815 53744
tri 55815 53610 56100 53895 sw
tri 56100 53610 56385 53895 ne
rect 56385 53612 58079 53895
tri 58079 53612 58363 53896 sw
tri 58363 53612 58647 53896 ne
rect 58647 53800 60151 53896
tri 60151 53800 60439 54088 sw
tri 60439 53800 60727 54088 ne
rect 60727 54000 62221 54088
tri 62221 54000 62507 54286 sw
tri 62507 54000 62793 54286 ne
rect 62793 54102 70613 54286
rect 70669 54102 71000 55302
rect 62793 54000 71000 54102
rect 60727 53800 62507 54000
tri 62507 53800 62707 54000 sw
rect 58647 53612 60439 53800
rect 56385 53610 58363 53612
rect 52028 53433 56100 53610
rect 47536 53361 51717 53433
rect 45458 53172 47249 53361
rect 43275 53083 45166 53172
rect 38929 52892 42982 53083
rect 34440 52840 38632 52892
rect 30000 52748 34152 52840
tri 30000 52654 30094 52748 ne
rect 30094 52660 34152 52748
tri 34152 52660 34332 52840 sw
tri 34440 52660 34620 52840 ne
rect 34620 52660 38632 52840
rect 30094 52654 34332 52660
tri 29800 52360 30094 52654 sw
tri 30094 52360 30388 52654 ne
rect 30388 52372 34332 52654
tri 34332 52372 34620 52660 sw
tri 34620 52372 34908 52660 ne
rect 34908 52595 38632 52660
tri 38632 52595 38929 52892 sw
tri 38929 52595 39226 52892 ne
rect 39226 52793 42982 52892
tri 42982 52793 43272 53083 sw
tri 43275 52793 43565 53083 ne
rect 43565 52880 45166 53083
tri 45166 52880 45458 53172 sw
tri 45458 52880 45750 53172 ne
rect 45750 53074 47249 53172
tri 47249 53074 47536 53361 sw
tri 47536 53074 47823 53361 ne
rect 47823 53122 51717 53361
tri 51717 53122 52028 53433 sw
tri 52028 53122 52339 53433 ne
rect 52339 53325 56100 53433
tri 56100 53325 56385 53610 sw
tri 56385 53325 56670 53610 ne
rect 56670 53328 58363 53610
tri 58363 53328 58647 53612 sw
tri 58647 53328 58931 53612 ne
rect 58931 53512 60439 53612
tri 60439 53512 60727 53800 sw
tri 60727 53512 61015 53800 ne
rect 61015 53722 71000 53800
rect 61015 53512 70613 53722
rect 58931 53328 60727 53512
rect 56670 53325 58647 53328
rect 52339 53150 56385 53325
tri 56385 53150 56560 53325 sw
tri 56670 53150 56845 53325 ne
rect 56845 53150 58647 53325
rect 52339 53122 56560 53150
rect 47823 53074 52028 53122
rect 45750 52880 47536 53074
rect 43565 52793 45458 52880
rect 39226 52595 43272 52793
rect 34908 52494 38929 52595
tri 38929 52494 39030 52595 sw
tri 39226 52494 39327 52595 ne
rect 39327 52500 43272 52595
tri 43272 52500 43565 52793 sw
tri 43565 52500 43858 52793 ne
rect 43858 52792 45458 52793
tri 45458 52792 45546 52880 sw
tri 45750 52792 45838 52880 ne
rect 45838 52792 47536 52880
rect 43858 52500 45546 52792
tri 45546 52500 45838 52792 sw
tri 45838 52500 46130 52792 ne
rect 46130 52787 47536 52792
tri 47536 52787 47823 53074 sw
tri 47823 52787 48110 53074 ne
rect 48110 52811 52028 53074
tri 52028 52811 52339 53122 sw
tri 52339 52811 52650 53122 ne
rect 52650 52865 56560 53122
tri 56560 52865 56845 53150 sw
tri 56845 52865 57130 53150 ne
rect 57130 53148 58647 53150
tri 58647 53148 58827 53328 sw
tri 58931 53148 59111 53328 ne
rect 59111 53224 60727 53328
tri 60727 53224 61015 53512 sw
tri 61015 53224 61303 53512 ne
rect 61303 53224 70613 53512
rect 59111 53148 61015 53224
rect 57130 52865 58827 53148
rect 52650 52811 56845 52865
rect 48110 52787 52339 52811
rect 46130 52500 47823 52787
tri 47823 52500 48110 52787 sw
tri 48110 52500 48397 52787 ne
rect 48397 52500 52339 52787
tri 52339 52500 52650 52811 sw
tri 52650 52500 52961 52811 ne
rect 52961 52580 56845 52811
tri 56845 52580 57130 52865 sw
tri 57130 52580 57415 52865 ne
rect 57415 52864 58827 52865
tri 58827 52864 59111 53148 sw
tri 59111 52864 59395 53148 ne
rect 59395 52976 61015 53148
tri 61015 52976 61263 53224 sw
tri 61303 52976 61551 53224 ne
rect 61551 52976 70613 53224
rect 59395 52864 61263 52976
rect 57415 52580 59111 52864
tri 59111 52580 59395 52864 sw
tri 59395 52580 59679 52864 ne
rect 59679 52688 61263 52864
tri 61263 52688 61551 52976 sw
tri 61551 52688 61839 52976 ne
rect 61839 52688 70613 52976
rect 59679 52580 61551 52688
rect 52961 52500 57130 52580
tri 57130 52500 57210 52580 sw
tri 57415 52500 57495 52580 ne
rect 57495 52500 59395 52580
rect 39327 52494 43565 52500
rect 34908 52372 39030 52494
rect 30388 52360 34620 52372
rect 26800 52066 30094 52360
tri 30094 52066 30388 52360 sw
tri 30388 52066 30682 52360 ne
rect 30682 52084 34620 52360
tri 34620 52084 34908 52372 sw
tri 34908 52084 35196 52372 ne
rect 35196 52197 39030 52372
tri 39030 52197 39327 52494 sw
tri 39327 52197 39624 52494 ne
rect 39624 52207 43565 52494
tri 43565 52207 43858 52500 sw
tri 43858 52207 44151 52500 ne
rect 44151 52208 45838 52500
tri 45838 52208 46130 52500 sw
tri 46130 52208 46422 52500 ne
rect 46422 52213 48110 52500
tri 48110 52213 48397 52500 sw
tri 48397 52213 48684 52500 ne
rect 48684 52213 52650 52500
rect 46422 52208 48397 52213
rect 44151 52207 46130 52208
rect 39624 52197 43858 52207
rect 35196 52084 39327 52197
rect 30682 52066 34908 52084
rect 26800 51998 30388 52066
tri 30388 51998 30456 52066 sw
tri 30682 51998 30750 52066 ne
rect 30750 51998 34908 52066
rect 26800 51704 30456 51998
tri 30456 51704 30750 51998 sw
tri 30750 51704 31044 51998 ne
rect 31044 51796 34908 51998
tri 34908 51796 35196 52084 sw
tri 35196 51796 35484 52084 ne
rect 35484 51900 39327 52084
tri 39327 51900 39624 52197 sw
tri 39624 51900 39921 52197 ne
rect 39921 51914 43858 52197
tri 43858 51914 44151 52207 sw
tri 44151 51914 44444 52207 ne
rect 44444 51916 46130 52207
tri 46130 51916 46422 52208 sw
tri 46422 51916 46714 52208 ne
rect 46714 51926 48397 52208
tri 48397 51926 48684 52213 sw
tri 48684 51926 48971 52213 ne
rect 48971 52189 52650 52213
tri 52650 52189 52961 52500 sw
tri 52961 52189 53272 52500 ne
rect 53272 52215 57210 52500
tri 57210 52215 57495 52500 sw
tri 57495 52215 57780 52500 ne
rect 57780 52484 59395 52500
tri 59395 52484 59491 52580 sw
tri 59679 52484 59775 52580 ne
rect 59775 52484 61551 52580
rect 57780 52215 59491 52484
rect 53272 52200 57495 52215
tri 57495 52200 57510 52215 sw
tri 57780 52200 57795 52215 ne
rect 57795 52200 59491 52215
tri 59491 52200 59775 52484 sw
tri 59775 52200 60059 52484 ne
rect 60059 52400 61551 52484
tri 61551 52400 61839 52688 sw
tri 61839 52400 62127 52688 ne
rect 62127 52522 70613 52688
rect 70669 52522 71000 53722
rect 62127 52400 71000 52522
rect 60059 52200 61839 52400
tri 61839 52200 62039 52400 sw
rect 53272 52189 57510 52200
rect 48971 51928 52961 52189
tri 52961 51928 53222 52189 sw
tri 53272 51928 53533 52189 ne
rect 53533 51928 57510 52189
rect 48971 51926 53222 51928
rect 46714 51916 48684 51926
rect 44444 51914 46422 51916
rect 39921 51906 44151 51914
tri 44151 51906 44159 51914 sw
tri 44444 51906 44452 51914 ne
rect 44452 51906 46422 51914
rect 39921 51900 44159 51906
rect 35484 51796 39624 51900
rect 31044 51704 35196 51796
rect 26800 51410 30750 51704
tri 30750 51410 31044 51704 sw
tri 31044 51410 31338 51704 ne
rect 31338 51508 35196 51704
tri 35196 51508 35484 51796 sw
tri 35484 51508 35772 51796 ne
rect 35772 51603 39624 51796
tri 39624 51603 39921 51900 sw
tri 39921 51603 40218 51900 ne
rect 40218 51613 44159 51900
tri 44159 51613 44452 51906 sw
tri 44452 51613 44745 51906 ne
rect 44745 51624 46422 51906
tri 46422 51624 46714 51916 sw
tri 46714 51624 47006 51916 ne
rect 47006 51880 48684 51916
tri 48684 51880 48730 51926 sw
tri 48971 51880 49017 51926 ne
rect 49017 51880 53222 51926
rect 47006 51624 48730 51880
rect 44745 51613 46714 51624
rect 40218 51603 44452 51613
rect 35772 51508 39921 51603
rect 31338 51410 35484 51508
tri 26600 51120 26800 51320 sw
tri 26800 51120 27090 51410 ne
rect 27090 51120 31044 51410
rect 25200 50830 26800 51120
tri 26800 50830 27090 51120 sw
tri 27090 50830 27380 51120 ne
rect 27380 51116 31044 51120
tri 31044 51116 31338 51410 sw
tri 31338 51116 31632 51410 ne
rect 31632 51220 35484 51410
tri 35484 51220 35772 51508 sw
tri 35772 51220 36060 51508 ne
rect 36060 51306 39921 51508
tri 39921 51306 40218 51603 sw
tri 40218 51306 40515 51603 ne
rect 40515 51320 44452 51603
tri 44452 51320 44745 51613 sw
tri 44745 51320 45038 51613 ne
rect 45038 51405 46714 51613
tri 46714 51405 46933 51624 sw
tri 47006 51484 47146 51624 ne
rect 47146 51593 48730 51624
tri 48730 51593 49017 51880 sw
tri 49017 51593 49304 51880 ne
rect 49304 51617 53222 51880
tri 53222 51617 53533 51928 sw
tri 53533 51617 53844 51928 ne
rect 53844 51915 57510 51928
tri 57510 51915 57795 52200 sw
tri 57795 51915 58080 52200 ne
rect 58080 51916 59775 52200
tri 59775 51916 60059 52200 sw
tri 60059 51916 60343 52200 ne
rect 60343 51916 71000 52200
rect 58080 51915 60059 51916
rect 53844 51630 57795 51915
tri 57795 51630 58080 51915 sw
tri 58080 51630 58365 51915 ne
rect 58365 51632 60059 51915
tri 60059 51632 60343 51916 sw
tri 60343 51632 60627 51916 ne
rect 60627 51632 71000 51916
rect 58365 51630 60343 51632
rect 53844 51617 58080 51630
rect 49304 51593 53533 51617
rect 47146 51484 49017 51593
rect 45038 51320 46933 51405
rect 40515 51306 44745 51320
tri 44745 51306 44759 51320 sw
tri 45038 51306 45052 51320 ne
rect 45052 51306 46933 51320
rect 36060 51220 40218 51306
rect 31632 51116 35772 51220
rect 27380 50830 31338 51116
rect 25200 50740 27090 50830
tri 25200 50651 25289 50740 ne
rect 25289 50651 27090 50740
tri 25000 50451 25200 50651 sw
tri 25289 50451 25489 50651 ne
rect 25489 50650 27090 50651
tri 27090 50650 27270 50830 sw
tri 27380 50650 27560 50830 ne
rect 27560 50822 31338 50830
tri 31338 50822 31632 51116 sw
tri 31632 50822 31926 51116 ne
rect 31926 50932 35772 51116
tri 35772 50932 36060 51220 sw
tri 36060 50932 36348 51220 ne
rect 36348 51009 40218 51220
tri 40218 51009 40515 51306 sw
tri 40515 51009 40812 51306 ne
rect 40812 51013 44759 51306
tri 44759 51013 45052 51306 sw
tri 45052 51013 45345 51306 ne
rect 45345 51192 46933 51306
tri 46933 51192 47146 51405 sw
tri 47146 51192 47438 51484 ne
rect 47438 51306 49017 51484
tri 49017 51306 49304 51593 sw
tri 49304 51306 49591 51593 ne
rect 49591 51306 53533 51593
tri 53533 51306 53844 51617 sw
tri 53844 51306 54155 51617 ne
rect 54155 51345 58080 51617
tri 58080 51345 58365 51630 sw
tri 58365 51345 58650 51630 ne
rect 58650 51368 60343 51630
tri 60343 51368 60607 51632 sw
tri 60627 51368 60891 51632 ne
rect 60891 51368 71000 51632
rect 58650 51345 60607 51368
rect 54155 51306 58365 51345
rect 47438 51192 49304 51306
rect 45345 51013 47146 51192
rect 40812 51009 45052 51013
rect 36348 50932 40515 51009
rect 31926 50822 36060 50932
rect 27560 50764 31632 50822
tri 31632 50764 31690 50822 sw
tri 31926 50764 31984 50822 ne
rect 31984 50764 36060 50822
rect 27560 50650 31690 50764
rect 25489 50451 27270 50650
rect 23600 50360 25200 50451
tri 25200 50360 25291 50451 sw
tri 25489 50360 25580 50451 ne
rect 25580 50360 27270 50451
tri 27270 50360 27560 50650 sw
tri 27560 50360 27850 50650 ne
rect 27850 50470 31690 50650
tri 31690 50470 31984 50764 sw
tri 31984 50470 32278 50764 ne
rect 32278 50644 36060 50764
tri 36060 50644 36348 50932 sw
tri 36348 50644 36636 50932 ne
rect 36636 50770 40515 50932
tri 40515 50770 40754 51009 sw
tri 40812 50770 41051 51009 ne
rect 41051 50900 45052 51009
tri 45052 50900 45165 51013 sw
tri 45345 50900 45458 51013 ne
rect 45458 50900 47146 51013
tri 47146 50900 47438 51192 sw
tri 47438 50900 47730 51192 ne
rect 47730 51019 49304 51192
tri 49304 51019 49591 51306 sw
tri 49591 51019 49878 51306 ne
rect 49878 51019 53844 51306
rect 47730 50900 49591 51019
rect 41051 50770 45165 50900
rect 36636 50644 40754 50770
rect 32278 50470 36348 50644
rect 27850 50360 31984 50470
rect 23600 50071 25291 50360
tri 25291 50071 25580 50360 sw
tri 25580 50071 25869 50360 ne
rect 25869 50071 27560 50360
tri 23600 49974 23697 50071 ne
rect 23697 49974 25580 50071
tri 23400 49677 23697 49974 sw
tri 23697 49677 23994 49974 ne
rect 23994 49918 25580 49974
tri 25580 49918 25733 50071 sw
tri 25869 49918 26022 50071 ne
rect 26022 50070 27560 50071
tri 27560 50070 27850 50360 sw
tri 27850 50070 28140 50360 ne
rect 28140 50176 31984 50360
tri 31984 50176 32278 50470 sw
tri 32278 50176 32572 50470 ne
rect 32572 50464 36348 50470
tri 36348 50464 36528 50644 sw
tri 36636 50464 36816 50644 ne
rect 36816 50473 40754 50644
tri 40754 50473 41051 50770 sw
tri 41051 50473 41348 50770 ne
rect 41348 50607 45165 50770
tri 45165 50607 45458 50900 sw
tri 45458 50607 45751 50900 ne
rect 45751 50812 47438 50900
tri 47438 50812 47526 50900 sw
tri 47730 50812 47818 50900 ne
rect 47818 50812 49591 50900
rect 45751 50607 47526 50812
rect 41348 50473 45458 50607
rect 36816 50464 41051 50473
rect 32572 50176 36528 50464
tri 36528 50176 36816 50464 sw
tri 36816 50176 37104 50464 ne
rect 37104 50176 41051 50464
tri 41051 50176 41348 50473 sw
tri 41348 50176 41645 50473 ne
rect 41645 50360 45458 50473
tri 45458 50360 45705 50607 sw
tri 45751 50360 45998 50607 ne
rect 45998 50520 47526 50607
tri 47526 50520 47818 50812 sw
tri 47818 50520 48110 50812 ne
rect 48110 50732 49591 50812
tri 49591 50732 49878 51019 sw
tri 49878 50732 50165 51019 ne
rect 50165 50995 53844 51019
tri 53844 50995 54155 51306 sw
tri 54155 50995 54466 51306 ne
rect 54466 51170 58365 51306
tri 58365 51170 58540 51345 sw
tri 58650 51170 58825 51345 ne
rect 58825 51170 60607 51345
rect 54466 50995 58540 51170
rect 50165 50732 54155 50995
rect 48110 50536 49878 50732
tri 49878 50536 50074 50732 sw
tri 50165 50536 50361 50732 ne
rect 50361 50684 54155 50732
tri 54155 50684 54466 50995 sw
tri 54466 50684 54777 50995 ne
rect 54777 50885 58540 50995
tri 58540 50885 58825 51170 sw
tri 58825 50885 59110 51170 ne
rect 59110 51084 60607 51170
tri 60607 51084 60891 51368 sw
tri 60891 51084 61175 51368 ne
rect 61175 51084 71000 51368
rect 59110 50885 60891 51084
rect 54777 50684 58825 50885
rect 50361 50536 54466 50684
rect 48110 50520 50074 50536
rect 45998 50360 47818 50520
rect 41645 50176 45705 50360
rect 28140 50070 32278 50176
rect 26022 49918 27850 50070
rect 23994 49677 25733 49918
rect 20400 49380 23697 49677
tri 23697 49380 23994 49677 sw
tri 23994 49380 24291 49677 ne
rect 24291 49629 25733 49677
tri 25733 49629 26022 49918 sw
tri 26022 49629 26311 49918 ne
rect 26311 49780 27850 49918
tri 27850 49780 28140 50070 sw
tri 28140 49780 28430 50070 ne
rect 28430 49882 32278 50070
tri 32278 49882 32572 50176 sw
tri 32572 49882 32866 50176 ne
rect 32866 49888 36816 50176
tri 36816 49888 37104 50176 sw
tri 37104 49888 37392 50176 ne
rect 37392 49888 41348 50176
rect 32866 49882 37104 49888
rect 28430 49780 32572 49882
rect 26311 49629 28140 49780
rect 24291 49380 26022 49629
rect 20400 49265 23994 49380
tri 23994 49265 24109 49380 sw
tri 24291 49265 24406 49380 ne
rect 24406 49340 26022 49380
tri 26022 49340 26311 49629 sw
tri 26311 49340 26600 49629 ne
rect 26600 49490 28140 49629
tri 28140 49490 28430 49780 sw
tri 28430 49490 28720 49780 ne
rect 28720 49588 32572 49780
tri 32572 49588 32866 49882 sw
tri 32866 49588 33160 49882 ne
rect 33160 49600 37104 49882
tri 37104 49600 37392 49888 sw
tri 37392 49600 37680 49888 ne
rect 37680 49879 41348 49888
tri 41348 49879 41645 50176 sw
tri 41645 49879 41942 50176 ne
rect 41942 50067 45705 50176
tri 45705 50067 45998 50360 sw
tri 45998 50067 46291 50360 ne
rect 46291 50228 47818 50360
tri 47818 50228 48110 50520 sw
tri 48110 50228 48402 50520 ne
rect 48402 50249 50074 50520
tri 50074 50249 50361 50536 sw
tri 50361 50249 50648 50536 ne
rect 50648 50373 54466 50536
tri 54466 50373 54777 50684 sw
tri 54777 50373 55088 50684 ne
rect 55088 50600 58825 50684
tri 58825 50600 59110 50885 sw
tri 59110 50600 59395 50885 ne
rect 59395 50800 60891 50885
tri 60891 50800 61175 51084 sw
tri 61175 50800 61459 51084 ne
rect 61459 50800 71000 51084
rect 59395 50600 61175 50800
tri 61175 50600 61375 50800 sw
rect 55088 50520 59110 50600
tri 59110 50520 59190 50600 sw
tri 59395 50520 59475 50600 ne
rect 59475 50520 71000 50600
rect 55088 50373 59190 50520
rect 50648 50249 54777 50373
rect 48402 50228 50361 50249
rect 46291 50067 48110 50228
rect 41942 49879 45998 50067
rect 37680 49600 41645 49879
rect 33160 49588 37392 49600
rect 28720 49490 32866 49588
rect 26600 49340 28430 49490
rect 24406 49265 26311 49340
rect 20400 48968 24109 49265
tri 24109 48968 24406 49265 sw
tri 24406 48968 24703 49265 ne
rect 24703 49051 26311 49265
tri 26311 49051 26600 49340 sw
tri 26600 49051 26889 49340 ne
rect 26889 49250 28430 49340
tri 28430 49250 28670 49490 sw
tri 28720 49250 28960 49490 ne
rect 28960 49294 32866 49490
tri 32866 49294 33160 49588 sw
tri 33160 49294 33454 49588 ne
rect 33454 49312 37392 49588
tri 37392 49312 37680 49600 sw
tri 37680 49312 37968 49600 ne
rect 37968 49582 41645 49600
tri 41645 49582 41942 49879 sw
tri 41942 49582 42239 49879 ne
rect 42239 49774 45998 49879
tri 45998 49774 46291 50067 sw
tri 46291 49774 46584 50067 ne
rect 46584 49936 48110 50067
tri 48110 49936 48402 50228 sw
tri 48402 49936 48694 50228 ne
rect 48694 49962 50361 50228
tri 50361 49962 50648 50249 sw
tri 50648 49962 50935 50249 ne
rect 50935 50062 54777 50249
tri 54777 50062 55088 50373 sw
tri 55088 50062 55399 50373 ne
rect 55399 50249 59190 50373
tri 59190 50249 59461 50520 sw
tri 59475 50249 59746 50520 ne
rect 59746 50249 71000 50520
rect 55399 50062 59461 50249
rect 50935 49962 55088 50062
rect 48694 49936 50648 49962
rect 46584 49774 48402 49936
rect 42239 49718 46291 49774
tri 46291 49718 46347 49774 sw
tri 46584 49718 46640 49774 ne
rect 46640 49718 48402 49774
rect 42239 49582 46347 49718
rect 37968 49312 41942 49582
rect 33454 49294 37680 49312
rect 28960 49250 33160 49294
rect 26889 49051 28670 49250
rect 24703 49049 26600 49051
tri 26600 49049 26602 49051 sw
tri 26889 49049 26891 49051 ne
rect 26891 49049 28670 49051
rect 24703 48968 26602 49049
rect 20400 48730 24406 48968
tri 20400 48648 20482 48730 ne
rect 20482 48671 24406 48730
tri 24406 48671 24703 48968 sw
tri 24703 48671 25000 48968 ne
rect 25000 48760 26602 48968
tri 26602 48760 26891 49049 sw
tri 26891 48760 27180 49049 ne
rect 27180 48960 28670 49049
tri 28670 48960 28960 49250 sw
tri 28960 48960 29250 49250 ne
rect 29250 49196 33160 49250
tri 33160 49196 33258 49294 sw
tri 33454 49196 33552 49294 ne
rect 33552 49196 37680 49294
rect 29250 48960 33258 49196
rect 27180 48760 28960 48960
rect 25000 48671 26891 48760
rect 20482 48648 24703 48671
tri 20200 48366 20482 48648 sw
tri 20482 48366 20764 48648 ne
rect 20764 48380 24703 48648
tri 24703 48380 24994 48671 sw
tri 25000 48380 25291 48671 ne
rect 25291 48669 26891 48671
tri 26891 48669 26982 48760 sw
tri 27180 48669 27271 48760 ne
rect 27271 48670 28960 48760
tri 28960 48670 29250 48960 sw
tri 29250 48670 29540 48960 ne
rect 29540 48902 33258 48960
tri 33258 48902 33552 49196 sw
tri 33552 48902 33846 49196 ne
rect 33846 49024 37680 49196
tri 37680 49024 37968 49312 sw
tri 37968 49024 38256 49312 ne
rect 38256 49285 41942 49312
tri 41942 49285 42239 49582 sw
tri 42239 49285 42536 49582 ne
rect 42536 49425 46347 49582
tri 46347 49425 46640 49718 sw
tri 46640 49425 46933 49718 ne
rect 46933 49644 48402 49718
tri 48402 49644 48694 49936 sw
tri 48694 49644 48986 49936 ne
rect 48986 49675 50648 49936
tri 50648 49675 50935 49962 sw
tri 50935 49675 51222 49962 ne
rect 51222 49784 55088 49962
tri 55088 49784 55366 50062 sw
tri 55399 49784 55677 50062 ne
rect 55677 49964 59461 50062
tri 59461 49964 59746 50249 sw
tri 59746 49964 60031 50249 ne
rect 60031 49964 71000 50249
rect 55677 49784 59746 49964
rect 51222 49675 55366 49784
rect 48986 49644 50935 49675
rect 46933 49504 48694 49644
tri 48694 49504 48834 49644 sw
tri 48986 49504 49126 49644 ne
rect 49126 49504 50935 49644
rect 46933 49425 48834 49504
rect 42536 49285 46640 49425
rect 38256 49271 42239 49285
tri 42239 49271 42253 49285 sw
tri 42536 49271 42550 49285 ne
rect 42550 49271 46640 49285
rect 38256 49024 42253 49271
rect 33846 48902 37968 49024
rect 29540 48670 33552 48902
rect 27271 48669 29250 48670
rect 25291 48380 26982 48669
tri 26982 48380 27271 48669 sw
tri 27271 48380 27560 48669 ne
rect 27560 48380 29250 48669
tri 29250 48380 29540 48670 sw
tri 29540 48380 29830 48670 ne
rect 29830 48608 33552 48670
tri 33552 48608 33846 48902 sw
tri 33846 48608 34140 48902 ne
rect 34140 48736 37968 48902
tri 37968 48736 38256 49024 sw
tri 38256 48736 38544 49024 ne
rect 38544 48974 42253 49024
tri 42253 48974 42550 49271 sw
tri 42550 48974 42847 49271 ne
rect 42847 49132 46640 49271
tri 46640 49132 46933 49425 sw
tri 46933 49132 47226 49425 ne
rect 47226 49212 48834 49425
tri 48834 49212 49126 49504 sw
tri 49126 49212 49418 49504 ne
rect 49418 49401 50935 49504
tri 50935 49401 51209 49675 sw
tri 51222 49401 51496 49675 ne
rect 51496 49473 55366 49675
tri 55366 49473 55677 49784 sw
tri 55677 49473 55988 49784 ne
rect 55988 49679 59746 49784
tri 59746 49679 60031 49964 sw
tri 60031 49679 60316 49964 ne
rect 60316 49679 71000 49964
rect 55988 49570 60031 49679
tri 60031 49570 60140 49679 sw
tri 60316 49570 60425 49679 ne
rect 60425 49570 71000 49679
rect 55988 49473 60140 49570
rect 51496 49401 55677 49473
rect 49418 49212 51209 49401
rect 47226 49132 49126 49212
rect 42847 48974 46933 49132
rect 38544 48736 42550 48974
rect 34140 48704 38256 48736
tri 38256 48704 38288 48736 sw
tri 38544 48704 38576 48736 ne
rect 38576 48704 42550 48736
rect 34140 48608 38288 48704
rect 29830 48380 33846 48608
rect 20764 48366 24994 48380
rect 17200 48084 20482 48366
tri 20482 48084 20764 48366 sw
tri 20764 48084 21046 48366 ne
rect 21046 48084 24994 48366
rect 17200 47802 20764 48084
tri 20764 47802 21046 48084 sw
tri 21046 47802 21328 48084 ne
rect 21328 48083 24994 48084
tri 24994 48083 25291 48380 sw
tri 25291 48083 25588 48380 ne
rect 25588 48091 27271 48380
tri 27271 48091 27560 48380 sw
tri 27560 48091 27849 48380 ne
rect 27849 48310 29540 48380
tri 29540 48310 29610 48380 sw
tri 29830 48310 29900 48380 ne
rect 29900 48314 33846 48380
tri 33846 48314 34140 48608 sw
tri 34140 48314 34434 48608 ne
rect 34434 48416 38288 48608
tri 38288 48416 38576 48704 sw
tri 38576 48416 38864 48704 ne
rect 38864 48677 42550 48704
tri 42550 48677 42847 48974 sw
tri 42847 48677 43144 48974 ne
rect 43144 48839 46933 48974
tri 46933 48839 47226 49132 sw
tri 47226 48839 47519 49132 ne
rect 47519 48920 49126 49132
tri 49126 48920 49418 49212 sw
tri 49418 48920 49710 49212 ne
rect 49710 49114 51209 49212
tri 51209 49114 51496 49401 sw
tri 51496 49114 51783 49401 ne
rect 51783 49162 55677 49401
tri 55677 49162 55988 49473 sw
tri 55988 49162 56299 49473 ne
rect 56299 49285 60140 49473
tri 60140 49285 60425 49570 sw
tri 60425 49285 60710 49570 ne
rect 60710 49285 71000 49570
rect 56299 49162 60425 49285
rect 51783 49114 55988 49162
rect 49710 48920 51496 49114
rect 47519 48839 49418 48920
rect 43144 48677 47226 48839
rect 38864 48416 42847 48677
rect 34434 48314 38576 48416
rect 29900 48310 34140 48314
rect 27849 48091 29610 48310
rect 25588 48083 27560 48091
rect 21328 48020 25291 48083
tri 25291 48020 25354 48083 sw
tri 25588 48020 25651 48083 ne
rect 25651 48020 27560 48083
rect 21328 47802 25354 48020
rect 17200 47754 21046 47802
tri 21046 47754 21094 47802 sw
tri 21328 47754 21376 47802 ne
rect 21376 47754 25354 47802
rect 17200 47472 21094 47754
tri 21094 47472 21376 47754 sw
tri 21376 47472 21658 47754 ne
rect 21658 47723 25354 47754
tri 25354 47723 25651 48020 sw
tri 25651 47723 25948 48020 ne
rect 25948 47802 27560 48020
tri 27560 47802 27849 48091 sw
tri 27849 47802 28138 48091 ne
rect 28138 48020 29610 48091
tri 29610 48020 29900 48310 sw
tri 29900 48020 30190 48310 ne
rect 30190 48020 34140 48310
tri 34140 48020 34434 48314 sw
tri 34434 48020 34728 48314 ne
rect 34728 48128 38576 48314
tri 38576 48128 38864 48416 sw
tri 38864 48128 39152 48416 ne
rect 39152 48380 42847 48416
tri 42847 48380 43144 48677 sw
tri 43144 48380 43441 48677 ne
rect 43441 48673 47226 48677
tri 47226 48673 47392 48839 sw
tri 47519 48673 47685 48839 ne
rect 47685 48832 49418 48839
tri 49418 48832 49506 48920 sw
tri 49710 48832 49798 48920 ne
rect 49798 48832 51496 48920
rect 47685 48673 49506 48832
rect 43441 48380 47392 48673
tri 47392 48380 47685 48673 sw
tri 47685 48380 47978 48673 ne
rect 47978 48540 49506 48673
tri 49506 48540 49798 48832 sw
tri 49798 48540 50090 48832 ne
rect 50090 48827 51496 48832
tri 51496 48827 51783 49114 sw
tri 51783 48827 52070 49114 ne
rect 52070 48851 55988 49114
tri 55988 48851 56299 49162 sw
tri 56299 48851 56610 49162 ne
rect 56610 49000 60425 49162
tri 60425 49000 60710 49285 sw
tri 60710 49200 60795 49285 ne
rect 60795 49200 71000 49285
rect 56610 48851 71000 49000
rect 52070 48827 56299 48851
rect 50090 48540 51783 48827
tri 51783 48540 52070 48827 sw
tri 52070 48540 52357 48827 ne
rect 52357 48540 56299 48827
tri 56299 48540 56610 48851 sw
tri 56610 48540 56921 48851 ne
rect 56921 48540 71000 48851
rect 47978 48380 49798 48540
rect 39152 48128 43144 48380
rect 34728 48020 38864 48128
rect 28138 47802 29900 48020
rect 25948 47723 27849 47802
rect 21658 47472 25651 47723
rect 17200 47404 21376 47472
tri 17200 47312 17292 47404 ne
rect 17292 47312 21376 47404
tri 17000 47020 17292 47312 sw
tri 17292 47020 17584 47312 ne
rect 17584 47190 21376 47312
tri 21376 47190 21658 47472 sw
tri 21658 47190 21940 47472 ne
rect 21940 47426 25651 47472
tri 25651 47426 25948 47723 sw
tri 25948 47426 26245 47723 ne
rect 26245 47513 27849 47723
tri 27849 47513 28138 47802 sw
tri 28138 47513 28427 47802 ne
rect 28427 47730 29900 47802
tri 29900 47730 30190 48020 sw
tri 30190 47730 30480 48020 ne
rect 30480 47730 34434 48020
rect 28427 47513 30190 47730
rect 26245 47426 28138 47513
rect 21940 47374 25948 47426
tri 25948 47374 26000 47426 sw
tri 26245 47374 26297 47426 ne
rect 26297 47374 28138 47426
rect 21940 47190 26000 47374
rect 17584 47020 21658 47190
rect 14000 46728 17292 47020
tri 17292 46728 17584 47020 sw
tri 17584 46728 17876 47020 ne
rect 17876 46908 21658 47020
tri 21658 46908 21940 47190 sw
tri 21940 46908 22222 47190 ne
rect 22222 47077 26000 47190
tri 26000 47077 26297 47374 sw
tri 26297 47077 26594 47374 ne
rect 26594 47358 28138 47374
tri 28138 47358 28293 47513 sw
tri 28427 47358 28582 47513 ne
rect 28582 47440 30190 47513
tri 30190 47440 30480 47730 sw
tri 30480 47440 30770 47730 ne
rect 30770 47726 34434 47730
tri 34434 47726 34728 48020 sw
tri 34728 47726 35022 48020 ne
rect 35022 47840 38864 48020
tri 38864 47840 39152 48128 sw
tri 39152 47840 39440 48128 ne
rect 39440 48083 43144 48128
tri 43144 48083 43441 48380 sw
tri 43441 48083 43738 48380 ne
rect 43738 48087 47685 48380
tri 47685 48087 47978 48380 sw
tri 47978 48087 48271 48380 ne
rect 48271 48248 49798 48380
tri 49798 48248 50090 48540 sw
tri 50090 48248 50382 48540 ne
rect 50382 48253 52070 48540
tri 52070 48253 52357 48540 sw
tri 52357 48253 52644 48540 ne
rect 52644 48253 56610 48540
rect 50382 48248 52357 48253
rect 48271 48087 50090 48248
rect 43738 48083 47978 48087
rect 39440 47840 43441 48083
rect 35022 47726 39152 47840
rect 30770 47440 34728 47726
rect 28582 47358 30480 47440
rect 26594 47077 28293 47358
rect 22222 46908 26297 47077
rect 17876 46728 21940 46908
rect 14000 46448 17584 46728
tri 17584 46448 17864 46728 sw
tri 17876 46448 18156 46728 ne
rect 18156 46626 21940 46728
tri 21940 46626 22222 46908 sw
tri 22222 46626 22504 46908 ne
rect 22504 46780 26297 46908
tri 26297 46780 26594 47077 sw
tri 26594 46780 26891 47077 ne
rect 26891 47069 28293 47077
tri 28293 47069 28582 47358 sw
tri 28582 47069 28871 47358 ne
rect 28871 47150 30480 47358
tri 30480 47150 30770 47440 sw
tri 30770 47150 31060 47440 ne
rect 31060 47432 34728 47440
tri 34728 47432 35022 47726 sw
tri 35022 47432 35316 47726 ne
rect 35316 47552 39152 47726
tri 39152 47552 39440 47840 sw
tri 39440 47552 39728 47840 ne
rect 39728 47786 43441 47840
tri 43441 47786 43738 48083 sw
tri 43738 47786 44035 48083 ne
rect 44035 47794 47978 48083
tri 47978 47794 48271 48087 sw
tri 48271 47794 48564 48087 ne
rect 48564 47956 50090 48087
tri 50090 47956 50382 48248 sw
tri 50382 47956 50674 48248 ne
rect 50674 47966 52357 48248
tri 52357 47966 52644 48253 sw
tri 52644 47966 52931 48253 ne
rect 52931 48229 56610 48253
tri 56610 48229 56921 48540 sw
tri 56921 48229 57232 48540 ne
rect 57232 48229 71000 48540
rect 52931 47966 56921 48229
rect 50674 47956 52644 47966
rect 48564 47794 50382 47956
rect 44035 47786 48271 47794
rect 39728 47552 43738 47786
rect 35316 47432 39440 47552
rect 31060 47150 35022 47432
rect 28871 47069 30770 47150
rect 26891 46780 28582 47069
tri 28582 46780 28871 47069 sw
tri 28871 46780 29160 47069 ne
rect 29160 46980 30770 47069
tri 30770 46980 30940 47150 sw
tri 31060 46980 31230 47150 ne
rect 31230 47138 35022 47150
tri 35022 47138 35316 47432 sw
tri 35316 47138 35610 47432 ne
rect 35610 47264 39440 47432
tri 39440 47264 39728 47552 sw
tri 39728 47264 40016 47552 ne
rect 40016 47489 43738 47552
tri 43738 47489 44035 47786 sw
tri 44035 47489 44332 47786 ne
rect 44332 47526 48271 47786
tri 48271 47526 48539 47794 sw
tri 48564 47526 48832 47794 ne
rect 48832 47664 50382 47794
tri 50382 47664 50674 47956 sw
tri 50674 47664 50966 47956 ne
rect 50966 47914 52644 47956
tri 52644 47914 52696 47966 sw
tri 52931 47914 52983 47966 ne
rect 52983 47918 56921 47966
tri 56921 47918 57232 48229 sw
tri 57232 47918 57543 48229 ne
rect 57543 47918 71000 48229
rect 52983 47914 57232 47918
rect 50966 47664 52696 47914
rect 48832 47526 50674 47664
rect 44332 47489 48539 47526
rect 40016 47264 44035 47489
rect 35610 47138 39728 47264
rect 31230 46988 35316 47138
tri 35316 46988 35466 47138 sw
tri 35610 46988 35760 47138 ne
rect 35760 46988 39728 47138
rect 31230 46980 35466 46988
rect 29160 46780 30940 46980
rect 22504 46626 26594 46780
rect 18156 46448 22222 46626
rect 14000 46156 17864 46448
tri 17864 46156 18156 46448 sw
tri 18156 46156 18448 46448 ne
rect 18448 46344 22222 46448
tri 22222 46344 22504 46626 sw
tri 22504 46344 22786 46626 ne
rect 22786 46483 26594 46626
tri 26594 46483 26891 46780 sw
tri 26891 46483 27188 46780 ne
rect 27188 46689 28871 46780
tri 28871 46689 28962 46780 sw
tri 29160 46689 29251 46780 ne
rect 29251 46690 30940 46780
tri 30940 46690 31230 46980 sw
tri 31230 46690 31520 46980 ne
rect 31520 46694 35466 46980
tri 35466 46694 35760 46988 sw
tri 35760 46694 36054 46988 ne
rect 36054 46976 39728 46988
tri 39728 46976 40016 47264 sw
tri 40016 46976 40304 47264 ne
rect 40304 47192 44035 47264
tri 44035 47192 44332 47489 sw
tri 44332 47192 44629 47489 ne
rect 44629 47233 48539 47489
tri 48539 47233 48832 47526 sw
tri 48832 47233 49125 47526 ne
rect 49125 47524 50674 47526
tri 50674 47524 50814 47664 sw
tri 50966 47524 51106 47664 ne
rect 51106 47627 52696 47664
tri 52696 47627 52983 47914 sw
tri 52983 47627 53270 47914 ne
rect 53270 47675 57232 47914
tri 57232 47675 57475 47918 sw
tri 57543 47675 57786 47918 ne
rect 57786 47675 71000 47918
rect 53270 47627 57475 47675
rect 51106 47524 52983 47627
rect 49125 47233 50814 47524
rect 44629 47192 48832 47233
rect 40304 47120 44332 47192
tri 44332 47120 44404 47192 sw
tri 44629 47120 44701 47192 ne
rect 44701 47120 48832 47192
rect 40304 46976 44404 47120
rect 36054 46694 40016 46976
rect 31520 46690 35760 46694
rect 29251 46689 31230 46690
rect 27188 46483 28962 46689
rect 22786 46400 26891 46483
tri 26891 46400 26974 46483 sw
tri 27188 46400 27271 46483 ne
rect 27271 46400 28962 46483
tri 28962 46400 29251 46689 sw
tri 29251 46400 29540 46689 ne
rect 29540 46400 31230 46689
tri 31230 46400 31520 46690 sw
tri 31520 46400 31810 46690 ne
rect 31810 46400 35760 46690
tri 35760 46400 36054 46694 sw
tri 36054 46400 36348 46694 ne
rect 36348 46688 40016 46694
tri 40016 46688 40304 46976 sw
tri 40304 46688 40592 46976 ne
rect 40592 46823 44404 46976
tri 44404 46823 44701 47120 sw
tri 44701 46823 44998 47120 ne
rect 44998 46940 48832 47120
tri 48832 46940 49125 47233 sw
tri 49125 46940 49418 47233 ne
rect 49418 47232 50814 47233
tri 50814 47232 51106 47524 sw
tri 51106 47232 51398 47524 ne
rect 51398 47340 52983 47524
tri 52983 47340 53270 47627 sw
tri 53270 47340 53557 47627 ne
rect 53557 47364 57475 47627
tri 57475 47364 57786 47675 sw
tri 57786 47364 58097 47675 ne
rect 58097 47364 71000 47675
rect 53557 47340 57786 47364
rect 51398 47232 53270 47340
rect 49418 46940 51106 47232
tri 51106 46940 51398 47232 sw
tri 51398 46940 51690 47232 ne
rect 51690 47053 53270 47232
tri 53270 47053 53557 47340 sw
tri 53557 47053 53844 47340 ne
rect 53844 47053 57786 47340
tri 57786 47053 58097 47364 sw
tri 58097 47053 58408 47364 ne
rect 58408 47053 71000 47364
rect 51690 46940 53557 47053
rect 44998 46823 49125 46940
rect 40592 46688 44701 46823
rect 36348 46400 40304 46688
tri 40304 46400 40592 46688 sw
tri 40592 46400 40880 46688 ne
rect 40880 46526 44701 46688
tri 44701 46526 44998 46823 sw
tri 44998 46526 45295 46823 ne
rect 45295 46647 49125 46823
tri 49125 46647 49418 46940 sw
tri 49418 46647 49711 46940 ne
rect 49711 46852 51398 46940
tri 51398 46852 51486 46940 sw
tri 51690 46852 51778 46940 ne
rect 51778 46852 53557 46940
rect 49711 46647 51486 46852
rect 45295 46526 49418 46647
rect 40880 46400 44998 46526
rect 22786 46344 26974 46400
rect 18448 46156 22504 46344
rect 14000 46068 18156 46156
tri 14000 43708 16360 46068 ne
rect 16360 45864 18156 46068
tri 18156 45864 18448 46156 sw
tri 18448 45864 18740 46156 ne
rect 18740 46146 22504 46156
tri 22504 46146 22702 46344 sw
tri 22786 46146 22984 46344 ne
rect 22984 46161 26974 46344
tri 26974 46161 27213 46400 sw
tri 27271 46161 27510 46400 ne
rect 27510 46161 29251 46400
rect 22984 46146 27213 46161
rect 18740 45864 22702 46146
tri 22702 45864 22984 46146 sw
tri 22984 45864 23266 46146 ne
rect 23266 45864 27213 46146
tri 27213 45864 27510 46161 sw
tri 27510 45864 27807 46161 ne
rect 27807 46111 29251 46161
tri 29251 46111 29540 46400 sw
tri 29540 46111 29829 46400 ne
rect 29829 46111 31520 46400
rect 27807 45864 29540 46111
rect 16360 45572 18448 45864
tri 18448 45572 18740 45864 sw
tri 18740 45572 19032 45864 ne
rect 19032 45582 22984 45864
tri 22984 45582 23266 45864 sw
tri 23266 45582 23548 45864 ne
rect 23548 45582 27510 45864
rect 19032 45572 23266 45582
rect 16360 45280 18740 45572
tri 18740 45280 19032 45572 sw
tri 19032 45280 19324 45572 ne
rect 19324 45300 23266 45572
tri 23266 45300 23548 45582 sw
tri 23548 45300 23830 45582 ne
rect 23830 45567 27510 45582
tri 27510 45567 27807 45864 sw
tri 27807 45567 28104 45864 ne
rect 28104 45822 29540 45864
tri 29540 45822 29829 46111 sw
tri 29829 45822 30118 46111 ne
rect 30118 46110 31520 46111
tri 31520 46110 31810 46400 sw
tri 31810 46110 32100 46400 ne
rect 32100 46110 36054 46400
rect 30118 45822 31810 46110
rect 28104 45567 29829 45822
rect 23830 45300 27807 45567
rect 19324 45280 23548 45300
rect 16360 44988 19032 45280
tri 19032 44988 19324 45280 sw
tri 19324 44988 19616 45280 ne
rect 19616 45018 23548 45280
tri 23548 45018 23830 45300 sw
tri 23830 45018 24112 45300 ne
rect 24112 45270 27807 45300
tri 27807 45270 28104 45567 sw
tri 28104 45270 28401 45567 ne
rect 28401 45533 29829 45567
tri 29829 45533 30118 45822 sw
tri 30118 45533 30407 45822 ne
rect 30407 45820 31810 45822
tri 31810 45820 32100 46110 sw
tri 32100 45820 32390 46110 ne
rect 32390 46106 36054 46110
tri 36054 46106 36348 46400 sw
tri 36348 46106 36642 46400 ne
rect 36642 46220 40592 46400
tri 40592 46220 40772 46400 sw
tri 40880 46220 41060 46400 ne
rect 41060 46229 44998 46400
tri 44998 46229 45295 46526 sw
tri 45295 46229 45592 46526 ne
rect 45592 46400 49418 46526
tri 49418 46400 49665 46647 sw
tri 49711 46400 49958 46647 ne
rect 49958 46560 51486 46647
tri 51486 46560 51778 46852 sw
tri 51778 46560 52070 46852 ne
rect 52070 46766 53557 46852
tri 53557 46766 53844 47053 sw
tri 53844 46766 54131 47053 ne
rect 54131 46766 58097 47053
rect 52070 46560 53844 46766
rect 49958 46400 51778 46560
rect 45592 46229 49665 46400
rect 41060 46220 45295 46229
rect 36642 46106 40772 46220
rect 32390 45820 36348 46106
rect 30407 45533 32100 45820
rect 28401 45378 30118 45533
tri 30118 45378 30273 45533 sw
tri 30407 45378 30562 45533 ne
rect 30562 45530 32100 45533
tri 32100 45530 32390 45820 sw
tri 32390 45530 32680 45820 ne
rect 32680 45812 36348 45820
tri 36348 45812 36642 46106 sw
tri 36642 45812 36936 46106 ne
rect 36936 45932 40772 46106
tri 40772 45932 41060 46220 sw
tri 41060 45932 41348 46220 ne
rect 41348 45932 45295 46220
tri 45295 45932 45592 46229 sw
tri 45592 45932 45889 46229 ne
rect 45889 46107 49665 46229
tri 49665 46107 49958 46400 sw
tri 49958 46107 50251 46400 ne
rect 50251 46268 51778 46400
tri 51778 46268 52070 46560 sw
tri 52070 46268 52362 46560 ne
rect 52362 46479 53844 46560
tri 53844 46479 54131 46766 sw
tri 54131 46479 54418 46766 ne
rect 54418 46742 58097 46766
tri 58097 46742 58408 47053 sw
tri 58408 46742 58719 47053 ne
rect 58719 46742 71000 47053
rect 54418 46479 58408 46742
rect 52362 46287 54131 46479
tri 54131 46287 54323 46479 sw
tri 54418 46287 54610 46479 ne
rect 54610 46431 58408 46479
tri 58408 46431 58719 46742 sw
tri 58719 46431 59030 46742 ne
rect 59030 46431 71000 46742
rect 54610 46421 58719 46431
tri 58719 46421 58729 46431 sw
tri 59030 46421 59040 46431 ne
rect 59040 46421 71000 46431
rect 54610 46287 58729 46421
rect 52362 46268 54323 46287
rect 50251 46107 52070 46268
rect 45889 45932 49958 46107
rect 36936 45812 41060 45932
rect 32680 45530 36642 45812
rect 30562 45378 32390 45530
rect 28401 45270 30273 45378
rect 24112 45018 28104 45270
rect 19616 44988 23830 45018
rect 16360 44876 19324 44988
tri 19324 44876 19436 44988 sw
tri 19616 44876 19728 44988 ne
rect 19728 44876 23830 44988
rect 16360 44584 19436 44876
tri 19436 44584 19728 44876 sw
tri 19728 44584 20020 44876 ne
rect 20020 44736 23830 44876
tri 23830 44736 24112 45018 sw
tri 24112 44736 24394 45018 ne
rect 24394 45014 28104 45018
tri 28104 45014 28360 45270 sw
tri 28401 45014 28657 45270 ne
rect 28657 45089 30273 45270
tri 30273 45089 30562 45378 sw
tri 30562 45089 30851 45378 ne
rect 30851 45290 32390 45378
tri 32390 45290 32630 45530 sw
tri 32680 45290 32920 45530 ne
rect 32920 45518 36642 45530
tri 36642 45518 36936 45812 sw
tri 36936 45518 37230 45812 ne
rect 37230 45644 41060 45812
tri 41060 45644 41348 45932 sw
tri 41348 45644 41636 45932 ne
rect 41636 45644 45592 45932
rect 37230 45518 41348 45644
rect 32920 45290 36936 45518
rect 30851 45089 32630 45290
rect 28657 45014 30562 45089
rect 24394 44736 28360 45014
rect 20020 44584 24112 44736
rect 16360 44292 19728 44584
tri 19728 44292 20020 44584 sw
tri 20020 44292 20312 44584 ne
rect 20312 44454 24112 44584
tri 24112 44454 24394 44736 sw
tri 24394 44454 24676 44736 ne
rect 24676 44717 28360 44736
tri 28360 44717 28657 45014 sw
tri 28657 44717 28954 45014 ne
rect 28954 44800 30562 45014
tri 30562 44800 30851 45089 sw
tri 30851 44800 31140 45089 ne
rect 31140 45000 32630 45089
tri 32630 45000 32920 45290 sw
tri 32920 45000 33210 45290 ne
rect 33210 45224 36936 45290
tri 36936 45224 37230 45518 sw
tri 37230 45224 37524 45518 ne
rect 37524 45356 41348 45518
tri 41348 45356 41636 45644 sw
tri 41636 45356 41924 45644 ne
rect 41924 45635 45592 45644
tri 45592 45635 45889 45932 sw
tri 45889 45635 46186 45932 ne
rect 46186 45814 49958 45932
tri 49958 45814 50251 46107 sw
tri 50251 45814 50544 46107 ne
rect 50544 45976 52070 46107
tri 52070 45976 52362 46268 sw
tri 52362 45976 52654 46268 ne
rect 52654 46000 54323 46268
tri 54323 46000 54610 46287 sw
tri 54610 46000 54897 46287 ne
rect 54897 46110 58729 46287
tri 58729 46110 59040 46421 sw
tri 59040 46110 59351 46421 ne
rect 59351 46110 71000 46421
rect 54897 46000 59040 46110
rect 52654 45976 54610 46000
rect 50544 45814 52362 45976
rect 46186 45767 50251 45814
tri 50251 45767 50298 45814 sw
tri 50544 45767 50591 45814 ne
rect 50591 45767 52362 45814
rect 46186 45635 50298 45767
rect 41924 45356 45889 45635
rect 37524 45224 41636 45356
rect 33210 45000 37230 45224
rect 31140 44800 32920 45000
rect 28954 44717 30851 44800
rect 24676 44454 28657 44717
rect 20312 44356 24394 44454
tri 24394 44356 24492 44454 sw
tri 24676 44356 24774 44454 ne
rect 24774 44420 28657 44454
tri 28657 44420 28954 44717 sw
tri 28954 44420 29251 44717 ne
rect 29251 44709 30851 44717
tri 30851 44709 30942 44800 sw
tri 31140 44709 31231 44800 ne
rect 31231 44710 32920 44800
tri 32920 44710 33210 45000 sw
tri 33210 44710 33500 45000 ne
rect 33500 44952 37230 45000
tri 37230 44952 37502 45224 sw
tri 37524 44952 37796 45224 ne
rect 37796 45068 41636 45224
tri 41636 45068 41924 45356 sw
tri 41924 45068 42212 45356 ne
rect 42212 45338 45889 45356
tri 45889 45338 46186 45635 sw
tri 46186 45338 46483 45635 ne
rect 46483 45474 50298 45635
tri 50298 45474 50591 45767 sw
tri 50591 45474 50884 45767 ne
rect 50884 45684 52362 45767
tri 52362 45684 52654 45976 sw
tri 52654 45684 52946 45976 ne
rect 52946 45713 54610 45976
tri 54610 45713 54897 46000 sw
tri 54897 45713 55184 46000 ne
rect 55184 45799 59040 46000
tri 59040 45799 59351 46110 sw
tri 59351 46000 59461 46110 ne
rect 59461 46000 71000 46110
rect 55184 45739 71000 45799
rect 55184 45713 70613 45739
rect 52946 45684 54897 45713
rect 50884 45544 52654 45684
tri 52654 45544 52794 45684 sw
tri 52946 45544 53086 45684 ne
rect 53086 45544 54897 45684
rect 50884 45474 52794 45544
rect 46483 45338 50591 45474
rect 42212 45068 46186 45338
rect 37796 44952 41924 45068
rect 33500 44710 37502 44952
rect 31231 44709 33210 44710
rect 29251 44420 30942 44709
tri 30942 44420 31231 44709 sw
tri 31231 44420 31520 44709 ne
rect 31520 44420 33210 44709
tri 33210 44420 33500 44710 sw
tri 33500 44420 33790 44710 ne
rect 33790 44658 37502 44710
tri 37502 44658 37796 44952 sw
tri 37796 44658 38090 44952 ne
rect 38090 44780 41924 44952
tri 41924 44780 42212 45068 sw
tri 42212 44780 42500 45068 ne
rect 42500 45041 46186 45068
tri 46186 45041 46483 45338 sw
tri 46483 45041 46780 45338 ne
rect 46780 45181 50591 45338
tri 50591 45181 50884 45474 sw
tri 50884 45181 51177 45474 ne
rect 51177 45252 52794 45474
tri 52794 45252 53086 45544 sw
tri 53086 45252 53378 45544 ne
rect 53378 45426 54897 45544
tri 54897 45426 55184 45713 sw
tri 55184 45426 55471 45713 ne
rect 55471 45426 70613 45713
rect 53378 45252 55184 45426
rect 51177 45181 53086 45252
rect 46780 45041 50884 45181
rect 42500 45014 46483 45041
tri 46483 45014 46510 45041 sw
tri 46780 45014 46807 45041 ne
rect 46807 45014 50884 45041
rect 42500 44780 46510 45014
rect 38090 44658 42212 44780
rect 33790 44420 37796 44658
rect 24774 44356 28954 44420
rect 20312 44292 24492 44356
rect 16360 44000 20020 44292
tri 20020 44000 20312 44292 sw
tri 20312 44000 20604 44292 ne
rect 20604 44074 24492 44292
tri 24492 44074 24774 44356 sw
tri 24774 44074 25056 44356 ne
rect 25056 44123 28954 44356
tri 28954 44123 29251 44420 sw
tri 29251 44123 29548 44420 ne
rect 29548 44131 31231 44420
tri 31231 44131 31520 44420 sw
tri 31520 44131 31809 44420 ne
rect 31809 44131 33500 44420
rect 29548 44123 31520 44131
rect 25056 44074 29251 44123
rect 20604 44000 24774 44074
rect 16360 43708 20312 44000
tri 20312 43708 20604 44000 sw
tri 20604 43708 20896 44000 ne
rect 20896 43792 24774 44000
tri 24774 43792 25056 44074 sw
tri 25056 43792 25338 44074 ne
rect 25338 44073 29251 44074
tri 29251 44073 29301 44123 sw
tri 29548 44073 29598 44123 ne
rect 29598 44073 31520 44123
rect 25338 43792 29301 44073
rect 20896 43708 25056 43792
tri 16360 39464 20604 43708 ne
tri 20604 43416 20896 43708 sw
tri 20896 43416 21188 43708 ne
rect 21188 43510 25056 43708
tri 25056 43510 25338 43792 sw
tri 25338 43510 25620 43792 ne
rect 25620 43776 29301 43792
tri 29301 43776 29598 44073 sw
tri 29598 43776 29895 44073 ne
rect 29895 43842 31520 44073
tri 31520 43842 31809 44131 sw
tri 31809 43842 32098 44131 ne
rect 32098 44130 33500 44131
tri 33500 44130 33790 44420 sw
tri 33790 44130 34080 44420 ne
rect 34080 44364 37796 44420
tri 37796 44364 38090 44658 sw
tri 38090 44364 38384 44658 ne
rect 38384 44492 42212 44658
tri 42212 44492 42500 44780 sw
tri 42500 44492 42788 44780 ne
rect 42788 44717 46510 44780
tri 46510 44717 46807 45014 sw
tri 46807 44717 47104 45014 ne
rect 47104 44888 50884 45014
tri 50884 44888 51177 45181 sw
tri 51177 44888 51470 45181 ne
rect 51470 44960 53086 45181
tri 53086 44960 53378 45252 sw
tri 53378 44960 53670 45252 ne
rect 53670 45154 55184 45252
tri 55184 45154 55456 45426 sw
tri 55471 45154 55743 45426 ne
rect 55743 45154 70613 45426
rect 53670 44960 55456 45154
rect 51470 44888 53378 44960
rect 47104 44717 51177 44888
rect 42788 44492 46807 44717
rect 38384 44460 42500 44492
tri 42500 44460 42532 44492 sw
tri 42788 44460 42820 44492 ne
rect 42820 44460 46807 44492
rect 38384 44364 42532 44460
rect 34080 44130 38090 44364
rect 32098 44066 33790 44130
tri 33790 44066 33854 44130 sw
tri 34080 44066 34144 44130 ne
rect 34144 44070 38090 44130
tri 38090 44070 38384 44364 sw
tri 38384 44070 38678 44364 ne
rect 38678 44172 42532 44364
tri 42532 44172 42820 44460 sw
tri 42820 44172 43108 44460 ne
rect 43108 44420 46807 44460
tri 46807 44420 47104 44717 sw
tri 47104 44420 47401 44717 ne
rect 47401 44595 51177 44717
tri 51177 44595 51470 44888 sw
tri 51470 44595 51763 44888 ne
rect 51763 44872 53378 44888
tri 53378 44872 53466 44960 sw
tri 53670 44872 53758 44960 ne
rect 53758 44872 55456 44960
rect 51763 44595 53466 44872
rect 47401 44420 51470 44595
tri 51470 44420 51645 44595 sw
tri 51763 44420 51938 44595 ne
rect 51938 44580 53466 44595
tri 53466 44580 53758 44872 sw
tri 53758 44580 54050 44872 ne
rect 54050 44867 55456 44872
tri 55456 44867 55743 45154 sw
tri 55743 44867 56030 45154 ne
rect 56030 44867 70613 45154
rect 54050 44580 55743 44867
tri 55743 44580 56030 44867 sw
tri 56030 44580 56317 44867 ne
rect 56317 44580 70613 44867
rect 51938 44420 53758 44580
rect 43108 44172 47104 44420
rect 38678 44070 42820 44172
rect 34144 44066 38384 44070
rect 32098 43842 33854 44066
rect 29895 43776 31809 43842
rect 25620 43510 29598 43776
rect 21188 43416 25338 43510
rect 20604 43124 20896 43416
tri 20896 43124 21188 43416 sw
tri 21188 43124 21480 43416 ne
rect 21480 43228 25338 43416
tri 25338 43228 25620 43510 sw
tri 25620 43228 25902 43510 ne
rect 25902 43479 29598 43510
tri 29598 43479 29895 43776 sw
tri 29895 43479 30192 43776 ne
rect 30192 43553 31809 43776
tri 31809 43553 32098 43842 sw
tri 32098 43553 32387 43842 ne
rect 32387 43776 33854 43842
tri 33854 43776 34144 44066 sw
tri 34144 43776 34434 44066 ne
rect 34434 43776 38384 44066
tri 38384 43776 38678 44070 sw
tri 38678 43776 38972 44070 ne
rect 38972 43884 42820 44070
tri 42820 43884 43108 44172 sw
tri 43108 43884 43396 44172 ne
rect 43396 44123 47104 44172
tri 47104 44123 47401 44420 sw
tri 47401 44123 47698 44420 ne
rect 47698 44127 51645 44420
tri 51645 44127 51938 44420 sw
tri 51938 44127 52231 44420 ne
rect 52231 44288 53758 44420
tri 53758 44288 54050 44580 sw
tri 54050 44288 54342 44580 ne
rect 54342 44293 56030 44580
tri 56030 44293 56317 44580 sw
tri 56317 44293 56604 44580 ne
rect 56604 44293 70613 44580
rect 54342 44288 56317 44293
rect 52231 44127 54050 44288
rect 47698 44123 51938 44127
rect 43396 43884 47401 44123
rect 38972 43776 43108 43884
rect 32387 43553 34144 43776
rect 30192 43479 32098 43553
rect 25902 43228 29895 43479
rect 21480 43124 25620 43228
rect 20604 42832 21188 43124
tri 21188 42832 21480 43124 sw
tri 21480 42832 21772 43124 ne
rect 21772 42946 25620 43124
tri 25620 42946 25902 43228 sw
tri 25902 42946 26184 43228 ne
rect 26184 43182 29895 43228
tri 29895 43182 30192 43479 sw
tri 30192 43182 30489 43479 ne
rect 30489 43398 32098 43479
tri 32098 43398 32253 43553 sw
tri 32387 43398 32542 43553 ne
rect 32542 43486 34144 43553
tri 34144 43486 34434 43776 sw
tri 34434 43486 34724 43776 ne
rect 34724 43486 38678 43776
rect 32542 43398 34434 43486
rect 30489 43182 32253 43398
rect 26184 43117 30192 43182
tri 30192 43117 30257 43182 sw
tri 30489 43117 30554 43182 ne
rect 30554 43117 32253 43182
rect 26184 42946 30257 43117
rect 21772 42832 25902 42946
rect 20604 42540 21480 42832
tri 21480 42540 21772 42832 sw
tri 21772 42540 22064 42832 ne
rect 22064 42664 25902 42832
tri 25902 42664 26184 42946 sw
tri 26184 42664 26466 42946 ne
rect 26466 42820 30257 42946
tri 30257 42820 30554 43117 sw
tri 30554 42820 30851 43117 ne
rect 30851 43109 32253 43117
tri 32253 43109 32542 43398 sw
tri 32542 43109 32831 43398 ne
rect 32831 43196 34434 43398
tri 34434 43196 34724 43486 sw
tri 34724 43196 35014 43486 ne
rect 35014 43482 38678 43486
tri 38678 43482 38972 43776 sw
tri 38972 43482 39266 43776 ne
rect 39266 43596 43108 43776
tri 43108 43596 43396 43884 sw
tri 43396 43596 43684 43884 ne
rect 43684 43826 47401 43884
tri 47401 43826 47698 44123 sw
tri 47698 43826 47995 44123 ne
rect 47995 43834 51938 44123
tri 51938 43834 52231 44127 sw
tri 52231 43834 52524 44127 ne
rect 52524 43996 54050 44127
tri 54050 43996 54342 44288 sw
tri 54342 43996 54634 44288 ne
rect 54634 44006 56317 44288
tri 56317 44006 56604 44293 sw
tri 56604 44006 56891 44293 ne
rect 56891 44006 70613 44293
rect 54634 43996 56604 44006
rect 52524 43834 54342 43996
rect 47995 43826 52231 43834
rect 43684 43596 47698 43826
rect 39266 43482 43396 43596
rect 35014 43196 38972 43482
rect 32831 43109 34724 43196
rect 30851 42820 32542 43109
tri 32542 42820 32831 43109 sw
tri 32831 42820 33120 43109 ne
rect 33120 43020 34724 43109
tri 34724 43020 34900 43196 sw
tri 35014 43020 35190 43196 ne
rect 35190 43188 38972 43196
tri 38972 43188 39266 43482 sw
tri 39266 43188 39560 43482 ne
rect 39560 43308 43396 43482
tri 43396 43308 43684 43596 sw
tri 43684 43308 43972 43596 ne
rect 43972 43529 47698 43596
tri 47698 43529 47995 43826 sw
tri 47995 43529 48292 43826 ne
rect 48292 43566 52231 43826
tri 52231 43566 52499 43834 sw
tri 52524 43566 52792 43834 ne
rect 52792 43704 54342 43834
tri 54342 43704 54634 43996 sw
tri 54634 43704 54926 43996 ne
rect 54926 43719 56604 43996
tri 56604 43719 56891 44006 sw
tri 56891 43719 57178 44006 ne
rect 57178 43719 70613 44006
rect 54926 43704 56891 43719
rect 52792 43566 54634 43704
rect 48292 43529 52499 43566
rect 43972 43308 47995 43529
rect 39560 43188 43684 43308
rect 35190 43028 39266 43188
tri 39266 43028 39426 43188 sw
tri 39560 43028 39720 43188 ne
rect 39720 43028 43684 43188
rect 35190 43020 39426 43028
rect 33120 42820 34900 43020
rect 26466 42664 30554 42820
rect 22064 42540 26184 42664
rect 20604 42496 21772 42540
tri 21772 42496 21816 42540 sw
tri 22064 42496 22108 42540 ne
rect 22108 42496 26184 42540
rect 20604 42204 21816 42496
tri 21816 42204 22108 42496 sw
tri 22108 42204 22400 42496 ne
rect 22400 42382 26184 42496
tri 26184 42382 26466 42664 sw
tri 26466 42382 26748 42664 ne
rect 26748 42523 30554 42664
tri 30554 42523 30851 42820 sw
tri 30851 42523 31148 42820 ne
rect 31148 42729 32831 42820
tri 32831 42729 32922 42820 sw
tri 33120 42729 33211 42820 ne
rect 33211 42730 34900 42820
tri 34900 42730 35190 43020 sw
tri 35190 42730 35480 43020 ne
rect 35480 42734 39426 43020
tri 39426 42734 39720 43028 sw
tri 39720 42734 40014 43028 ne
rect 40014 43020 43684 43028
tri 43684 43020 43972 43308 sw
tri 43972 43020 44260 43308 ne
rect 44260 43232 47995 43308
tri 47995 43232 48292 43529 sw
tri 48292 43232 48589 43529 ne
rect 48589 43273 52499 43529
tri 52499 43273 52792 43566 sw
tri 52792 43273 53085 43566 ne
rect 53085 43564 54634 43566
tri 54634 43564 54774 43704 sw
tri 54926 43564 55066 43704 ne
rect 55066 43661 56891 43704
tri 56891 43661 56949 43719 sw
tri 57178 43661 57236 43719 ne
rect 57236 43661 70613 43719
rect 55066 43564 56949 43661
rect 53085 43273 54774 43564
rect 48589 43232 52792 43273
rect 44260 43173 48292 43232
tri 48292 43173 48351 43232 sw
tri 48589 43173 48648 43232 ne
rect 48648 43173 52792 43232
rect 44260 43020 48351 43173
rect 40014 42734 43972 43020
rect 35480 42730 39720 42734
rect 33211 42729 35190 42730
rect 31148 42523 32922 42729
rect 26748 42440 30851 42523
tri 30851 42440 30934 42523 sw
tri 31148 42440 31231 42523 ne
rect 31231 42440 32922 42523
tri 32922 42440 33211 42729 sw
tri 33211 42440 33500 42729 ne
rect 33500 42440 35190 42729
tri 35190 42440 35480 42730 sw
tri 35480 42440 35770 42730 ne
rect 35770 42440 39720 42730
tri 39720 42440 40014 42734 sw
tri 40014 42440 40308 42734 ne
rect 40308 42732 43972 42734
tri 43972 42732 44260 43020 sw
tri 44260 42732 44548 43020 ne
rect 44548 42876 48351 43020
tri 48351 42876 48648 43173 sw
tri 48648 42876 48945 43173 ne
rect 48945 42980 52792 43173
tri 52792 42980 53085 43273 sw
tri 53085 42980 53378 43273 ne
rect 53378 43272 54774 43273
tri 54774 43272 55066 43564 sw
tri 55066 43272 55358 43564 ne
rect 55358 43374 56949 43564
tri 56949 43374 57236 43661 sw
tri 57236 43374 57523 43661 ne
rect 57523 43374 70613 43661
rect 55358 43272 57236 43374
rect 53378 42980 55066 43272
tri 55066 42980 55358 43272 sw
tri 55358 42980 55650 43272 ne
rect 55650 43087 57236 43272
tri 57236 43087 57523 43374 sw
tri 57523 43087 57810 43374 ne
rect 57810 43087 70613 43374
rect 55650 42980 57523 43087
rect 48945 42876 53085 42980
rect 44548 42732 48648 42876
rect 40308 42444 44260 42732
tri 44260 42444 44548 42732 sw
tri 44548 42444 44836 42732 ne
rect 44836 42579 48648 42732
tri 48648 42579 48945 42876 sw
tri 48945 42579 49242 42876 ne
rect 49242 42687 53085 42876
tri 53085 42687 53378 42980 sw
tri 53378 42687 53671 42980 ne
rect 53671 42800 55358 42980
tri 55358 42800 55538 42980 sw
tri 55650 42800 55830 42980 ne
rect 55830 42800 57523 42980
tri 57523 42800 57810 43087 sw
tri 57810 42800 58097 43087 ne
rect 58097 42875 70613 43087
rect 70669 42875 71000 45739
rect 58097 42800 71000 42875
rect 53671 42687 55538 42800
rect 49242 42579 53378 42687
rect 44836 42444 48945 42579
rect 40308 42440 44548 42444
rect 26748 42382 30934 42440
rect 22400 42204 26466 42382
rect 20604 41912 22108 42204
tri 22108 41912 22400 42204 sw
tri 22400 41912 22692 42204 ne
rect 22692 42100 26466 42204
tri 26466 42100 26748 42382 sw
tri 26748 42100 27030 42382 ne
rect 27030 42143 30934 42382
tri 30934 42143 31231 42440 sw
tri 31231 42143 31528 42440 ne
rect 31528 42151 33211 42440
tri 33211 42151 33500 42440 sw
tri 33500 42151 33789 42440 ne
rect 33789 42151 35480 42440
rect 31528 42143 33500 42151
rect 27030 42100 31231 42143
rect 22692 41912 26748 42100
rect 20604 41620 22400 41912
tri 22400 41620 22692 41912 sw
tri 22692 41620 22984 41912 ne
rect 22984 41902 26748 41912
tri 26748 41902 26946 42100 sw
tri 27030 41902 27228 42100 ne
rect 27228 41917 31231 42100
tri 31231 41917 31457 42143 sw
tri 31528 41917 31754 42143 ne
rect 31754 41917 33500 42143
rect 27228 41902 31457 41917
rect 22984 41620 26946 41902
tri 26946 41620 27228 41902 sw
tri 27228 41620 27510 41902 ne
rect 27510 41620 31457 41902
tri 31457 41620 31754 41917 sw
tri 31754 41620 32051 41917 ne
rect 32051 41862 33500 41917
tri 33500 41862 33789 42151 sw
tri 33789 41862 34078 42151 ne
rect 34078 42150 35480 42151
tri 35480 42150 35770 42440 sw
tri 35770 42150 36060 42440 ne
rect 36060 42150 40014 42440
rect 34078 41862 35770 42150
rect 32051 41620 33789 41862
rect 20604 41328 22692 41620
tri 22692 41328 22984 41620 sw
tri 22984 41328 23276 41620 ne
rect 23276 41338 27228 41620
tri 27228 41338 27510 41620 sw
tri 27510 41338 27792 41620 ne
rect 27792 41338 31754 41620
rect 23276 41328 27510 41338
rect 20604 41036 22984 41328
tri 22984 41036 23276 41328 sw
tri 23276 41036 23568 41328 ne
rect 23568 41056 27510 41328
tri 27510 41056 27792 41338 sw
tri 27792 41056 28074 41338 ne
rect 28074 41323 31754 41338
tri 31754 41323 32051 41620 sw
tri 32051 41323 32348 41620 ne
rect 32348 41573 33789 41620
tri 33789 41573 34078 41862 sw
tri 34078 41573 34367 41862 ne
rect 34367 41860 35770 41862
tri 35770 41860 36060 42150 sw
tri 36060 41860 36350 42150 ne
rect 36350 42146 40014 42150
tri 40014 42146 40308 42440 sw
tri 40308 42146 40602 42440 ne
rect 40602 42156 44548 42440
tri 44548 42156 44836 42444 sw
tri 44836 42156 45124 42444 ne
rect 45124 42282 48945 42444
tri 48945 42282 49242 42579 sw
tri 49242 42282 49539 42579 ne
rect 49539 42440 53378 42579
tri 53378 42440 53625 42687 sw
tri 53671 42440 53918 42687 ne
rect 53918 42600 55538 42687
tri 55538 42600 55738 42800 sw
tri 55830 42600 56030 42800 ne
rect 56030 42600 57810 42800
tri 57810 42600 58010 42800 sw
rect 53918 42440 55738 42600
rect 49539 42282 53625 42440
rect 45124 42156 49242 42282
rect 40602 42146 44836 42156
rect 36350 41860 40308 42146
rect 34367 41573 36060 41860
rect 32348 41418 34078 41573
tri 34078 41418 34233 41573 sw
tri 34367 41418 34522 41573 ne
rect 34522 41570 36060 41573
tri 36060 41570 36350 41860 sw
tri 36350 41570 36640 41860 ne
rect 36640 41852 40308 41860
tri 40308 41852 40602 42146 sw
tri 40602 41852 40896 42146 ne
rect 40896 41976 44836 42146
tri 44836 41976 45016 42156 sw
tri 45124 41976 45304 42156 ne
rect 45304 41985 49242 42156
tri 49242 41985 49539 42282 sw
tri 49539 41985 49836 42282 ne
rect 49836 42147 53625 42282
tri 53625 42147 53918 42440 sw
tri 53918 42147 54211 42440 ne
rect 54211 42308 55738 42440
tri 55738 42308 56030 42600 sw
tri 56030 42308 56322 42600 ne
rect 56322 42497 71000 42600
rect 56322 42308 70613 42497
rect 54211 42147 56030 42308
rect 49836 41985 53918 42147
rect 45304 41976 49539 41985
rect 40896 41852 45016 41976
rect 36640 41570 40602 41852
rect 34522 41418 36350 41570
rect 32348 41323 34233 41418
rect 28074 41056 32051 41323
rect 23568 41036 27792 41056
rect 20604 40744 23276 41036
tri 23276 40744 23568 41036 sw
tri 23568 40744 23860 41036 ne
rect 23860 40774 27792 41036
tri 27792 40774 28074 41056 sw
tri 28074 40774 28356 41056 ne
rect 28356 41026 32051 41056
tri 32051 41026 32348 41323 sw
tri 32348 41026 32645 41323 ne
rect 32645 41129 34233 41323
tri 34233 41129 34522 41418 sw
tri 34522 41129 34811 41418 ne
rect 34811 41330 36350 41418
tri 36350 41330 36590 41570 sw
tri 36640 41330 36880 41570 ne
rect 36880 41558 40602 41570
tri 40602 41558 40896 41852 sw
tri 40896 41558 41190 41852 ne
rect 41190 41688 45016 41852
tri 45016 41688 45304 41976 sw
tri 45304 41688 45592 41976 ne
rect 45592 41688 49539 41976
tri 49539 41688 49836 41985 sw
tri 49836 41688 50133 41985 ne
rect 50133 41854 53918 41985
tri 53918 41854 54211 42147 sw
tri 54211 41854 54504 42147 ne
rect 54504 42016 56030 42147
tri 56030 42016 56322 42308 sw
tri 56322 42016 56614 42308 ne
rect 56614 42016 70613 42308
rect 54504 41854 56322 42016
rect 50133 41688 54211 41854
rect 41190 41558 45304 41688
rect 36880 41330 40896 41558
rect 34811 41129 36590 41330
rect 32645 41026 34522 41129
rect 28356 40774 32348 41026
rect 23860 40744 28074 40774
rect 20604 40632 23568 40744
tri 23568 40632 23680 40744 sw
tri 23860 40632 23972 40744 ne
rect 23972 40632 28074 40744
rect 20604 40340 23680 40632
tri 23680 40340 23972 40632 sw
tri 23972 40340 24264 40632 ne
rect 24264 40492 28074 40632
tri 28074 40492 28356 40774 sw
tri 28356 40492 28638 40774 ne
rect 28638 40757 32348 40774
tri 32348 40757 32617 41026 sw
tri 32645 40757 32914 41026 ne
rect 32914 40840 34522 41026
tri 34522 40840 34811 41129 sw
tri 34811 40840 35100 41129 ne
rect 35100 41040 36590 41129
tri 36590 41040 36880 41330 sw
tri 36880 41040 37170 41330 ne
rect 37170 41264 40896 41330
tri 40896 41264 41190 41558 sw
tri 41190 41264 41484 41558 ne
rect 41484 41400 45304 41558
tri 45304 41400 45592 41688 sw
tri 45592 41400 45880 41688 ne
rect 45880 41400 49836 41688
rect 41484 41264 45592 41400
rect 37170 41040 41190 41264
rect 35100 40840 36880 41040
rect 32914 40757 34811 40840
rect 28638 40492 32617 40757
rect 24264 40340 28356 40492
rect 20604 40048 23972 40340
tri 23972 40048 24264 40340 sw
tri 24264 40048 24556 40340 ne
rect 24556 40210 28356 40340
tri 28356 40210 28638 40492 sw
tri 28638 40210 28920 40492 ne
rect 28920 40460 32617 40492
tri 32617 40460 32914 40757 sw
tri 32914 40460 33211 40757 ne
rect 33211 40749 34811 40757
tri 34811 40749 34902 40840 sw
tri 35100 40749 35191 40840 ne
rect 35191 40750 36880 40840
tri 36880 40750 37170 41040 sw
tri 37170 40750 37460 41040 ne
rect 37460 41002 41190 41040
tri 41190 41002 41452 41264 sw
tri 41484 41002 41746 41264 ne
rect 41746 41112 45592 41264
tri 45592 41112 45880 41400 sw
tri 45880 41112 46168 41400 ne
rect 46168 41391 49836 41400
tri 49836 41391 50133 41688 sw
tri 50133 41391 50430 41688 ne
rect 50430 41586 54211 41688
tri 54211 41586 54479 41854 sw
tri 54504 41586 54772 41854 ne
rect 54772 41784 56322 41854
tri 56322 41784 56554 42016 sw
tri 56614 41784 56846 42016 ne
rect 56846 41784 70613 42016
rect 54772 41586 56554 41784
rect 50430 41391 54479 41586
rect 46168 41112 50133 41391
rect 41746 41002 45880 41112
rect 37460 40750 41452 41002
rect 35191 40749 37170 40750
rect 33211 40460 34902 40749
tri 34902 40460 35191 40749 sw
tri 35191 40460 35480 40749 ne
rect 35480 40460 37170 40749
tri 37170 40460 37460 40750 sw
tri 37460 40460 37750 40750 ne
rect 37750 40708 41452 40750
tri 41452 40708 41746 41002 sw
tri 41746 40708 42040 41002 ne
rect 42040 40824 45880 41002
tri 45880 40824 46168 41112 sw
tri 46168 40824 46456 41112 ne
rect 46456 41094 50133 41112
tri 50133 41094 50430 41391 sw
tri 50430 41094 50727 41391 ne
rect 50727 41293 54479 41391
tri 54479 41293 54772 41586 sw
tri 54772 41293 55065 41586 ne
rect 55065 41492 56554 41586
tri 56554 41492 56846 41784 sw
tri 56846 41492 57138 41784 ne
rect 57138 41492 70613 41784
rect 55065 41293 56846 41492
rect 50727 41094 54772 41293
rect 46456 41054 50430 41094
tri 50430 41054 50470 41094 sw
tri 50727 41054 50767 41094 ne
rect 50767 41054 54772 41094
rect 46456 40824 50470 41054
rect 42040 40708 46168 40824
rect 37750 40460 41746 40708
rect 28920 40210 32914 40460
rect 24556 40112 28638 40210
tri 28638 40112 28736 40210 sw
tri 28920 40112 29018 40210 ne
rect 29018 40163 32914 40210
tri 32914 40163 33211 40460 sw
tri 33211 40163 33508 40460 ne
rect 33508 40171 35191 40460
tri 35191 40171 35480 40460 sw
tri 35480 40171 35769 40460 ne
rect 35769 40171 37460 40460
rect 33508 40163 35480 40171
rect 29018 40112 33211 40163
rect 24556 40048 28736 40112
rect 20604 39756 24264 40048
tri 24264 39756 24556 40048 sw
tri 24556 39756 24848 40048 ne
rect 24848 39830 28736 40048
tri 28736 39830 29018 40112 sw
tri 29018 39830 29300 40112 ne
rect 29300 39866 33211 40112
tri 33211 39866 33508 40163 sw
tri 33508 39866 33805 40163 ne
rect 33805 39882 35480 40163
tri 35480 39882 35769 40171 sw
tri 35769 39882 36058 40171 ne
rect 36058 40170 37460 40171
tri 37460 40170 37750 40460 sw
tri 37750 40170 38040 40460 ne
rect 38040 40414 41746 40460
tri 41746 40414 42040 40708 sw
tri 42040 40414 42334 40708 ne
rect 42334 40536 46168 40708
tri 46168 40536 46456 40824 sw
tri 46456 40536 46744 40824 ne
rect 46744 40757 50470 40824
tri 50470 40757 50767 41054 sw
tri 50767 40757 51064 41054 ne
rect 51064 41000 54772 41054
tri 54772 41000 55065 41293 sw
tri 55065 41000 55358 41293 ne
rect 55358 41200 56846 41293
tri 56846 41200 57138 41492 sw
tri 57138 41200 57430 41492 ne
rect 57430 41297 70613 41492
rect 70669 41297 71000 42497
rect 57430 41200 71000 41297
rect 55358 41000 57138 41200
tri 57138 41000 57338 41200 sw
rect 51064 40937 55065 41000
tri 55065 40937 55128 41000 sw
tri 55358 40937 55421 41000 ne
rect 55421 40937 71000 41000
rect 51064 40757 55128 40937
rect 46744 40536 50767 40757
rect 42334 40414 46456 40536
rect 38040 40170 42040 40414
rect 36058 40112 37750 40170
tri 37750 40112 37808 40170 sw
tri 38040 40112 38098 40170 ne
rect 38098 40120 42040 40170
tri 42040 40120 42334 40414 sw
tri 42334 40120 42628 40414 ne
rect 42628 40248 46456 40414
tri 46456 40248 46744 40536 sw
tri 46744 40248 47032 40536 ne
rect 47032 40460 50767 40536
tri 50767 40460 51064 40757 sw
tri 51064 40460 51361 40757 ne
rect 51361 40644 55128 40757
tri 55128 40644 55421 40937 sw
tri 55421 40644 55714 40937 ne
rect 55714 40644 71000 40937
rect 51361 40460 55421 40644
rect 47032 40248 51064 40460
rect 42628 40216 46744 40248
tri 46744 40216 46776 40248 sw
tri 47032 40216 47064 40248 ne
rect 47064 40216 51064 40248
rect 42628 40120 46776 40216
rect 38098 40112 42334 40120
rect 36058 39882 37808 40112
rect 33805 39866 35769 39882
rect 29300 39830 33508 39866
rect 24848 39756 29018 39830
rect 20604 39464 24556 39756
tri 24556 39464 24848 39756 sw
tri 24848 39464 25140 39756 ne
rect 25140 39548 29018 39756
tri 29018 39548 29300 39830 sw
tri 29300 39548 29582 39830 ne
rect 29582 39829 33508 39830
tri 33508 39829 33545 39866 sw
tri 33805 39829 33842 39866 ne
rect 33842 39829 35769 39866
rect 29582 39548 33545 39829
rect 25140 39464 29300 39548
tri 20604 35220 24848 39464 ne
tri 24848 39172 25140 39464 sw
tri 25140 39172 25432 39464 ne
rect 25432 39266 29300 39464
tri 29300 39266 29582 39548 sw
tri 29582 39266 29864 39548 ne
rect 29864 39532 33545 39548
tri 33545 39532 33842 39829 sw
tri 33842 39532 34139 39829 ne
rect 34139 39593 35769 39829
tri 35769 39593 36058 39882 sw
tri 36058 39593 36347 39882 ne
rect 36347 39822 37808 39882
tri 37808 39822 38098 40112 sw
tri 38098 39822 38388 40112 ne
rect 38388 39826 42334 40112
tri 42334 39826 42628 40120 sw
tri 42628 39826 42922 40120 ne
rect 42922 39928 46776 40120
tri 46776 39928 47064 40216 sw
tri 47064 39928 47352 40216 ne
rect 47352 40163 51064 40216
tri 51064 40163 51361 40460 sw
tri 51361 40163 51658 40460 ne
rect 51658 40351 55421 40460
tri 55421 40351 55714 40644 sw
tri 55714 40351 56007 40644 ne
rect 56007 40351 71000 40644
rect 51658 40163 55714 40351
rect 47352 39928 51361 40163
rect 42922 39826 47064 39928
rect 38388 39822 42628 39826
rect 36347 39593 38098 39822
rect 34139 39532 36058 39593
rect 29864 39266 33842 39532
rect 25432 39172 29582 39266
rect 24848 38880 25140 39172
tri 25140 38880 25432 39172 sw
tri 25432 38880 25724 39172 ne
rect 25724 38984 29582 39172
tri 29582 38984 29864 39266 sw
tri 29864 38984 30146 39266 ne
rect 30146 39235 33842 39266
tri 33842 39235 34139 39532 sw
tri 34139 39235 34436 39532 ne
rect 34436 39438 36058 39532
tri 36058 39438 36213 39593 sw
tri 36347 39438 36502 39593 ne
rect 36502 39532 38098 39593
tri 38098 39532 38388 39822 sw
tri 38388 39532 38678 39822 ne
rect 38678 39532 42628 39822
tri 42628 39532 42922 39826 sw
tri 42922 39532 43216 39826 ne
rect 43216 39640 47064 39826
tri 47064 39640 47352 39928 sw
tri 47352 39640 47640 39928 ne
rect 47640 39866 51361 39928
tri 51361 39866 51658 40163 sw
tri 51658 39866 51955 40163 ne
rect 51955 40058 55714 40163
tri 55714 40058 56007 40351 sw
tri 56007 40058 56300 40351 ne
rect 56300 40058 71000 40351
rect 51955 39986 56007 40058
tri 56007 39986 56079 40058 sw
tri 56300 39986 56372 40058 ne
rect 56372 39986 71000 40058
rect 51955 39866 56079 39986
rect 47640 39640 51658 39866
rect 43216 39532 47352 39640
rect 36502 39438 38388 39532
rect 34436 39235 36213 39438
rect 30146 39157 34139 39235
tri 34139 39157 34217 39235 sw
tri 34436 39157 34514 39235 ne
rect 34514 39157 36213 39235
rect 30146 38984 34217 39157
rect 25724 38880 29864 38984
rect 24848 38588 25432 38880
tri 25432 38588 25724 38880 sw
tri 25724 38588 26016 38880 ne
rect 26016 38702 29864 38880
tri 29864 38702 30146 38984 sw
tri 30146 38702 30428 38984 ne
rect 30428 38860 34217 38984
tri 34217 38860 34514 39157 sw
tri 34514 38860 34811 39157 ne
rect 34811 39149 36213 39157
tri 36213 39149 36502 39438 sw
tri 36502 39149 36791 39438 ne
rect 36791 39242 38388 39438
tri 38388 39242 38678 39532 sw
tri 38678 39242 38968 39532 ne
rect 38968 39242 42922 39532
rect 36791 39149 38678 39242
rect 34811 38860 36502 39149
tri 36502 38860 36791 39149 sw
tri 36791 38860 37080 39149 ne
rect 37080 38952 38678 39149
tri 38678 38952 38968 39242 sw
tri 38968 38952 39258 39242 ne
rect 39258 39238 42922 39242
tri 42922 39238 43216 39532 sw
tri 43216 39238 43510 39532 ne
rect 43510 39352 47352 39532
tri 47352 39352 47640 39640 sw
tri 47640 39352 47928 39640 ne
rect 47928 39569 51658 39640
tri 51658 39569 51955 39866 sw
tri 51955 39569 52252 39866 ne
rect 52252 39693 56079 39866
tri 56079 39693 56372 39986 sw
tri 56372 39693 56665 39986 ne
rect 56665 39693 71000 39986
rect 52252 39569 56372 39693
rect 47928 39352 51955 39569
rect 43510 39238 47640 39352
rect 39258 38952 43216 39238
rect 37080 38860 38968 38952
rect 30428 38702 34514 38860
rect 26016 38588 30146 38702
rect 24848 38296 25724 38588
tri 25724 38296 26016 38588 sw
tri 26016 38296 26308 38588 ne
rect 26308 38420 30146 38588
tri 30146 38420 30428 38702 sw
tri 30428 38420 30710 38702 ne
rect 30710 38563 34514 38702
tri 34514 38563 34811 38860 sw
tri 34811 38563 35108 38860 ne
rect 35108 38769 36791 38860
tri 36791 38769 36882 38860 sw
tri 37080 38769 37171 38860 ne
rect 37171 38770 38968 38860
tri 38968 38770 39150 38952 sw
tri 39258 38770 39440 38952 ne
rect 39440 38944 43216 38952
tri 43216 38944 43510 39238 sw
tri 43510 38944 43804 39238 ne
rect 43804 39064 47640 39238
tri 47640 39064 47928 39352 sw
tri 47928 39064 48216 39352 ne
rect 48216 39272 51955 39352
tri 51955 39272 52252 39569 sw
tri 52252 39272 52549 39569 ne
rect 52549 39400 56372 39569
tri 56372 39400 56665 39693 sw
tri 56665 39600 56758 39693 ne
rect 56758 39600 71000 39693
rect 52549 39332 71000 39400
rect 52549 39272 70613 39332
rect 48216 39064 52252 39272
rect 43804 38944 47928 39064
rect 39440 38774 43510 38944
tri 43510 38774 43680 38944 sw
tri 43804 38774 43974 38944 ne
rect 43974 38776 47928 38944
tri 47928 38776 48216 39064 sw
tri 48216 38776 48504 39064 ne
rect 48504 38975 52252 39064
tri 52252 38975 52549 39272 sw
tri 52549 38975 52846 39272 ne
rect 52846 38975 70613 39272
rect 48504 38929 52549 38975
tri 52549 38929 52595 38975 sw
tri 52846 38929 52892 38975 ne
rect 52892 38929 70613 38975
rect 48504 38776 52595 38929
rect 43974 38774 48216 38776
rect 39440 38770 43680 38774
rect 37171 38769 39150 38770
rect 35108 38563 36882 38769
rect 30710 38480 34811 38563
tri 34811 38480 34894 38563 sw
tri 35108 38480 35191 38563 ne
rect 35191 38480 36882 38563
tri 36882 38480 37171 38769 sw
tri 37171 38480 37460 38769 ne
rect 37460 38480 39150 38769
tri 39150 38480 39440 38770 sw
tri 39440 38480 39730 38770 ne
rect 39730 38480 43680 38770
tri 43680 38480 43974 38774 sw
tri 43974 38480 44268 38774 ne
rect 44268 38488 48216 38774
tri 48216 38488 48504 38776 sw
tri 48504 38488 48792 38776 ne
rect 48792 38632 52595 38776
tri 52595 38632 52892 38929 sw
tri 52892 38632 53189 38929 ne
rect 53189 38632 70613 38929
rect 48792 38488 52892 38632
rect 44268 38480 48504 38488
rect 30710 38420 34894 38480
rect 26308 38296 30428 38420
rect 24848 38252 26016 38296
tri 26016 38252 26060 38296 sw
tri 26308 38252 26352 38296 ne
rect 26352 38252 30428 38296
rect 24848 37960 26060 38252
tri 26060 37960 26352 38252 sw
tri 26352 37960 26644 38252 ne
rect 26644 38138 30428 38252
tri 30428 38138 30710 38420 sw
tri 30710 38138 30992 38420 ne
rect 30992 38183 34894 38420
tri 34894 38183 35191 38480 sw
tri 35191 38183 35488 38480 ne
rect 35488 38191 37171 38480
tri 37171 38191 37460 38480 sw
tri 37460 38191 37749 38480 ne
rect 37749 38191 39440 38480
rect 35488 38183 37460 38191
rect 30992 38138 35191 38183
rect 26644 37960 30710 38138
rect 24848 37668 26352 37960
tri 26352 37668 26644 37960 sw
tri 26644 37668 26936 37960 ne
rect 26936 37856 30710 37960
tri 30710 37856 30992 38138 sw
tri 30992 37856 31274 38138 ne
rect 31274 37970 35191 38138
tri 35191 37970 35404 38183 sw
tri 35488 37970 35701 38183 ne
rect 35701 37970 37460 38183
rect 31274 37856 35404 37970
rect 26936 37668 30992 37856
rect 24848 37376 26644 37668
tri 26644 37376 26936 37668 sw
tri 26936 37376 27228 37668 ne
rect 27228 37658 30992 37668
tri 30992 37658 31190 37856 sw
tri 31274 37658 31472 37856 ne
rect 31472 37673 35404 37856
tri 35404 37673 35701 37970 sw
tri 35701 37673 35998 37970 ne
rect 35998 37902 37460 37970
tri 37460 37902 37749 38191 sw
tri 37749 37902 38038 38191 ne
rect 38038 38190 39440 38191
tri 39440 38190 39730 38480 sw
tri 39730 38190 40020 38480 ne
rect 40020 38190 43974 38480
rect 38038 37902 39730 38190
rect 35998 37673 37749 37902
rect 31472 37658 35701 37673
rect 27228 37376 31190 37658
tri 31190 37376 31472 37658 sw
tri 31472 37376 31754 37658 ne
rect 31754 37376 35701 37658
tri 35701 37376 35998 37673 sw
tri 35998 37376 36295 37673 ne
rect 36295 37613 37749 37673
tri 37749 37613 38038 37902 sw
tri 38038 37613 38327 37902 ne
rect 38327 37900 39730 37902
tri 39730 37900 40020 38190 sw
tri 40020 37900 40310 38190 ne
rect 40310 38186 43974 38190
tri 43974 38186 44268 38480 sw
tri 44268 38186 44562 38480 ne
rect 44562 38200 48504 38480
tri 48504 38200 48792 38488 sw
tri 48792 38200 49080 38488 ne
rect 49080 38335 52892 38488
tri 52892 38335 53189 38632 sw
tri 53189 38335 53486 38632 ne
rect 53486 38335 70613 38632
rect 49080 38200 53189 38335
rect 44562 38186 48792 38200
rect 40310 37900 44268 38186
rect 38327 37613 40020 37900
rect 36295 37458 38038 37613
tri 38038 37458 38193 37613 sw
tri 38327 37458 38482 37613 ne
rect 38482 37610 40020 37613
tri 40020 37610 40310 37900 sw
tri 40310 37610 40600 37900 ne
rect 40600 37892 44268 37900
tri 44268 37892 44562 38186 sw
tri 44562 37892 44856 38186 ne
rect 44856 37912 48792 38186
tri 48792 37912 49080 38200 sw
tri 49080 37912 49368 38200 ne
rect 49368 38038 53189 38200
tri 53189 38038 53486 38335 sw
tri 53486 38038 53783 38335 ne
rect 53783 38038 70613 38335
rect 49368 37912 53486 38038
rect 44856 37892 49080 37912
rect 40600 37610 44562 37892
rect 38482 37458 40310 37610
rect 36295 37376 38193 37458
rect 24848 37084 26936 37376
tri 26936 37084 27228 37376 sw
tri 27228 37084 27520 37376 ne
rect 27520 37094 31472 37376
tri 31472 37094 31754 37376 sw
tri 31754 37094 32036 37376 ne
rect 32036 37094 35998 37376
rect 27520 37084 31754 37094
rect 24848 36792 27228 37084
tri 27228 36792 27520 37084 sw
tri 27520 36792 27812 37084 ne
rect 27812 36812 31754 37084
tri 31754 36812 32036 37094 sw
tri 32036 36812 32318 37094 ne
rect 32318 37079 35998 37094
tri 35998 37079 36295 37376 sw
tri 36295 37079 36592 37376 ne
rect 36592 37169 38193 37376
tri 38193 37169 38482 37458 sw
tri 38482 37169 38771 37458 ne
rect 38771 37370 40310 37458
tri 40310 37370 40550 37610 sw
tri 40600 37370 40840 37610 ne
rect 40840 37598 44562 37610
tri 44562 37598 44856 37892 sw
tri 44856 37598 45150 37892 ne
rect 45150 37732 49080 37892
tri 49080 37732 49260 37912 sw
tri 49368 37732 49548 37912 ne
rect 49548 37741 53486 37912
tri 53486 37741 53783 38038 sw
tri 53783 37741 54080 38038 ne
rect 54080 37741 70613 38038
rect 49548 37732 53783 37741
rect 45150 37598 49260 37732
rect 40840 37370 44856 37598
rect 38771 37169 40550 37370
rect 36592 37079 38482 37169
rect 32318 36812 36295 37079
rect 27812 36792 32036 36812
rect 24848 36500 27520 36792
tri 27520 36500 27812 36792 sw
tri 27812 36500 28104 36792 ne
rect 28104 36530 32036 36792
tri 32036 36530 32318 36812 sw
tri 32318 36530 32600 36812 ne
rect 32600 36797 36295 36812
tri 36295 36797 36577 37079 sw
tri 36592 36797 36874 37079 ne
rect 36874 36880 38482 37079
tri 38482 36880 38771 37169 sw
tri 38771 36880 39060 37169 ne
rect 39060 37080 40550 37169
tri 40550 37080 40840 37370 sw
tri 40840 37080 41130 37370 ne
rect 41130 37304 44856 37370
tri 44856 37304 45150 37598 sw
tri 45150 37304 45444 37598 ne
rect 45444 37444 49260 37598
tri 49260 37444 49548 37732 sw
tri 49548 37444 49836 37732 ne
rect 49836 37444 53783 37732
tri 53783 37444 54080 37741 sw
tri 54080 37444 54377 37741 ne
rect 54377 37444 70613 37741
rect 45444 37304 49548 37444
rect 41130 37080 45150 37304
rect 39060 36880 40840 37080
rect 36874 36797 38771 36880
rect 32600 36530 36577 36797
rect 28104 36500 32318 36530
rect 24848 36388 27812 36500
tri 27812 36388 27924 36500 sw
tri 28104 36388 28216 36500 ne
rect 28216 36388 32318 36500
rect 24848 36096 27924 36388
tri 27924 36096 28216 36388 sw
tri 28216 36096 28508 36388 ne
rect 28508 36248 32318 36388
tri 32318 36248 32600 36530 sw
tri 32600 36248 32882 36530 ne
rect 32882 36500 36577 36530
tri 36577 36500 36874 36797 sw
tri 36874 36500 37171 36797 ne
rect 37171 36789 38771 36797
tri 38771 36789 38862 36880 sw
tri 39060 36789 39151 36880 ne
rect 39151 36790 40840 36880
tri 40840 36790 41130 37080 sw
tri 41130 36790 41420 37080 ne
rect 41420 37010 45150 37080
tri 45150 37010 45444 37304 sw
tri 45444 37010 45738 37304 ne
rect 45738 37156 49548 37304
tri 49548 37156 49836 37444 sw
tri 49836 37156 50124 37444 ne
rect 50124 37156 54080 37444
rect 45738 37010 49836 37156
rect 41420 36790 45444 37010
rect 39151 36789 41130 36790
rect 37171 36500 38862 36789
tri 38862 36500 39151 36789 sw
tri 39151 36500 39440 36789 ne
rect 39440 36500 41130 36789
tri 41130 36500 41420 36790 sw
tri 41420 36500 41710 36790 ne
rect 41710 36758 45444 36790
tri 45444 36758 45696 37010 sw
tri 45738 36758 45990 37010 ne
rect 45990 36868 49836 37010
tri 49836 36868 50124 37156 sw
tri 50124 36868 50412 37156 ne
rect 50412 37147 54080 37156
tri 54080 37147 54377 37444 sw
tri 54377 37147 54674 37444 ne
rect 54674 37147 70613 37444
rect 50412 36868 54377 37147
rect 45990 36758 50124 36868
rect 41710 36500 45696 36758
rect 32882 36248 36874 36500
rect 28508 36096 32600 36248
rect 24848 35804 28216 36096
tri 28216 35804 28508 36096 sw
tri 28508 35804 28800 36096 ne
rect 28800 35966 32600 36096
tri 32600 35966 32882 36248 sw
tri 32882 35966 33164 36248 ne
rect 33164 36203 36874 36248
tri 36874 36203 37171 36500 sw
tri 37171 36203 37468 36500 ne
rect 37468 36211 39151 36500
tri 39151 36211 39440 36500 sw
tri 39440 36211 39729 36500 ne
rect 39729 36211 41420 36500
rect 37468 36203 39440 36211
rect 33164 35966 37171 36203
rect 28800 35868 32882 35966
tri 32882 35868 32980 35966 sw
tri 33164 35868 33262 35966 ne
rect 33262 35906 37171 35966
tri 37171 35906 37468 36203 sw
tri 37468 35906 37765 36203 ne
rect 37765 35922 39440 36203
tri 39440 35922 39729 36211 sw
tri 39729 35922 40018 36211 ne
rect 40018 36210 41420 36211
tri 41420 36210 41710 36500 sw
tri 41710 36210 42000 36500 ne
rect 42000 36464 45696 36500
tri 45696 36464 45990 36758 sw
tri 45990 36464 46284 36758 ne
rect 46284 36580 50124 36758
tri 50124 36580 50412 36868 sw
tri 50412 36580 50700 36868 ne
rect 50700 36850 54377 36868
tri 54377 36850 54674 37147 sw
tri 54674 36850 54971 37147 ne
rect 54971 36850 70613 37147
rect 50700 36794 54674 36850
tri 54674 36794 54730 36850 sw
tri 54971 36794 55027 36850 ne
rect 55027 36794 70613 36850
rect 50700 36580 54730 36794
rect 46284 36464 50412 36580
rect 42000 36210 45990 36464
rect 40018 35922 41710 36210
rect 37765 35906 39729 35922
rect 33262 35882 37468 35906
tri 37468 35882 37492 35906 sw
tri 37765 35882 37789 35906 ne
rect 37789 35882 39729 35906
rect 33262 35868 37492 35882
rect 28800 35804 32980 35868
rect 24848 35512 28508 35804
tri 28508 35512 28800 35804 sw
tri 28800 35512 29092 35804 ne
rect 29092 35586 32980 35804
tri 32980 35586 33262 35868 sw
tri 33262 35586 33544 35868 ne
rect 33544 35586 37492 35868
rect 29092 35512 33262 35586
rect 24848 35220 28800 35512
tri 28800 35220 29092 35512 sw
tri 29092 35220 29384 35512 ne
rect 29384 35304 33262 35512
tri 33262 35304 33544 35586 sw
tri 33544 35304 33826 35586 ne
rect 33826 35585 37492 35586
tri 37492 35585 37789 35882 sw
tri 37789 35585 38086 35882 ne
rect 38086 35633 39729 35882
tri 39729 35633 40018 35922 sw
tri 40018 35633 40307 35922 ne
rect 40307 35920 41710 35922
tri 41710 35920 42000 36210 sw
tri 42000 35920 42290 36210 ne
rect 42290 36170 45990 36210
tri 45990 36170 46284 36464 sw
tri 46284 36170 46578 36464 ne
rect 46578 36292 50412 36464
tri 50412 36292 50700 36580 sw
tri 50700 36292 50988 36580 ne
rect 50988 36497 54730 36580
tri 54730 36497 55027 36794 sw
tri 55027 36497 55324 36794 ne
rect 55324 36497 70613 36794
rect 50988 36292 55027 36497
rect 46578 36170 50700 36292
rect 42290 35920 46284 36170
rect 40307 35868 42000 35920
tri 42000 35868 42052 35920 sw
tri 42290 35868 42342 35920 ne
rect 42342 35876 46284 35920
tri 46284 35876 46578 36170 sw
tri 46578 35876 46872 36170 ne
rect 46872 36004 50700 36170
tri 50700 36004 50988 36292 sw
tri 50988 36004 51276 36292 ne
rect 51276 36200 55027 36292
tri 55027 36200 55324 36497 sw
tri 55324 36400 55421 36497 ne
rect 55421 36468 70613 36497
rect 70669 36468 71000 39332
rect 55421 36400 71000 36468
rect 51276 36132 71000 36200
rect 51276 36004 70613 36132
rect 46872 35972 50988 36004
tri 50988 35972 51020 36004 sw
tri 51276 35972 51308 36004 ne
rect 51308 35972 70613 36004
rect 46872 35876 51020 35972
rect 42342 35868 46578 35876
rect 40307 35633 42052 35868
rect 38086 35585 40018 35633
rect 33826 35304 37789 35585
rect 29384 35220 33544 35304
tri 24848 30976 29092 35220 ne
tri 29092 34928 29384 35220 sw
tri 29384 34928 29676 35220 ne
rect 29676 35022 33544 35220
tri 33544 35022 33826 35304 sw
tri 33826 35022 34108 35304 ne
rect 34108 35288 37789 35304
tri 37789 35288 38086 35585 sw
tri 38086 35288 38383 35585 ne
rect 38383 35409 40018 35585
tri 40018 35409 40242 35633 sw
tri 40307 35478 40462 35633 ne
rect 40462 35578 42052 35633
tri 42052 35578 42342 35868 sw
tri 42342 35578 42632 35868 ne
rect 42632 35582 46578 35868
tri 46578 35582 46872 35876 sw
tri 46872 35582 47166 35876 ne
rect 47166 35684 51020 35876
tri 51020 35684 51308 35972 sw
tri 51308 35684 51596 35972 ne
rect 51596 35684 70613 35972
rect 47166 35582 51308 35684
rect 42632 35578 46872 35582
rect 40462 35478 42342 35578
rect 38383 35288 40242 35409
rect 34108 35022 38086 35288
rect 29676 34928 33826 35022
rect 29092 34636 29384 34928
tri 29384 34636 29676 34928 sw
tri 29676 34636 29968 34928 ne
rect 29968 34740 33826 34928
tri 33826 34740 34108 35022 sw
tri 34108 34740 34390 35022 ne
rect 34390 34991 38086 35022
tri 38086 34991 38383 35288 sw
tri 38383 34991 38680 35288 ne
rect 38680 35189 40242 35288
tri 40242 35189 40462 35409 sw
tri 40462 35189 40751 35478 ne
rect 40751 35288 42342 35478
tri 42342 35288 42632 35578 sw
tri 42632 35288 42922 35578 ne
rect 42922 35288 46872 35578
tri 46872 35288 47166 35582 sw
tri 47166 35288 47460 35582 ne
rect 47460 35396 51308 35582
tri 51308 35396 51596 35684 sw
tri 51596 35396 51884 35684 ne
rect 51884 35396 70613 35684
rect 47460 35288 51596 35396
rect 40751 35189 42632 35288
rect 38680 34991 40462 35189
rect 34390 34900 38383 34991
tri 38383 34900 38474 34991 sw
tri 38680 34900 38771 34991 ne
rect 38771 34900 40462 34991
tri 40462 34900 40751 35189 sw
tri 40751 34900 41040 35189 ne
rect 41040 34998 42632 35189
tri 42632 34998 42922 35288 sw
tri 42922 34998 43212 35288 ne
rect 43212 34998 47166 35288
rect 41040 34900 42922 34998
rect 34390 34740 38474 34900
rect 29968 34636 34108 34740
rect 29092 34344 29676 34636
tri 29676 34344 29968 34636 sw
tri 29968 34344 30260 34636 ne
rect 30260 34458 34108 34636
tri 34108 34458 34390 34740 sw
tri 34390 34458 34672 34740 ne
rect 34672 34603 38474 34740
tri 38474 34603 38771 34900 sw
tri 38771 34603 39068 34900 ne
rect 39068 34809 40751 34900
tri 40751 34809 40842 34900 sw
tri 41040 34809 41131 34900 ne
rect 41131 34809 42922 34900
rect 39068 34603 40842 34809
rect 34672 34520 38771 34603
tri 38771 34520 38854 34603 sw
tri 39068 34520 39151 34603 ne
rect 39151 34520 40842 34603
tri 40842 34520 41131 34809 sw
tri 41131 34520 41420 34809 ne
rect 41420 34708 42922 34809
tri 42922 34708 43212 34998 sw
tri 43212 34708 43502 34998 ne
rect 43502 34994 47166 34998
tri 47166 34994 47460 35288 sw
tri 47460 34994 47754 35288 ne
rect 47754 35108 51596 35288
tri 51596 35108 51884 35396 sw
tri 51884 35108 52172 35396 ne
rect 52172 35108 70613 35396
rect 47754 34994 51884 35108
rect 43502 34708 47460 34994
rect 41420 34534 43212 34708
tri 43212 34534 43386 34708 sw
tri 43502 34534 43676 34708 ne
rect 43676 34700 47460 34708
tri 47460 34700 47754 34994 sw
tri 47754 34700 48048 34994 ne
rect 48048 34820 51884 34994
tri 51884 34820 52172 35108 sw
tri 52172 34820 52460 35108 ne
rect 52460 34820 70613 35108
rect 48048 34700 52172 34820
rect 43676 34538 47754 34700
tri 47754 34538 47916 34700 sw
tri 48048 34538 48210 34700 ne
rect 48210 34538 52172 34700
rect 43676 34534 47916 34538
rect 41420 34520 43386 34534
rect 34672 34458 38854 34520
rect 30260 34344 34390 34458
rect 29092 34052 29968 34344
tri 29968 34052 30260 34344 sw
tri 30260 34052 30552 34344 ne
rect 30552 34176 34390 34344
tri 34390 34176 34672 34458 sw
tri 34672 34176 34954 34458 ne
rect 34954 34223 38854 34458
tri 38854 34223 39151 34520 sw
tri 39151 34223 39448 34520 ne
rect 39448 34231 41131 34520
tri 41131 34231 41420 34520 sw
tri 41420 34231 41709 34520 ne
rect 41709 34244 43386 34520
tri 43386 34244 43676 34534 sw
tri 43676 34244 43966 34534 ne
rect 43966 34244 47916 34534
tri 47916 34244 48210 34538 sw
tri 48210 34244 48504 34538 ne
rect 48504 34532 52172 34538
tri 52172 34532 52460 34820 sw
tri 52460 34532 52748 34820 ne
rect 52748 34532 70613 34820
rect 48504 34244 52460 34532
tri 52460 34244 52748 34532 sw
tri 52748 34244 53036 34532 ne
rect 53036 34244 70613 34532
rect 41709 34231 43676 34244
rect 39448 34223 41420 34231
rect 34954 34176 39151 34223
rect 30552 34052 34672 34176
rect 29092 34008 30260 34052
tri 30260 34008 30304 34052 sw
tri 30552 34008 30596 34052 ne
rect 30596 34008 34672 34052
rect 29092 33716 30304 34008
tri 30304 33716 30596 34008 sw
tri 30596 33716 30888 34008 ne
rect 30888 33894 34672 34008
tri 34672 33894 34954 34176 sw
tri 34954 33894 35236 34176 ne
rect 35236 33926 39151 34176
tri 39151 33926 39448 34223 sw
tri 39448 33926 39745 34223 ne
rect 39745 33942 41420 34223
tri 41420 33942 41709 34231 sw
tri 41709 33942 41998 34231 ne
rect 41998 33954 43676 34231
tri 43676 33954 43966 34244 sw
tri 43966 33954 44256 34244 ne
rect 44256 33954 48210 34244
rect 41998 33942 43966 33954
rect 39745 33926 41709 33942
rect 35236 33894 39448 33926
rect 30888 33716 34954 33894
rect 29092 33424 30596 33716
tri 30596 33424 30888 33716 sw
tri 30888 33424 31180 33716 ne
rect 31180 33612 34954 33716
tri 34954 33612 35236 33894 sw
tri 35236 33612 35518 33894 ne
rect 35518 33726 39448 33894
tri 39448 33726 39648 33926 sw
tri 39745 33726 39945 33926 ne
rect 39945 33726 41709 33926
rect 35518 33612 39648 33726
rect 31180 33424 35236 33612
rect 29092 33132 30888 33424
tri 30888 33132 31180 33424 sw
tri 31180 33132 31472 33424 ne
rect 31472 33414 35236 33424
tri 35236 33414 35434 33612 sw
tri 35518 33414 35716 33612 ne
rect 35716 33429 39648 33612
tri 39648 33429 39945 33726 sw
tri 39945 33429 40242 33726 ne
rect 40242 33653 41709 33726
tri 41709 33653 41998 33942 sw
tri 41998 33653 42287 33942 ne
rect 42287 33664 43966 33942
tri 43966 33664 44256 33954 sw
tri 44256 33664 44546 33954 ne
rect 44546 33950 48210 33954
tri 48210 33950 48504 34244 sw
tri 48504 33950 48798 34244 ne
rect 48798 33956 52748 34244
tri 52748 33956 53036 34244 sw
tri 53036 33956 53324 34244 ne
rect 53324 33956 70613 34244
rect 48798 33950 53036 33956
rect 44546 33664 48504 33950
rect 42287 33653 44256 33664
rect 40242 33498 41998 33653
tri 41998 33498 42153 33653 sw
tri 42287 33498 42442 33653 ne
rect 42442 33498 44256 33653
rect 40242 33429 42153 33498
rect 35716 33414 39945 33429
rect 31472 33132 35434 33414
tri 35434 33132 35716 33414 sw
tri 35716 33132 35998 33414 ne
rect 35998 33132 39945 33414
tri 39945 33132 40242 33429 sw
tri 40242 33132 40539 33429 ne
rect 40539 33209 42153 33429
tri 42153 33209 42442 33498 sw
tri 42442 33209 42731 33498 ne
rect 42731 33410 44256 33498
tri 44256 33410 44510 33664 sw
tri 44546 33410 44800 33664 ne
rect 44800 33656 48504 33664
tri 48504 33656 48798 33950 sw
tri 48798 33656 49092 33950 ne
rect 49092 33668 53036 33950
tri 53036 33668 53324 33956 sw
tri 53324 33668 53612 33956 ne
rect 53612 33668 70613 33956
rect 49092 33656 53324 33668
rect 44800 33410 48798 33656
rect 42731 33209 44510 33410
rect 40539 33132 42442 33209
rect 29092 32840 31180 33132
tri 31180 32840 31472 33132 sw
tri 31472 32840 31764 33132 ne
rect 31764 32850 35716 33132
tri 35716 32850 35998 33132 sw
tri 35998 32850 36280 33132 ne
rect 36280 32850 40242 33132
rect 31764 32840 35998 32850
rect 29092 32548 31472 32840
tri 31472 32548 31764 32840 sw
tri 31764 32548 32056 32840 ne
rect 32056 32568 35998 32840
tri 35998 32568 36280 32850 sw
tri 36280 32568 36562 32850 ne
rect 36562 32835 40242 32850
tri 40242 32835 40539 33132 sw
tri 40539 32835 40836 33132 ne
rect 40836 32920 42442 33132
tri 42442 32920 42731 33209 sw
tri 42731 32920 43020 33209 ne
rect 43020 33120 44510 33209
tri 44510 33120 44800 33410 sw
tri 44800 33120 45090 33410 ne
rect 45090 33362 48798 33410
tri 48798 33362 49092 33656 sw
tri 49092 33362 49386 33656 ne
rect 49386 33576 53324 33656
tri 53324 33576 53416 33668 sw
tri 53612 33576 53704 33668 ne
rect 53704 33576 70613 33668
rect 49386 33362 53416 33576
rect 45090 33120 49092 33362
rect 43020 32920 44800 33120
rect 40836 32835 42731 32920
rect 36562 32568 40539 32835
rect 32056 32548 36280 32568
rect 29092 32256 31764 32548
tri 31764 32256 32056 32548 sw
tri 32056 32256 32348 32548 ne
rect 32348 32286 36280 32548
tri 36280 32286 36562 32568 sw
tri 36562 32286 36844 32568 ne
rect 36844 32540 40539 32568
tri 40539 32540 40834 32835 sw
tri 40836 32540 41131 32835 ne
rect 41131 32829 42731 32835
tri 42731 32829 42822 32920 sw
tri 43020 32829 43111 32920 ne
rect 43111 32830 44800 32920
tri 44800 32830 45090 33120 sw
tri 45090 32830 45380 33120 ne
rect 45380 33068 49092 33120
tri 49092 33068 49386 33362 sw
tri 49386 33068 49680 33362 ne
rect 49680 33288 53416 33362
tri 53416 33288 53704 33576 sw
tri 53704 33288 53992 33576 ne
rect 53992 33288 70613 33576
rect 49680 33068 53704 33288
rect 45380 32830 49386 33068
rect 43111 32829 45090 32830
rect 41131 32540 42822 32829
tri 42822 32540 43111 32829 sw
tri 43111 32540 43400 32829 ne
rect 43400 32540 45090 32829
tri 45090 32540 45380 32830 sw
tri 45380 32540 45670 32830 ne
rect 45670 32774 49386 32830
tri 49386 32774 49680 33068 sw
tri 49680 32774 49974 33068 ne
rect 49974 33000 53704 33068
tri 53704 33000 53992 33288 sw
tri 53992 33200 54080 33288 ne
rect 54080 33268 70613 33288
rect 70669 33268 71000 36132
rect 54080 33200 71000 33268
rect 49974 32920 71000 33000
rect 49974 32774 70613 32920
rect 45670 32540 49680 32774
rect 36844 32286 40834 32540
rect 32348 32256 36562 32286
rect 29092 32144 32056 32256
tri 32056 32144 32168 32256 sw
tri 32348 32144 32460 32256 ne
rect 32460 32144 36562 32256
rect 29092 31852 32168 32144
tri 32168 31852 32460 32144 sw
tri 32460 31852 32752 32144 ne
rect 32752 32004 36562 32144
tri 36562 32004 36844 32286 sw
tri 36844 32004 37126 32286 ne
rect 37126 32243 40834 32286
tri 40834 32243 41131 32540 sw
tri 41131 32243 41428 32540 ne
rect 41428 32251 43111 32540
tri 43111 32251 43400 32540 sw
tri 43400 32251 43689 32540 ne
rect 43689 32251 45380 32540
rect 41428 32243 43400 32251
rect 37126 32004 41131 32243
rect 32752 31852 36844 32004
rect 29092 31560 32460 31852
tri 32460 31560 32752 31852 sw
tri 32752 31560 33044 31852 ne
rect 33044 31722 36844 31852
tri 36844 31722 37126 32004 sw
tri 37126 31722 37408 32004 ne
rect 37408 31946 41131 32004
tri 41131 31946 41428 32243 sw
tri 41428 31946 41725 32243 ne
rect 41725 31962 43400 32243
tri 43400 31962 43689 32251 sw
tri 43689 31962 43978 32251 ne
rect 43978 32250 45380 32251
tri 45380 32250 45670 32540 sw
tri 45670 32250 45960 32540 ne
rect 45960 32514 49680 32540
tri 49680 32514 49940 32774 sw
tri 49974 32514 50234 32774 ne
rect 50234 32514 70613 32774
rect 45960 32250 49940 32514
rect 43978 31962 45670 32250
rect 41725 31946 43689 31962
rect 37408 31722 41428 31946
rect 33044 31624 37126 31722
tri 37126 31624 37224 31722 sw
tri 37408 31624 37506 31722 ne
rect 37506 31649 41428 31722
tri 41428 31649 41725 31946 sw
tri 41725 31649 42022 31946 ne
rect 42022 31673 43689 31946
tri 43689 31673 43978 31962 sw
tri 43978 31673 44267 31962 ne
rect 44267 31960 45670 31962
tri 45670 31960 45960 32250 sw
tri 45960 31960 46250 32250 ne
rect 46250 32220 49940 32250
tri 49940 32220 50234 32514 sw
tri 50234 32220 50528 32514 ne
rect 50528 32220 70613 32514
rect 46250 31960 50234 32220
rect 44267 31914 45960 31960
tri 45960 31914 46006 31960 sw
tri 46250 31914 46296 31960 ne
rect 46296 31926 50234 31960
tri 50234 31926 50528 32220 sw
tri 50528 31926 50822 32220 ne
rect 50822 31926 70613 32220
rect 46296 31914 50528 31926
rect 44267 31673 46006 31914
rect 42022 31649 43978 31673
rect 37506 31624 41725 31649
rect 33044 31560 37224 31624
rect 29092 31268 32752 31560
tri 32752 31268 33044 31560 sw
tri 33044 31268 33336 31560 ne
rect 33336 31342 37224 31560
tri 37224 31342 37506 31624 sw
tri 37506 31342 37788 31624 ne
rect 37788 31534 41725 31624
tri 41725 31534 41840 31649 sw
tri 42022 31534 42137 31649 ne
rect 42137 31534 43978 31649
rect 37788 31342 41840 31534
rect 33336 31268 37506 31342
rect 29092 30976 33044 31268
tri 33044 30976 33336 31268 sw
tri 33336 30976 33628 31268 ne
rect 33628 31060 37506 31268
tri 37506 31060 37788 31342 sw
tri 37788 31060 38070 31342 ne
rect 38070 31237 41840 31342
tri 41840 31237 42137 31534 sw
tri 42137 31237 42434 31534 ne
rect 42434 31518 43978 31534
tri 43978 31518 44133 31673 sw
tri 44267 31518 44422 31673 ne
rect 44422 31624 46006 31673
tri 46006 31624 46296 31914 sw
tri 46296 31624 46586 31914 ne
rect 46586 31632 50528 31914
tri 50528 31632 50822 31926 sw
tri 50822 31632 51116 31926 ne
rect 51116 31632 70613 31926
rect 46586 31624 50822 31632
rect 44422 31518 46296 31624
rect 42434 31237 44133 31518
rect 38070 31060 42137 31237
rect 33628 30976 37788 31060
tri 29092 26732 33336 30976 ne
tri 33336 30684 33628 30976 sw
tri 33628 30684 33920 30976 ne
rect 33920 30778 37788 30976
tri 37788 30778 38070 31060 sw
tri 38070 30778 38352 31060 ne
rect 38352 30940 42137 31060
tri 42137 30940 42434 31237 sw
tri 42434 30940 42731 31237 ne
rect 42731 31229 44133 31237
tri 44133 31229 44422 31518 sw
tri 44422 31229 44711 31518 ne
rect 44711 31334 46296 31518
tri 46296 31334 46586 31624 sw
tri 46586 31334 46876 31624 ne
rect 46876 31338 50822 31624
tri 50822 31338 51116 31632 sw
tri 51116 31338 51410 31632 ne
rect 51410 31338 70613 31632
rect 46876 31334 51116 31338
rect 44711 31229 46586 31334
rect 42731 30940 44422 31229
tri 44422 30940 44711 31229 sw
tri 44711 30940 45000 31229 ne
rect 45000 31044 46586 31229
tri 46586 31044 46876 31334 sw
tri 46876 31044 47166 31334 ne
rect 47166 31044 51116 31334
tri 51116 31044 51410 31338 sw
tri 51410 31044 51704 31338 ne
rect 51704 31044 70613 31338
rect 45000 30940 46876 31044
rect 38352 30778 42434 30940
rect 33920 30684 38070 30778
rect 33336 30392 33628 30684
tri 33628 30392 33920 30684 sw
tri 33920 30392 34212 30684 ne
rect 34212 30496 38070 30684
tri 38070 30496 38352 30778 sw
tri 38352 30496 38634 30778 ne
rect 38634 30643 42434 30778
tri 42434 30643 42731 30940 sw
tri 42731 30643 43028 30940 ne
rect 43028 30849 44711 30940
tri 44711 30849 44802 30940 sw
tri 45000 30849 45091 30940 ne
rect 45091 30849 46876 30940
rect 43028 30643 44802 30849
rect 38634 30560 42731 30643
tri 42731 30560 42814 30643 sw
tri 43028 30560 43111 30643 ne
rect 43111 30560 44802 30643
tri 44802 30560 45091 30849 sw
tri 45091 30560 45380 30849 ne
rect 45380 30754 46876 30849
tri 46876 30754 47166 31044 sw
tri 47166 30754 47456 31044 ne
rect 47456 30754 51410 31044
rect 45380 30560 47166 30754
rect 38634 30496 42814 30560
rect 34212 30392 38352 30496
rect 33336 30100 33920 30392
tri 33920 30100 34212 30392 sw
tri 34212 30100 34504 30392 ne
rect 34504 30214 38352 30392
tri 38352 30214 38634 30496 sw
tri 38634 30214 38916 30496 ne
rect 38916 30263 42814 30496
tri 42814 30263 43111 30560 sw
tri 43111 30263 43408 30560 ne
rect 43408 30271 45091 30560
tri 45091 30271 45380 30560 sw
tri 45380 30271 45669 30560 ne
rect 45669 30464 47166 30560
tri 47166 30464 47456 30754 sw
tri 47456 30464 47746 30754 ne
rect 47746 30750 51410 30754
tri 51410 30750 51704 31044 sw
tri 51704 30750 51998 31044 ne
rect 51998 30750 70613 31044
rect 47746 30464 51704 30750
rect 45669 30290 47456 30464
tri 47456 30290 47630 30464 sw
tri 47746 30290 47920 30464 ne
rect 47920 30456 51704 30464
tri 51704 30456 51998 30750 sw
tri 51998 30456 52292 30750 ne
rect 52292 30456 70613 30750
rect 47920 30388 51998 30456
tri 51998 30388 52066 30456 sw
tri 52292 30388 52360 30456 ne
rect 52360 30388 70613 30456
rect 47920 30290 52066 30388
rect 45669 30271 47630 30290
rect 43408 30263 45380 30271
rect 38916 30214 43111 30263
rect 34504 30100 38634 30214
rect 33336 29808 34212 30100
tri 34212 29808 34504 30100 sw
tri 34504 29808 34796 30100 ne
rect 34796 29932 38634 30100
tri 38634 29932 38916 30214 sw
tri 38916 29932 39198 30214 ne
rect 39198 29966 43111 30214
tri 43111 29966 43408 30263 sw
tri 43408 29966 43705 30263 ne
rect 43705 29982 45380 30263
tri 45380 29982 45669 30271 sw
tri 45669 29982 45958 30271 ne
rect 45958 30000 47630 30271
tri 47630 30000 47920 30290 sw
tri 47920 30000 48210 30290 ne
rect 48210 30094 52066 30290
tri 52066 30094 52360 30388 sw
tri 52360 30094 52654 30388 ne
rect 52654 30094 70613 30388
rect 48210 30000 52360 30094
rect 45958 29982 47920 30000
rect 43705 29966 45669 29982
rect 39198 29932 43408 29966
rect 34796 29808 38916 29932
rect 33336 29764 34504 29808
tri 34504 29764 34548 29808 sw
tri 34796 29764 34840 29808 ne
rect 34840 29764 38916 29808
rect 33336 29472 34548 29764
tri 34548 29472 34840 29764 sw
tri 34840 29472 35132 29764 ne
rect 35132 29650 38916 29764
tri 38916 29650 39198 29932 sw
tri 39198 29650 39480 29932 ne
rect 39480 29779 43408 29932
tri 43408 29779 43595 29966 sw
tri 43705 29779 43892 29966 ne
rect 43892 29779 45669 29966
rect 39480 29650 43595 29779
rect 35132 29472 39198 29650
rect 33336 29180 34840 29472
tri 34840 29180 35132 29472 sw
tri 35132 29180 35424 29472 ne
rect 35424 29368 39198 29472
tri 39198 29368 39480 29650 sw
tri 39480 29368 39762 29650 ne
rect 39762 29482 43595 29650
tri 43595 29482 43892 29779 sw
tri 43892 29482 44189 29779 ne
rect 44189 29693 45669 29779
tri 45669 29693 45958 29982 sw
tri 45958 29693 46247 29982 ne
rect 46247 29710 47920 29982
tri 47920 29710 48210 30000 sw
tri 48210 29710 48500 30000 ne
rect 48500 29800 52360 30000
tri 52360 29800 52654 30094 sw
tri 52654 30000 52748 30094 ne
rect 52748 30056 70613 30094
rect 70669 30056 71000 32920
rect 52748 30000 71000 30056
rect 48500 29752 71000 29800
rect 48500 29710 70613 29752
rect 46247 29693 48210 29710
rect 44189 29538 45958 29693
tri 45958 29538 46113 29693 sw
tri 46247 29538 46402 29693 ne
rect 46402 29538 48210 29693
rect 44189 29482 46113 29538
rect 39762 29368 43892 29482
rect 35424 29180 39480 29368
rect 33336 28888 35132 29180
tri 35132 28888 35424 29180 sw
tri 35424 28888 35716 29180 ne
rect 35716 29170 39480 29180
tri 39480 29170 39678 29368 sw
tri 39762 29170 39960 29368 ne
rect 39960 29185 43892 29368
tri 43892 29185 44189 29482 sw
tri 44189 29185 44486 29482 ne
rect 44486 29249 46113 29482
tri 46113 29249 46402 29538 sw
tri 46402 29249 46691 29538 ne
rect 46691 29420 48210 29538
tri 48210 29420 48500 29710 sw
tri 48500 29420 48790 29710 ne
rect 48790 29420 70613 29710
rect 46691 29249 48500 29420
rect 44486 29185 46402 29249
rect 39960 29170 44189 29185
rect 35716 28888 39678 29170
tri 39678 28888 39960 29170 sw
tri 39960 28888 40242 29170 ne
rect 40242 28888 44189 29170
tri 44189 28888 44486 29185 sw
tri 44486 28888 44783 29185 ne
rect 44783 28960 46402 29185
tri 46402 28960 46691 29249 sw
tri 46691 28960 46980 29249 ne
rect 46980 29160 48500 29249
tri 48500 29160 48760 29420 sw
tri 48790 29160 49050 29420 ne
rect 49050 29160 70613 29420
rect 46980 28960 48760 29160
rect 44783 28888 46691 28960
rect 33336 28596 35424 28888
tri 35424 28596 35716 28888 sw
tri 35716 28596 36008 28888 ne
rect 36008 28606 39960 28888
tri 39960 28606 40242 28888 sw
tri 40242 28606 40524 28888 ne
rect 40524 28606 44486 28888
rect 36008 28596 40242 28606
rect 33336 28304 35716 28596
tri 35716 28304 36008 28596 sw
tri 36008 28304 36300 28596 ne
rect 36300 28324 40242 28596
tri 40242 28324 40524 28606 sw
tri 40524 28324 40806 28606 ne
rect 40806 28591 44486 28606
tri 44486 28591 44783 28888 sw
tri 44783 28591 45080 28888 ne
rect 45080 28869 46691 28888
tri 46691 28869 46782 28960 sw
tri 46980 28869 47071 28960 ne
rect 47071 28870 48760 28960
tri 48760 28870 49050 29160 sw
tri 49050 28870 49340 29160 ne
rect 49340 28870 70613 29160
rect 47071 28869 49050 28870
rect 45080 28591 46782 28869
rect 40806 28580 44783 28591
tri 44783 28580 44794 28591 sw
tri 45080 28580 45091 28591 ne
rect 45091 28580 46782 28591
tri 46782 28580 47071 28869 sw
tri 47071 28580 47360 28869 ne
rect 47360 28580 49050 28869
tri 49050 28580 49340 28870 sw
tri 49340 28580 49630 28870 ne
rect 49630 28580 70613 28870
rect 40806 28324 44794 28580
rect 36300 28304 40524 28324
rect 33336 28012 36008 28304
tri 36008 28012 36300 28304 sw
tri 36300 28012 36592 28304 ne
rect 36592 28042 40524 28304
tri 40524 28042 40806 28324 sw
tri 40806 28042 41088 28324 ne
rect 41088 28283 44794 28324
tri 44794 28283 45091 28580 sw
tri 45091 28283 45388 28580 ne
rect 45388 28291 47071 28580
tri 47071 28291 47360 28580 sw
tri 47360 28291 47649 28580 ne
rect 47649 28291 49340 28580
rect 45388 28283 47360 28291
rect 41088 28042 45091 28283
rect 36592 28012 40806 28042
rect 33336 27900 36300 28012
tri 36300 27900 36412 28012 sw
tri 36592 27900 36704 28012 ne
rect 36704 27900 40806 28012
rect 33336 27608 36412 27900
tri 36412 27608 36704 27900 sw
tri 36704 27608 36996 27900 ne
rect 36996 27760 40806 27900
tri 40806 27760 41088 28042 sw
tri 41088 27760 41370 28042 ne
rect 41370 27986 45091 28042
tri 45091 27986 45388 28283 sw
tri 45388 27986 45685 28283 ne
rect 45685 28002 47360 28283
tri 47360 28002 47649 28291 sw
tri 47649 28002 47938 28291 ne
rect 47938 28290 49340 28291
tri 49340 28290 49630 28580 sw
tri 49630 28290 49920 28580 ne
rect 49920 28290 70613 28580
rect 47938 28002 49630 28290
rect 45685 27986 47649 28002
rect 41370 27760 45388 27986
rect 36996 27608 41088 27760
rect 33336 27316 36704 27608
tri 36704 27316 36996 27608 sw
tri 36996 27316 37288 27608 ne
rect 37288 27478 41088 27608
tri 41088 27478 41370 27760 sw
tri 41370 27478 41652 27760 ne
rect 41652 27689 45388 27760
tri 45388 27689 45685 27986 sw
tri 45685 27689 45982 27986 ne
rect 45982 27713 47649 27986
tri 47649 27713 47938 28002 sw
tri 47938 27713 48227 28002 ne
rect 48227 28000 49630 28002
tri 49630 28000 49920 28290 sw
tri 49920 28000 50210 28290 ne
rect 50210 28000 70613 28290
rect 48227 27713 49920 28000
rect 45982 27689 47938 27713
rect 41652 27574 45685 27689
tri 45685 27574 45800 27689 sw
tri 45982 27574 46097 27689 ne
rect 46097 27574 47938 27689
rect 41652 27478 45800 27574
rect 37288 27380 41370 27478
tri 41370 27380 41468 27478 sw
tri 41652 27380 41750 27478 ne
rect 41750 27380 45800 27478
rect 37288 27316 41468 27380
rect 33336 27024 36996 27316
tri 36996 27024 37288 27316 sw
tri 37288 27024 37580 27316 ne
rect 37580 27098 41468 27316
tri 41468 27098 41750 27380 sw
tri 41750 27098 42032 27380 ne
rect 42032 27277 45800 27380
tri 45800 27277 46097 27574 sw
tri 46097 27277 46394 27574 ne
rect 46394 27558 47938 27574
tri 47938 27558 48093 27713 sw
tri 48227 27558 48382 27713 ne
rect 48382 27710 49920 27713
tri 49920 27710 50210 28000 sw
tri 50210 27710 50500 28000 ne
rect 50500 27710 70613 28000
rect 48382 27670 50210 27710
tri 50210 27670 50250 27710 sw
tri 50500 27670 50540 27710 ne
rect 50540 27670 70613 27710
rect 48382 27558 50250 27670
rect 46394 27277 48093 27558
rect 42032 27098 46097 27277
rect 37580 27024 41750 27098
rect 33336 26732 37288 27024
tri 37288 26732 37580 27024 sw
tri 37580 26732 37872 27024 ne
rect 37872 26816 41750 27024
tri 41750 26816 42032 27098 sw
tri 42032 26816 42314 27098 ne
rect 42314 26980 46097 27098
tri 46097 26980 46394 27277 sw
tri 46394 26980 46691 27277 ne
rect 46691 27269 48093 27277
tri 48093 27269 48382 27558 sw
tri 48382 27269 48671 27558 ne
rect 48671 27380 50250 27558
tri 50250 27380 50540 27670 sw
tri 50540 27380 50830 27670 ne
rect 50830 27380 70613 27670
rect 48671 27269 50540 27380
rect 46691 26980 48382 27269
tri 48382 26980 48671 27269 sw
tri 48671 26980 48960 27269 ne
rect 48960 27090 50540 27269
tri 50540 27090 50830 27380 sw
tri 50830 27090 51120 27380 ne
rect 51120 27090 70613 27380
rect 48960 26980 50830 27090
rect 42314 26816 46394 26980
rect 37872 26732 42032 26816
tri 33336 22488 37580 26732 ne
tri 37580 26440 37872 26732 sw
tri 37872 26440 38164 26732 ne
rect 38164 26534 42032 26732
tri 42032 26534 42314 26816 sw
tri 42314 26534 42596 26816 ne
rect 42596 26683 46394 26816
tri 46394 26683 46691 26980 sw
tri 46691 26683 46988 26980 ne
rect 46988 26800 48671 26980
tri 48671 26800 48851 26980 sw
tri 48960 26800 49140 26980 ne
rect 49140 26800 50830 26980
tri 50830 26800 51120 27090 sw
tri 51120 26800 51410 27090 ne
rect 51410 26888 70613 27090
rect 70669 26888 71000 29752
rect 51410 26800 71000 26888
rect 46988 26683 48851 26800
rect 42596 26600 46691 26683
tri 46691 26600 46774 26683 sw
tri 46988 26600 47071 26683 ne
rect 47071 26600 48851 26683
tri 48851 26600 49051 26800 sw
tri 49140 26600 49340 26800 ne
rect 49340 26600 51120 26800
tri 51120 26600 51320 26800 sw
rect 42596 26534 46774 26600
rect 38164 26440 42314 26534
rect 37580 26148 37872 26440
tri 37872 26148 38164 26440 sw
tri 38164 26148 38456 26440 ne
rect 38456 26252 42314 26440
tri 42314 26252 42596 26534 sw
tri 42596 26252 42878 26534 ne
rect 42878 26303 46774 26534
tri 46774 26303 47071 26600 sw
tri 47071 26303 47368 26600 ne
rect 47368 26311 49051 26600
tri 49051 26311 49340 26600 sw
tri 49340 26311 49629 26600 ne
rect 49629 26311 71000 26600
rect 47368 26303 49340 26311
rect 42878 26252 47071 26303
rect 38456 26148 42596 26252
rect 37580 25856 38164 26148
tri 38164 25856 38456 26148 sw
tri 38456 25856 38748 26148 ne
rect 38748 25970 42596 26148
tri 42596 25970 42878 26252 sw
tri 42878 25970 43160 26252 ne
rect 43160 26006 47071 26252
tri 47071 26006 47368 26303 sw
tri 47368 26006 47665 26303 ne
rect 47665 26022 49340 26303
tri 49340 26022 49629 26311 sw
tri 49629 26022 49918 26311 ne
rect 49918 26022 71000 26311
rect 47665 26006 49629 26022
rect 43160 25970 47368 26006
rect 38748 25856 42878 25970
rect 37580 25564 38456 25856
tri 38456 25564 38748 25856 sw
tri 38748 25564 39040 25856 ne
rect 39040 25688 42878 25856
tri 42878 25688 43160 25970 sw
tri 43160 25688 43442 25970 ne
rect 43442 25709 47368 25970
tri 47368 25709 47665 26006 sw
tri 47665 25709 47962 26006 ne
rect 47962 25778 49629 26006
tri 49629 25778 49873 26022 sw
tri 49918 25778 50162 26022 ne
rect 50162 25778 71000 26022
rect 47962 25709 49873 25778
rect 43442 25688 47665 25709
rect 39040 25564 43160 25688
rect 37580 25520 38748 25564
tri 38748 25520 38792 25564 sw
tri 39040 25520 39084 25564 ne
rect 39084 25520 43160 25564
rect 37580 25228 38792 25520
tri 38792 25228 39084 25520 sw
tri 39084 25228 39376 25520 ne
rect 39376 25406 43160 25520
tri 43160 25406 43442 25688 sw
tri 43442 25406 43724 25688 ne
rect 43724 25594 47665 25688
tri 47665 25594 47780 25709 sw
tri 47962 25594 48077 25709 ne
rect 48077 25594 49873 25709
rect 43724 25406 47780 25594
rect 39376 25228 43442 25406
rect 37580 24936 39084 25228
tri 39084 24936 39376 25228 sw
tri 39376 24936 39668 25228 ne
rect 39668 25124 43442 25228
tri 43442 25124 43724 25406 sw
tri 43724 25124 44006 25406 ne
rect 44006 25297 47780 25406
tri 47780 25297 48077 25594 sw
tri 48077 25297 48374 25594 ne
rect 48374 25489 49873 25594
tri 49873 25489 50162 25778 sw
tri 50162 25489 50451 25778 ne
rect 50451 25489 71000 25778
rect 48374 25297 50162 25489
rect 44006 25124 48077 25297
rect 39668 24936 43724 25124
rect 37580 24644 39376 24936
tri 39376 24644 39668 24936 sw
tri 39668 24644 39960 24936 ne
rect 39960 24926 43724 24936
tri 43724 24926 43922 25124 sw
tri 44006 24926 44204 25124 ne
rect 44204 25000 48077 25124
tri 48077 25000 48374 25297 sw
tri 48374 25000 48671 25297 ne
rect 48671 25200 50162 25297
tri 50162 25200 50451 25489 sw
tri 50451 25200 50740 25489 ne
rect 50740 25200 71000 25489
rect 48671 25000 50451 25200
tri 50451 25000 50651 25200 sw
rect 44204 24941 48374 25000
tri 48374 24941 48433 25000 sw
tri 48671 24941 48730 25000 ne
rect 48730 24941 71000 25000
rect 44204 24926 48433 24941
rect 39960 24644 43922 24926
tri 43922 24644 44204 24926 sw
tri 44204 24644 44486 24926 ne
rect 44486 24644 48433 24926
tri 48433 24644 48730 24941 sw
tri 48730 24644 49027 24941 ne
rect 49027 24906 71000 24941
rect 49027 24644 70613 24906
rect 37580 24352 39668 24644
tri 39668 24352 39960 24644 sw
tri 39960 24352 40252 24644 ne
rect 40252 24362 44204 24644
tri 44204 24362 44486 24644 sw
tri 44486 24362 44768 24644 ne
rect 44768 24362 48730 24644
rect 40252 24352 44486 24362
rect 37580 24060 39960 24352
tri 39960 24060 40252 24352 sw
tri 40252 24060 40544 24352 ne
rect 40544 24080 44486 24352
tri 44486 24080 44768 24362 sw
tri 44768 24080 45050 24362 ne
rect 45050 24347 48730 24362
tri 48730 24347 49027 24644 sw
tri 49027 24347 49324 24644 ne
rect 49324 24347 70613 24644
rect 45050 24080 49027 24347
rect 40544 24060 44768 24080
rect 37580 23768 40252 24060
tri 40252 23768 40544 24060 sw
tri 40544 23768 40836 24060 ne
rect 40836 23798 44768 24060
tri 44768 23798 45050 24080 sw
tri 45050 23798 45332 24080 ne
rect 45332 24050 49027 24080
tri 49027 24050 49324 24347 sw
tri 49324 24050 49621 24347 ne
rect 49621 24050 70613 24347
rect 45332 23994 49324 24050
tri 49324 23994 49380 24050 sw
tri 49621 23994 49677 24050 ne
rect 49677 23994 70613 24050
rect 45332 23798 49380 23994
rect 40836 23768 45050 23798
rect 37580 23656 40544 23768
tri 40544 23656 40656 23768 sw
tri 40836 23656 40948 23768 ne
rect 40948 23656 45050 23768
rect 37580 23364 40656 23656
tri 40656 23364 40948 23656 sw
tri 40948 23364 41240 23656 ne
rect 41240 23516 45050 23656
tri 45050 23516 45332 23798 sw
tri 45332 23516 45614 23798 ne
rect 45614 23697 49380 23798
tri 49380 23697 49677 23994 sw
tri 49677 23697 49974 23994 ne
rect 49974 23706 70613 23994
rect 70669 23706 71000 24906
rect 49974 23697 71000 23706
rect 45614 23516 49677 23697
rect 41240 23364 45332 23516
rect 37580 23072 40948 23364
tri 40948 23072 41240 23364 sw
tri 41240 23072 41532 23364 ne
rect 41532 23234 45332 23364
tri 45332 23234 45614 23516 sw
tri 45614 23234 45896 23516 ne
rect 45896 23400 49677 23516
tri 49677 23400 49974 23697 sw
tri 49974 23600 50071 23697 ne
rect 50071 23600 71000 23697
rect 45896 23234 71000 23400
rect 41532 23136 45614 23234
tri 45614 23136 45712 23234 sw
tri 45896 23136 45994 23234 ne
rect 45994 23136 71000 23234
rect 41532 23072 45712 23136
rect 37580 22780 41240 23072
tri 41240 22780 41532 23072 sw
tri 41532 22780 41824 23072 ne
rect 41824 22854 45712 23072
tri 45712 22854 45994 23136 sw
tri 45994 22854 46276 23136 ne
rect 46276 22854 71000 23136
rect 41824 22780 45994 22854
rect 37580 22488 41532 22780
tri 41532 22488 41824 22780 sw
tri 41824 22488 42116 22780 ne
rect 42116 22572 45994 22780
tri 45994 22572 46276 22854 sw
tri 46276 22572 46558 22854 ne
rect 46558 22572 71000 22854
rect 42116 22488 46276 22572
tri 37580 18244 41824 22488 ne
tri 41824 22196 42116 22488 sw
tri 42116 22196 42408 22488 ne
rect 42408 22290 46276 22488
tri 46276 22290 46558 22572 sw
tri 46558 22290 46840 22572 ne
rect 46840 22290 71000 22572
rect 42408 22196 46558 22290
rect 41824 21904 42116 22196
tri 42116 21904 42408 22196 sw
tri 42408 21904 42700 22196 ne
rect 42700 22008 46558 22196
tri 46558 22008 46840 22290 sw
tri 46840 22008 47122 22290 ne
rect 47122 22008 71000 22290
rect 42700 21904 46840 22008
rect 41824 21612 42408 21904
tri 42408 21612 42700 21904 sw
tri 42700 21612 42992 21904 ne
rect 42992 21726 46840 21904
tri 46840 21726 47122 22008 sw
tri 47122 21726 47404 22008 ne
rect 47404 21726 71000 22008
rect 42992 21612 47122 21726
rect 41824 21320 42700 21612
tri 42700 21320 42992 21612 sw
tri 42992 21320 43284 21612 ne
rect 43284 21444 47122 21612
tri 47122 21444 47404 21726 sw
tri 47404 21444 47686 21726 ne
rect 47686 21444 71000 21726
rect 43284 21320 47404 21444
rect 41824 21276 42992 21320
tri 42992 21276 43036 21320 sw
tri 43284 21276 43328 21320 ne
rect 43328 21276 47404 21320
rect 41824 20984 43036 21276
tri 43036 20984 43328 21276 sw
tri 43328 20984 43620 21276 ne
rect 43620 21162 47404 21276
tri 47404 21162 47686 21444 sw
tri 47686 21162 47968 21444 ne
rect 47968 21162 71000 21444
rect 43620 20984 47686 21162
rect 41824 20692 43328 20984
tri 43328 20692 43620 20984 sw
tri 43620 20692 43912 20984 ne
rect 43912 20880 47686 20984
tri 47686 20880 47968 21162 sw
tri 47968 20880 48250 21162 ne
rect 48250 20880 71000 21162
rect 43912 20764 47968 20880
tri 47968 20764 48084 20880 sw
tri 48250 20764 48366 20880 ne
rect 48366 20764 71000 20880
rect 43912 20692 48084 20764
rect 41824 20400 43620 20692
tri 43620 20400 43912 20692 sw
tri 43912 20400 44204 20692 ne
rect 44204 20482 48084 20692
tri 48084 20482 48366 20764 sw
tri 48366 20482 48648 20764 ne
rect 48648 20482 71000 20764
rect 44204 20400 48366 20482
rect 41824 20108 43912 20400
tri 43912 20108 44204 20400 sw
tri 44204 20108 44496 20400 ne
rect 44496 20200 48366 20400
tri 48366 20200 48648 20482 sw
tri 48648 20400 48730 20482 ne
rect 48730 20400 71000 20482
rect 44496 20108 71000 20200
rect 41824 19816 44204 20108
tri 44204 19816 44496 20108 sw
tri 44496 19816 44788 20108 ne
rect 44788 19816 71000 20108
rect 41824 19524 44496 19816
tri 44496 19524 44788 19816 sw
tri 44788 19524 45080 19816 ne
rect 45080 19524 71000 19816
rect 41824 19412 44788 19524
tri 44788 19412 44900 19524 sw
tri 45080 19412 45192 19524 ne
rect 45192 19412 71000 19524
rect 41824 19120 44900 19412
tri 44900 19120 45192 19412 sw
tri 45192 19120 45484 19412 ne
rect 45484 19120 71000 19412
rect 41824 18828 45192 19120
tri 45192 18828 45484 19120 sw
tri 45484 18828 45776 19120 ne
rect 45776 18828 71000 19120
rect 41824 18536 45484 18828
tri 45484 18536 45776 18828 sw
tri 45776 18536 46068 18828 ne
rect 46068 18536 71000 18828
rect 41824 18244 45776 18536
tri 45776 18244 46068 18536 sw
tri 46068 18244 46360 18536 ne
rect 46360 18244 71000 18536
tri 41824 14000 46068 18244 ne
tri 46068 17952 46360 18244 sw
tri 46360 17952 46652 18244 ne
rect 46652 17952 71000 18244
rect 46068 17660 46360 17952
tri 46360 17660 46652 17952 sw
tri 46652 17660 46944 17952 ne
rect 46944 17660 71000 17952
rect 46068 17584 46652 17660
tri 46652 17584 46728 17660 sw
tri 46944 17584 47020 17660 ne
rect 47020 17584 71000 17660
rect 46068 17292 46728 17584
tri 46728 17292 47020 17584 sw
tri 47020 17292 47312 17584 ne
rect 47312 17292 71000 17584
rect 46068 17000 47020 17292
tri 47020 17000 47312 17292 sw
tri 47312 17200 47404 17292 ne
rect 47404 17200 71000 17292
rect 46068 14000 71000 17000
use M1_PSUB_CDNS_40661953145669  M1_PSUB_CDNS_40661953145669_0
timestamp 1755005639
transform -1 0 58007 0 -1 13194
box 0 0 1 1
use M1_PSUB_CDNS_40661953145670  M1_PSUB_CDNS_40661953145670_0
timestamp 1755005639
transform 0 -1 69871 1 0 70385
box 0 0 1 1
use M1_PSUB_CDNS_40661953145671  M1_PSUB_CDNS_40661953145671_0
timestamp 1755005639
transform 1 0 70235 0 1 69871
box 0 0 1 1
use M1_PSUB_CDNS_40661953145672  M1_PSUB_CDNS_40661953145672_0
timestamp 1755005639
transform 0 -1 70899 1 0 41649
box 0 0 1 1
use M1_PSUB_CDNS_40661953145672  M1_PSUB_CDNS_40661953145672_1
timestamp 1755005639
transform 1 0 41636 0 1 70900
box 0 0 1 1
use M1_PSUB_CDNS_40661953145673  M1_PSUB_CDNS_40661953145673_0
timestamp 1755005639
transform 0 -1 13194 1 0 58004
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_0
timestamp 1755005639
transform 1 0 42317 0 1 15761
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_1
timestamp 1755005639
transform 1 0 42185 0 1 15893
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_2
timestamp 1755005639
transform 1 0 42977 0 1 15101
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_3
timestamp 1755005639
transform 1 0 44873 0 1 13233
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_4
timestamp 1755005639
transform 1 0 44693 0 1 13385
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_5
timestamp 1755005639
transform 1 0 44561 0 1 13517
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_6
timestamp 1755005639
transform 1 0 44429 0 1 13649
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_7
timestamp 1755005639
transform 1 0 44297 0 1 13781
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_8
timestamp 1755005639
transform 1 0 44165 0 1 13913
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_9
timestamp 1755005639
transform 1 0 44033 0 1 14045
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_10
timestamp 1755005639
transform 1 0 43901 0 1 14177
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_11
timestamp 1755005639
transform 1 0 43769 0 1 14309
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_12
timestamp 1755005639
transform 1 0 43637 0 1 14441
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_13
timestamp 1755005639
transform 1 0 43505 0 1 14573
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_14
timestamp 1755005639
transform 1 0 43373 0 1 14705
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_15
timestamp 1755005639
transform 1 0 43241 0 1 14837
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_16
timestamp 1755005639
transform 1 0 43109 0 1 14969
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_17
timestamp 1755005639
transform 1 0 42845 0 1 15233
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_18
timestamp 1755005639
transform 1 0 42713 0 1 15365
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_19
timestamp 1755005639
transform 1 0 42581 0 1 15497
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_20
timestamp 1755005639
transform 1 0 42449 0 1 15629
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_21
timestamp 1755005639
transform 1 0 33605 0 1 24473
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_22
timestamp 1755005639
transform 1 0 39017 0 1 19061
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_23
timestamp 1755005639
transform 1 0 38885 0 1 19193
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_24
timestamp 1755005639
transform 1 0 38753 0 1 19325
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_25
timestamp 1755005639
transform 1 0 38621 0 1 19457
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_26
timestamp 1755005639
transform 1 0 38489 0 1 19589
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_27
timestamp 1755005639
transform 1 0 38357 0 1 19721
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_28
timestamp 1755005639
transform 1 0 33737 0 1 24341
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_29
timestamp 1755005639
transform 1 0 33869 0 1 24209
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_30
timestamp 1755005639
transform 1 0 34001 0 1 24077
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_31
timestamp 1755005639
transform 1 0 34133 0 1 23945
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_32
timestamp 1755005639
transform 1 0 34265 0 1 23813
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_33
timestamp 1755005639
transform 1 0 34397 0 1 23681
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_34
timestamp 1755005639
transform 1 0 34529 0 1 23549
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_35
timestamp 1755005639
transform 1 0 34661 0 1 23417
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_36
timestamp 1755005639
transform 1 0 34793 0 1 23285
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_37
timestamp 1755005639
transform 1 0 33209 0 1 24869
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_38
timestamp 1755005639
transform 1 0 39413 0 1 18665
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_39
timestamp 1755005639
transform 1 0 41261 0 1 16817
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_40
timestamp 1755005639
transform 1 0 36245 0 1 21833
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_41
timestamp 1755005639
transform 1 0 37301 0 1 20777
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_42
timestamp 1755005639
transform 1 0 37169 0 1 20909
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_43
timestamp 1755005639
transform 1 0 37037 0 1 21041
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_44
timestamp 1755005639
transform 1 0 36905 0 1 21173
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_45
timestamp 1755005639
transform 1 0 36773 0 1 21305
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_46
timestamp 1755005639
transform 1 0 36641 0 1 21437
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_47
timestamp 1755005639
transform 1 0 36509 0 1 21569
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_48
timestamp 1755005639
transform 1 0 36377 0 1 21701
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_49
timestamp 1755005639
transform 1 0 32945 0 1 25133
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_50
timestamp 1755005639
transform 1 0 32813 0 1 25265
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_51
timestamp 1755005639
transform 1 0 32681 0 1 25397
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_52
timestamp 1755005639
transform 1 0 32549 0 1 25529
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_53
timestamp 1755005639
transform 1 0 32417 0 1 25661
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_54
timestamp 1755005639
transform 1 0 32285 0 1 25793
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_55
timestamp 1755005639
transform 1 0 32153 0 1 25925
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_56
timestamp 1755005639
transform 1 0 32021 0 1 26057
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_57
timestamp 1755005639
transform 1 0 31889 0 1 26189
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_58
timestamp 1755005639
transform 1 0 31757 0 1 26321
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_59
timestamp 1755005639
transform 1 0 31625 0 1 26453
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_60
timestamp 1755005639
transform 1 0 31493 0 1 26585
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_61
timestamp 1755005639
transform 1 0 31361 0 1 26717
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_62
timestamp 1755005639
transform 1 0 31229 0 1 26849
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_63
timestamp 1755005639
transform 1 0 33077 0 1 25001
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_64
timestamp 1755005639
transform 1 0 30965 0 1 27113
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_65
timestamp 1755005639
transform 1 0 30833 0 1 27245
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_66
timestamp 1755005639
transform 1 0 30701 0 1 27377
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_67
timestamp 1755005639
transform 1 0 31097 0 1 26981
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_68
timestamp 1755005639
transform 1 0 36113 0 1 21965
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_69
timestamp 1755005639
transform 1 0 35981 0 1 22097
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_70
timestamp 1755005639
transform 1 0 35849 0 1 22229
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_71
timestamp 1755005639
transform 1 0 35717 0 1 22361
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_72
timestamp 1755005639
transform 1 0 35585 0 1 22493
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_73
timestamp 1755005639
transform 1 0 35453 0 1 22625
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_74
timestamp 1755005639
transform 1 0 35321 0 1 22757
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_75
timestamp 1755005639
transform 1 0 35189 0 1 22889
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_76
timestamp 1755005639
transform 1 0 34925 0 1 23153
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_77
timestamp 1755005639
transform 1 0 41921 0 1 16157
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_78
timestamp 1755005639
transform 1 0 41789 0 1 16289
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_79
timestamp 1755005639
transform 1 0 41657 0 1 16421
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_80
timestamp 1755005639
transform 1 0 41525 0 1 16553
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_81
timestamp 1755005639
transform 1 0 41393 0 1 16685
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_82
timestamp 1755005639
transform 1 0 39281 0 1 18797
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_83
timestamp 1755005639
transform 1 0 41129 0 1 16949
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_84
timestamp 1755005639
transform 1 0 40997 0 1 17081
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_85
timestamp 1755005639
transform 1 0 40865 0 1 17213
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_86
timestamp 1755005639
transform 1 0 40733 0 1 17345
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_87
timestamp 1755005639
transform 1 0 40601 0 1 17477
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_88
timestamp 1755005639
transform 1 0 40469 0 1 17609
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_89
timestamp 1755005639
transform 1 0 40337 0 1 17741
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_90
timestamp 1755005639
transform 1 0 40205 0 1 17873
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_91
timestamp 1755005639
transform 1 0 40073 0 1 18005
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_92
timestamp 1755005639
transform 1 0 39941 0 1 18137
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_93
timestamp 1755005639
transform 1 0 39809 0 1 18269
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_94
timestamp 1755005639
transform 1 0 39677 0 1 18401
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_95
timestamp 1755005639
transform 1 0 38225 0 1 19853
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_96
timestamp 1755005639
transform 1 0 38093 0 1 19985
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_97
timestamp 1755005639
transform 1 0 37961 0 1 20117
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_98
timestamp 1755005639
transform 1 0 37829 0 1 20249
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_99
timestamp 1755005639
transform 1 0 37697 0 1 20381
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_100
timestamp 1755005639
transform 1 0 37565 0 1 20513
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_101
timestamp 1755005639
transform 1 0 37433 0 1 20645
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_102
timestamp 1755005639
transform 1 0 39545 0 1 18533
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_103
timestamp 1755005639
transform 1 0 35057 0 1 23021
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_104
timestamp 1755005639
transform 1 0 39149 0 1 18929
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_105
timestamp 1755005639
transform 1 0 33341 0 1 24737
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_106
timestamp 1755005639
transform 1 0 33473 0 1 24605
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_107
timestamp 1755005639
transform 1 0 18689 0 1 39389
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_108
timestamp 1755005639
transform 1 0 23969 0 1 34109
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_109
timestamp 1755005639
transform 1 0 23045 0 1 35033
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_110
timestamp 1755005639
transform 1 0 23309 0 1 34769
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_111
timestamp 1755005639
transform 1 0 23441 0 1 34637
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_112
timestamp 1755005639
transform 1 0 23573 0 1 34505
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_113
timestamp 1755005639
transform 1 0 23705 0 1 34373
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_114
timestamp 1755005639
transform 1 0 23837 0 1 34241
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_115
timestamp 1755005639
transform 1 0 24101 0 1 33977
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_116
timestamp 1755005639
transform 1 0 24233 0 1 33845
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_117
timestamp 1755005639
transform 1 0 24365 0 1 33713
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_118
timestamp 1755005639
transform 1 0 24497 0 1 33581
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_119
timestamp 1755005639
transform 1 0 24629 0 1 33449
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_120
timestamp 1755005639
transform 1 0 24761 0 1 33317
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_121
timestamp 1755005639
transform 1 0 25025 0 1 33053
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_122
timestamp 1755005639
transform 1 0 23177 0 1 34901
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_123
timestamp 1755005639
transform 1 0 22913 0 1 35165
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_124
timestamp 1755005639
transform 1 0 22781 0 1 35297
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_125
timestamp 1755005639
transform 1 0 22649 0 1 35429
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_126
timestamp 1755005639
transform 1 0 22517 0 1 35561
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_127
timestamp 1755005639
transform 1 0 22385 0 1 35693
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_128
timestamp 1755005639
transform 1 0 22253 0 1 35825
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_129
timestamp 1755005639
transform 1 0 22121 0 1 35957
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_130
timestamp 1755005639
transform 1 0 21989 0 1 36089
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_131
timestamp 1755005639
transform 1 0 21857 0 1 36221
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_132
timestamp 1755005639
transform 1 0 21725 0 1 36353
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_133
timestamp 1755005639
transform 1 0 21593 0 1 36485
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_134
timestamp 1755005639
transform 1 0 21461 0 1 36617
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_135
timestamp 1755005639
transform 1 0 21329 0 1 36749
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_136
timestamp 1755005639
transform 1 0 21065 0 1 37013
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_137
timestamp 1755005639
transform 1 0 24893 0 1 33185
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_138
timestamp 1755005639
transform 1 0 18557 0 1 39521
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_139
timestamp 1755005639
transform 1 0 18425 0 1 39653
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_140
timestamp 1755005639
transform 1 0 18293 0 1 39785
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_141
timestamp 1755005639
transform 1 0 18161 0 1 39917
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_142
timestamp 1755005639
transform 1 0 16973 0 1 41105
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_143
timestamp 1755005639
transform 1 0 18029 0 1 40049
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_144
timestamp 1755005639
transform 1 0 17897 0 1 40181
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_145
timestamp 1755005639
transform 1 0 17765 0 1 40313
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_146
timestamp 1755005639
transform 1 0 17633 0 1 40445
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_147
timestamp 1755005639
transform 1 0 17501 0 1 40577
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_148
timestamp 1755005639
transform 1 0 17369 0 1 40709
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_149
timestamp 1755005639
transform 1 0 27401 0 1 30677
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_150
timestamp 1755005639
transform 1 0 27269 0 1 30809
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_151
timestamp 1755005639
transform 1 0 27137 0 1 30941
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_152
timestamp 1755005639
transform 1 0 21197 0 1 36881
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_153
timestamp 1755005639
transform 1 0 26873 0 1 31205
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_154
timestamp 1755005639
transform 1 0 26741 0 1 31337
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_155
timestamp 1755005639
transform 1 0 26609 0 1 31469
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_156
timestamp 1755005639
transform 1 0 26477 0 1 31601
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_157
timestamp 1755005639
transform 1 0 26345 0 1 31733
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_158
timestamp 1755005639
transform 1 0 26213 0 1 31865
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_159
timestamp 1755005639
transform 1 0 26081 0 1 31997
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_160
timestamp 1755005639
transform 1 0 25949 0 1 32129
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_161
timestamp 1755005639
transform 1 0 25817 0 1 32261
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_162
timestamp 1755005639
transform 1 0 25685 0 1 32393
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_163
timestamp 1755005639
transform 1 0 25553 0 1 32525
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_164
timestamp 1755005639
transform 1 0 25421 0 1 32657
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_165
timestamp 1755005639
transform 1 0 25289 0 1 32789
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_166
timestamp 1755005639
transform 1 0 25157 0 1 32921
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_167
timestamp 1755005639
transform 1 0 27005 0 1 31073
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_168
timestamp 1755005639
transform 1 0 17105 0 1 40973
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_169
timestamp 1755005639
transform 1 0 16841 0 1 41237
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_170
timestamp 1755005639
transform 1 0 16709 0 1 41369
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_171
timestamp 1755005639
transform 1 0 16577 0 1 41501
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_172
timestamp 1755005639
transform 1 0 16445 0 1 41633
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_173
timestamp 1755005639
transform 1 0 16313 0 1 41765
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_174
timestamp 1755005639
transform 1 0 16181 0 1 41897
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_175
timestamp 1755005639
transform 1 0 19085 0 1 38993
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_176
timestamp 1755005639
transform 1 0 20933 0 1 37145
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_177
timestamp 1755005639
transform 1 0 20801 0 1 37277
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_178
timestamp 1755005639
transform 1 0 20669 0 1 37409
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_179
timestamp 1755005639
transform 1 0 20537 0 1 37541
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_180
timestamp 1755005639
transform 1 0 20405 0 1 37673
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_181
timestamp 1755005639
transform 1 0 20273 0 1 37805
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_182
timestamp 1755005639
transform 1 0 20141 0 1 37937
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_183
timestamp 1755005639
transform 1 0 20009 0 1 38069
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_184
timestamp 1755005639
transform 1 0 19877 0 1 38201
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_185
timestamp 1755005639
transform 1 0 19745 0 1 38333
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_186
timestamp 1755005639
transform 1 0 19613 0 1 38465
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_187
timestamp 1755005639
transform 1 0 19481 0 1 38597
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_188
timestamp 1755005639
transform 1 0 19349 0 1 38729
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_189
timestamp 1755005639
transform 1 0 19217 0 1 38861
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_190
timestamp 1755005639
transform 1 0 17237 0 1 40841
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_191
timestamp 1755005639
transform 1 0 18953 0 1 39125
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_192
timestamp 1755005639
transform 1 0 18821 0 1 39257
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_193
timestamp 1755005639
transform 1 0 29117 0 1 28961
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_194
timestamp 1755005639
transform 1 0 28985 0 1 29093
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_195
timestamp 1755005639
transform 1 0 28721 0 1 29357
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_196
timestamp 1755005639
transform 1 0 28589 0 1 29489
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_197
timestamp 1755005639
transform 1 0 28457 0 1 29621
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_198
timestamp 1755005639
transform 1 0 28325 0 1 29753
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_199
timestamp 1755005639
transform 1 0 28193 0 1 29885
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_200
timestamp 1755005639
transform 1 0 28061 0 1 30017
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_201
timestamp 1755005639
transform 1 0 27929 0 1 30149
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_202
timestamp 1755005639
transform 1 0 27797 0 1 30281
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_203
timestamp 1755005639
transform 1 0 27665 0 1 30413
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_204
timestamp 1755005639
transform 1 0 29249 0 1 28829
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_205
timestamp 1755005639
transform 1 0 28853 0 1 29225
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_206
timestamp 1755005639
transform 1 0 29513 0 1 28565
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_207
timestamp 1755005639
transform 1 0 30437 0 1 27641
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_208
timestamp 1755005639
transform 1 0 30305 0 1 27773
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_209
timestamp 1755005639
transform 1 0 30173 0 1 27905
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_210
timestamp 1755005639
transform 1 0 30041 0 1 28037
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_211
timestamp 1755005639
transform 1 0 29909 0 1 28169
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_212
timestamp 1755005639
transform 1 0 29777 0 1 28301
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_213
timestamp 1755005639
transform 1 0 29645 0 1 28433
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_214
timestamp 1755005639
transform 1 0 29381 0 1 28697
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_215
timestamp 1755005639
transform 1 0 27533 0 1 30545
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_216
timestamp 1755005639
transform 1 0 30569 0 1 27509
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_217
timestamp 1755005639
transform 1 0 13937 0 1 44141
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_218
timestamp 1755005639
transform 1 0 13805 0 1 44273
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_219
timestamp 1755005639
transform 1 0 13673 0 1 44405
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_220
timestamp 1755005639
transform 1 0 13541 0 1 44537
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_221
timestamp 1755005639
transform 1 0 13409 0 1 44669
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_222
timestamp 1755005639
transform 1 0 13277 0 1 44801
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_223
timestamp 1755005639
transform 1 0 15125 0 1 42953
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_224
timestamp 1755005639
transform 1 0 15917 0 1 42161
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_225
timestamp 1755005639
transform 1 0 15785 0 1 42293
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_226
timestamp 1755005639
transform 1 0 15653 0 1 42425
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_227
timestamp 1755005639
transform 1 0 15521 0 1 42557
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_228
timestamp 1755005639
transform 1 0 15389 0 1 42689
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_229
timestamp 1755005639
transform 1 0 15257 0 1 42821
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_230
timestamp 1755005639
transform 1 0 14993 0 1 43085
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_231
timestamp 1755005639
transform 1 0 14861 0 1 43217
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_232
timestamp 1755005639
transform 1 0 14729 0 1 43349
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_233
timestamp 1755005639
transform 1 0 14597 0 1 43481
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_234
timestamp 1755005639
transform 1 0 14465 0 1 43613
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_235
timestamp 1755005639
transform 1 0 14333 0 1 43745
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_236
timestamp 1755005639
transform 1 0 14201 0 1 43877
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_237
timestamp 1755005639
transform 1 0 14069 0 1 44009
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_238
timestamp 1755005639
transform 1 0 16049 0 1 42029
box 0 0 1 1
use M1_PSUB_CDNS_40661953145674  M1_PSUB_CDNS_40661953145674_239
timestamp 1755005639
transform 1 0 42053 0 1 16025
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_0
timestamp 1755005639
transform 1 0 70641 0 1 24306
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_1
timestamp 1755005639
transform 1 0 70641 0 1 67516
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_2
timestamp 1755005639
transform 1 0 70641 0 1 59520
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_3
timestamp 1755005639
transform 1 0 70641 0 1 54702
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_4
timestamp 1755005639
transform 1 0 70641 0 1 53122
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_5
timestamp 1755005639
transform 1 0 70641 0 1 56310
box 0 0 1 1
use M3_M2_CDNS_40661953145675  M3_M2_CDNS_40661953145675_6
timestamp 1755005639
transform 1 0 70641 0 1 41897
box 0 0 1 1
use M3_M2_CDNS_40661953145676  M3_M2_CDNS_40661953145676_0
timestamp 1755005639
transform 1 0 70641 0 1 28320
box 0 0 1 1
use M3_M2_CDNS_40661953145676  M3_M2_CDNS_40661953145676_1
timestamp 1755005639
transform 1 0 70641 0 1 31488
box 0 0 1 1
use M3_M2_CDNS_40661953145676  M3_M2_CDNS_40661953145676_2
timestamp 1755005639
transform 1 0 70641 0 1 34700
box 0 0 1 1
use M3_M2_CDNS_40661953145676  M3_M2_CDNS_40661953145676_3
timestamp 1755005639
transform 1 0 70641 0 1 37900
box 0 0 1 1
use M3_M2_CDNS_40661953145676  M3_M2_CDNS_40661953145676_4
timestamp 1755005639
transform 1 0 70641 0 1 44307
box 0 0 1 1
<< labels >>
rlabel metal3 s 70454 64211 70454 64211 4 VSS
port 1 nsew
rlabel metal3 s 70454 62776 70454 62776 4 VDD
port 2 nsew
rlabel metal3 s 70454 61011 70454 61011 4 DVSS
port 3 nsew
rlabel metal3 s 70454 65976 70454 65976 4 DVSS
port 3 nsew
rlabel metal3 s 70454 69002 70454 69002 4 DVSS
port 3 nsew
rlabel metal3 s 70454 67411 70454 67411 4 DVDD
port 4 nsew
rlabel metal3 s 70454 59576 70454 59576 4 DVDD
port 4 nsew
rlabel metal3 s 70454 57811 70454 57811 4 DVSS
port 3 nsew
rlabel metal3 s 70454 56376 70454 56376 4 DVDD
port 4 nsew
rlabel metal3 s 70454 54611 70454 54611 4 DVDD
port 4 nsew
rlabel metal3 s 70454 53176 70454 53176 4 DVDD
port 4 nsew
rlabel metal3 s 70559 51411 70559 51411 4 VDD
port 2 nsew
rlabel metal3 s 70559 49976 70559 49976 4 VSS
port 1 nsew
rlabel metal3 s 70454 47548 70454 47548 4 DVSS
port 3 nsew
rlabel metal3 s 70454 44321 70454 44321 4 DVDD
port 4 nsew
rlabel metal3 s 70454 40295 70454 40295 4 DVSS
port 3 nsew
rlabel metal3 s 70454 41930 70454 41930 4 DVDD
port 4 nsew
rlabel metal3 s 70454 37912 70454 37912 4 DVDD
port 4 nsew
rlabel metal3 s 70454 34676 70454 34676 4 DVDD
port 4 nsew
rlabel metal3 s 70454 31562 70454 31562 4 DVDD
port 4 nsew
rlabel metal3 s 70454 28347 70454 28347 4 DVDD
port 4 nsew
rlabel metal3 s 70454 26053 70454 26053 4 DVSS
port 3 nsew
rlabel metal3 s 70454 24237 70454 24237 4 DVDD
port 4 nsew
rlabel metal3 s 70454 21860 70454 21860 4 DVSS
port 3 nsew
rlabel metal3 s 70385 18874 70385 18874 4 DVSS
port 3 nsew
rlabel metal3 s 70432 15703 70432 15703 4 DVSS
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 71000 71000
string GDS_END 17209510
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17191198
string path 329.850 1126.950 329.850 1122.100 1122.100 329.850 1155.475 329.850 
<< end >>
