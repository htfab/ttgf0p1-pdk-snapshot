magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< metal1 >>
rect 3 4188 203 4200
rect 3 4136 15 4188
rect 67 4136 139 4188
rect 191 4136 203 4188
rect 3 4064 203 4136
rect 3 4012 15 4064
rect 67 4012 139 4064
rect 191 4012 203 4064
rect 3 3940 203 4012
rect 3 3888 15 3940
rect 67 3888 139 3940
rect 191 3888 203 3940
rect 3 3816 203 3888
rect 3 3764 15 3816
rect 67 3764 139 3816
rect 191 3764 203 3816
rect 3 3692 203 3764
rect 3 3640 15 3692
rect 67 3640 139 3692
rect 191 3640 203 3692
rect 3 3568 203 3640
rect 3 3516 15 3568
rect 67 3516 139 3568
rect 191 3516 203 3568
rect 3 3444 203 3516
rect 3 3392 15 3444
rect 67 3392 139 3444
rect 191 3392 203 3444
rect 3 3320 203 3392
rect 3 3268 15 3320
rect 67 3268 139 3320
rect 191 3268 203 3320
rect 3 3256 203 3268
rect 1020 4188 1220 4200
rect 1020 4136 1032 4188
rect 1084 4136 1156 4188
rect 1208 4136 1220 4188
rect 1020 4064 1220 4136
rect 1020 4012 1032 4064
rect 1084 4012 1156 4064
rect 1208 4012 1220 4064
rect 1020 3940 1220 4012
rect 1020 3888 1032 3940
rect 1084 3888 1156 3940
rect 1208 3888 1220 3940
rect 1020 3816 1220 3888
rect 1020 3764 1032 3816
rect 1084 3764 1156 3816
rect 1208 3764 1220 3816
rect 1020 3692 1220 3764
rect 1020 3640 1032 3692
rect 1084 3640 1156 3692
rect 1208 3640 1220 3692
rect 1020 3568 1220 3640
rect 1020 3516 1032 3568
rect 1084 3516 1156 3568
rect 1208 3516 1220 3568
rect 1020 3444 1220 3516
rect 1020 3392 1032 3444
rect 1084 3392 1156 3444
rect 1208 3392 1220 3444
rect 1020 3320 1220 3392
rect 1020 3268 1032 3320
rect 1084 3268 1156 3320
rect 1208 3268 1220 3320
rect 1020 3256 1220 3268
<< via1 >>
rect 15 4136 67 4188
rect 139 4136 191 4188
rect 15 4012 67 4064
rect 139 4012 191 4064
rect 15 3888 67 3940
rect 139 3888 191 3940
rect 15 3764 67 3816
rect 139 3764 191 3816
rect 15 3640 67 3692
rect 139 3640 191 3692
rect 15 3516 67 3568
rect 139 3516 191 3568
rect 15 3392 67 3444
rect 139 3392 191 3444
rect 15 3268 67 3320
rect 139 3268 191 3320
rect 1032 4136 1084 4188
rect 1156 4136 1208 4188
rect 1032 4012 1084 4064
rect 1156 4012 1208 4064
rect 1032 3888 1084 3940
rect 1156 3888 1208 3940
rect 1032 3764 1084 3816
rect 1156 3764 1208 3816
rect 1032 3640 1084 3692
rect 1156 3640 1208 3692
rect 1032 3516 1084 3568
rect 1156 3516 1208 3568
rect 1032 3392 1084 3444
rect 1156 3392 1208 3444
rect 1032 3268 1084 3320
rect 1156 3268 1208 3320
<< metal2 >>
rect 495 6371 719 7462
rect 495 6315 516 6371
rect 572 6315 640 6371
rect 696 6315 719 6371
rect 495 6247 719 6315
rect 495 6191 516 6247
rect 572 6191 640 6247
rect 696 6191 719 6247
rect 495 6123 719 6191
rect 495 6067 516 6123
rect 572 6067 640 6123
rect 696 6067 719 6123
rect -8 5681 216 5708
rect -8 5625 16 5681
rect 72 5625 140 5681
rect 196 5625 216 5681
rect -8 5557 216 5625
rect -8 5501 16 5557
rect 72 5501 140 5557
rect 196 5501 216 5557
rect -8 5433 216 5501
rect -8 5377 16 5433
rect 72 5377 140 5433
rect 196 5377 216 5433
rect -8 4667 216 5377
rect -8 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 216 4667
rect -8 4543 216 4611
rect -8 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 216 4543
rect -8 4419 216 4487
rect -8 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 216 4419
rect -8 4188 216 4363
rect -8 4136 15 4188
rect 67 4136 139 4188
rect 191 4136 216 4188
rect -8 4064 216 4136
rect -8 4012 15 4064
rect 67 4012 139 4064
rect 191 4012 216 4064
rect -8 3940 216 4012
rect -8 3888 15 3940
rect 67 3888 139 3940
rect 191 3888 216 3940
rect -8 3816 216 3888
rect -8 3764 15 3816
rect 67 3764 139 3816
rect 191 3764 216 3816
rect -8 3692 216 3764
rect -8 3640 15 3692
rect 67 3640 139 3692
rect 191 3640 216 3692
rect -8 3568 216 3640
rect -8 3516 15 3568
rect 67 3516 139 3568
rect 191 3516 216 3568
rect -8 3444 216 3516
rect -8 3392 15 3444
rect 67 3392 139 3444
rect 191 3392 216 3444
rect -8 3320 216 3392
rect -8 3268 15 3320
rect 67 3268 139 3320
rect 191 3268 216 3320
rect 495 4034 719 6067
rect 495 3978 516 4034
rect 572 3978 640 4034
rect 696 3978 719 4034
rect 495 3910 719 3978
rect 495 3854 516 3910
rect 572 3854 640 3910
rect 696 3854 719 3910
rect 495 3786 719 3854
rect 495 3730 516 3786
rect 572 3730 640 3786
rect 696 3730 719 3786
rect 495 3662 719 3730
rect 495 3606 516 3662
rect 572 3606 640 3662
rect 696 3606 719 3662
rect 495 3538 719 3606
rect 495 3482 516 3538
rect 572 3482 640 3538
rect 696 3482 719 3538
rect 495 3414 719 3482
rect 495 3358 516 3414
rect 572 3358 640 3414
rect 696 3358 719 3414
rect 495 3313 719 3358
rect 1011 5681 1235 5708
rect 1011 5625 1033 5681
rect 1089 5625 1157 5681
rect 1213 5625 1235 5681
rect 1011 5557 1235 5625
rect 1011 5501 1033 5557
rect 1089 5501 1157 5557
rect 1213 5501 1235 5557
rect 1011 5433 1235 5501
rect 1011 5377 1033 5433
rect 1089 5377 1157 5433
rect 1213 5377 1235 5433
rect 1011 4667 1235 5377
rect 1011 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1235 4667
rect 1011 4543 1235 4611
rect 1011 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1235 4543
rect 1011 4419 1235 4487
rect 1011 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1235 4419
rect 1011 4188 1235 4363
rect 1011 4136 1032 4188
rect 1084 4136 1156 4188
rect 1208 4136 1235 4188
rect 1011 4064 1235 4136
rect 1011 4012 1032 4064
rect 1084 4012 1156 4064
rect 1208 4012 1235 4064
rect 1011 3940 1235 4012
rect 1011 3888 1032 3940
rect 1084 3888 1156 3940
rect 1208 3888 1235 3940
rect 1011 3816 1235 3888
rect 1011 3764 1032 3816
rect 1084 3764 1156 3816
rect 1208 3764 1235 3816
rect 1011 3692 1235 3764
rect 1011 3640 1032 3692
rect 1084 3640 1156 3692
rect 1208 3640 1235 3692
rect 1011 3568 1235 3640
rect 1011 3516 1032 3568
rect 1084 3516 1156 3568
rect 1208 3516 1235 3568
rect 1011 3444 1235 3516
rect 1011 3392 1032 3444
rect 1084 3392 1156 3444
rect 1208 3392 1235 3444
rect 1011 3320 1235 3392
rect -8 3065 216 3268
rect 1011 3268 1032 3320
rect 1084 3268 1156 3320
rect 1208 3268 1235 3320
rect 1011 3065 1235 3268
<< via2 >>
rect 516 6315 572 6371
rect 640 6315 696 6371
rect 516 6191 572 6247
rect 640 6191 696 6247
rect 516 6067 572 6123
rect 640 6067 696 6123
rect 16 5625 72 5681
rect 140 5625 196 5681
rect 16 5501 72 5557
rect 140 5501 196 5557
rect 16 5377 72 5433
rect 140 5377 196 5433
rect 16 4611 72 4667
rect 140 4611 196 4667
rect 16 4487 72 4543
rect 140 4487 196 4543
rect 16 4363 72 4419
rect 140 4363 196 4419
rect 516 3978 572 4034
rect 640 3978 696 4034
rect 516 3854 572 3910
rect 640 3854 696 3910
rect 516 3730 572 3786
rect 640 3730 696 3786
rect 516 3606 572 3662
rect 640 3606 696 3662
rect 516 3482 572 3538
rect 640 3482 696 3538
rect 516 3358 572 3414
rect 640 3358 696 3414
rect 1033 5625 1089 5681
rect 1157 5625 1213 5681
rect 1033 5501 1089 5557
rect 1157 5501 1213 5557
rect 1033 5377 1089 5433
rect 1157 5377 1213 5433
rect 1033 4611 1089 4667
rect 1157 4611 1213 4667
rect 1033 4487 1089 4543
rect 1157 4487 1213 4543
rect 1033 4363 1089 4419
rect 1157 4363 1213 4419
<< metal3 >>
rect 506 6371 706 6381
rect 506 6315 516 6371
rect 572 6315 640 6371
rect 696 6315 706 6371
rect 506 6247 706 6315
rect 506 6191 516 6247
rect 572 6191 640 6247
rect 696 6191 706 6247
rect 506 6123 706 6191
rect 506 6067 516 6123
rect 572 6067 640 6123
rect 696 6067 706 6123
rect 506 6057 706 6067
rect 6 5681 206 5691
rect 6 5625 16 5681
rect 72 5625 140 5681
rect 196 5625 206 5681
rect 6 5557 206 5625
rect 6 5501 16 5557
rect 72 5501 140 5557
rect 196 5501 206 5557
rect 6 5433 206 5501
rect 6 5377 16 5433
rect 72 5377 140 5433
rect 196 5377 206 5433
rect 6 5367 206 5377
rect 1023 5681 1223 5691
rect 1023 5625 1033 5681
rect 1089 5625 1157 5681
rect 1213 5625 1223 5681
rect 1023 5557 1223 5625
rect 1023 5501 1033 5557
rect 1089 5501 1157 5557
rect 1213 5501 1223 5557
rect 1023 5433 1223 5501
rect 1023 5377 1033 5433
rect 1089 5377 1157 5433
rect 1213 5377 1223 5433
rect 1023 5367 1223 5377
rect 6 4667 206 4677
rect 6 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 206 4667
rect 6 4543 206 4611
rect 6 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 206 4543
rect 6 4419 206 4487
rect 6 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 206 4419
rect 6 4353 206 4363
rect 1023 4667 1223 4677
rect 1023 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1223 4667
rect 1023 4543 1223 4611
rect 1023 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1223 4543
rect 1023 4419 1223 4487
rect 1023 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1223 4419
rect 1023 4353 1223 4363
rect 506 4034 706 4044
rect 506 3978 516 4034
rect 572 3978 640 4034
rect 696 3978 706 4034
rect 506 3910 706 3978
rect 506 3854 516 3910
rect 572 3854 640 3910
rect 696 3854 706 3910
rect 506 3786 706 3854
rect 506 3730 516 3786
rect 572 3730 640 3786
rect 696 3730 706 3786
rect 506 3662 706 3730
rect 506 3606 516 3662
rect 572 3606 640 3662
rect 696 3606 706 3662
rect 506 3538 706 3606
rect 506 3482 516 3538
rect 572 3482 640 3538
rect 696 3482 706 3538
rect 506 3414 706 3482
rect 506 3358 516 3414
rect 572 3358 640 3414
rect 696 3358 706 3414
rect 506 3348 706 3358
use M2_M14310591302097_512x8m81  M2_M14310591302097_512x8m81_0
timestamp 1755005639
transform 1 0 1120 0 1 3728
box 0 0 1 1
use M2_M14310591302097_512x8m81  M2_M14310591302097_512x8m81_1
timestamp 1755005639
transform 1 0 103 0 1 3728
box 0 0 1 1
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_0
timestamp 1755005639
transform 1 0 606 0 1 6219
box 0 0 1 1
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_1
timestamp 1755005639
transform 1 0 1123 0 1 4515
box 0 0 1 1
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_2
timestamp 1755005639
transform 1 0 1123 0 1 5529
box 0 0 1 1
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_3
timestamp 1755005639
transform 1 0 106 0 1 5529
box 0 0 1 1
use M3_M24310591302095_512x8m81  M3_M24310591302095_512x8m81_4
timestamp 1755005639
transform 1 0 106 0 1 4515
box 0 0 1 1
use M3_M243105913020102_512x8m81  M3_M243105913020102_512x8m81_0
timestamp 1755005639
transform 1 0 606 0 1 3696
box 0 0 1 1
<< properties >>
string GDS_END 1128834
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 1128222
<< end >>
