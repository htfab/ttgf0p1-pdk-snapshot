magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 3670 1094
<< pwell >>
rect -86 -86 3670 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 716 175 836 315
rect 940 175 1060 315
rect 1164 175 1284 315
rect 1332 175 1452 315
rect 1500 175 1620 315
rect 1764 175 1884 315
rect 2003 175 2123 315
rect 2231 175 2351 315
rect 2455 175 2575 315
rect 2679 175 2799 315
rect 2939 175 3059 333
rect 3307 69 3427 333
<< mvpmos >>
rect 132 573 232 849
rect 336 573 436 849
rect 684 573 784 773
rect 888 573 988 773
rect 1092 573 1192 773
rect 1296 573 1396 773
rect 1500 573 1600 773
rect 1848 635 1948 835
rect 2052 635 2152 835
rect 2256 635 2356 835
rect 2475 635 2575 835
rect 2723 635 2823 911
rect 2927 635 3027 911
rect 3307 573 3407 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 468 274 497 320
rect 543 274 556 320
rect 2859 315 2939 333
rect 468 175 556 274
rect 628 234 716 315
rect 628 188 641 234
rect 687 188 716 234
rect 628 175 716 188
rect 836 302 940 315
rect 836 256 865 302
rect 911 256 940 302
rect 836 175 940 256
rect 1060 302 1164 315
rect 1060 256 1089 302
rect 1135 256 1164 302
rect 1060 175 1164 256
rect 1284 175 1332 315
rect 1452 175 1500 315
rect 1620 234 1764 315
rect 1620 188 1649 234
rect 1695 188 1764 234
rect 1620 175 1764 188
rect 1884 302 2003 315
rect 1884 256 1927 302
rect 1973 256 2003 302
rect 1884 175 2003 256
rect 2123 302 2231 315
rect 2123 256 2156 302
rect 2202 256 2231 302
rect 2123 175 2231 256
rect 2351 302 2455 315
rect 2351 256 2380 302
rect 2426 256 2455 302
rect 2351 175 2455 256
rect 2575 234 2679 315
rect 2575 188 2604 234
rect 2650 188 2679 234
rect 2575 175 2679 188
rect 2799 175 2939 315
rect 3059 320 3147 333
rect 3059 274 3088 320
rect 3134 274 3147 320
rect 3059 175 3147 274
rect 3219 320 3307 333
rect 3219 180 3232 320
rect 3278 180 3307 320
rect 3219 69 3307 180
rect 3427 222 3515 333
rect 3427 82 3456 222
rect 3502 82 3515 222
rect 3427 69 3515 82
<< mvpdiff >>
rect 44 739 132 849
rect 44 599 57 739
rect 103 599 132 739
rect 44 573 132 599
rect 232 836 336 849
rect 232 696 261 836
rect 307 696 336 836
rect 232 573 336 696
rect 436 726 524 849
rect 2635 898 2723 911
rect 2635 852 2648 898
rect 2694 852 2723 898
rect 2635 835 2723 852
rect 1760 822 1848 835
rect 436 586 465 726
rect 511 586 524 726
rect 436 573 524 586
rect 596 760 684 773
rect 596 714 609 760
rect 655 714 684 760
rect 596 573 684 714
rect 784 726 888 773
rect 784 586 813 726
rect 859 586 888 726
rect 784 573 888 586
rect 988 726 1092 773
rect 988 586 1017 726
rect 1063 586 1092 726
rect 988 573 1092 586
rect 1192 760 1296 773
rect 1192 620 1221 760
rect 1267 620 1296 760
rect 1192 573 1296 620
rect 1396 760 1500 773
rect 1396 714 1425 760
rect 1471 714 1500 760
rect 1396 573 1500 714
rect 1600 760 1688 773
rect 1600 620 1629 760
rect 1675 620 1688 760
rect 1760 682 1773 822
rect 1819 682 1848 822
rect 1760 635 1848 682
rect 1948 788 2052 835
rect 1948 648 1977 788
rect 2023 648 2052 788
rect 1948 635 2052 648
rect 2152 788 2256 835
rect 2152 648 2181 788
rect 2227 648 2256 788
rect 2152 635 2256 648
rect 2356 694 2475 835
rect 2356 648 2385 694
rect 2431 648 2475 694
rect 2356 635 2475 648
rect 2575 635 2723 835
rect 2823 694 2927 911
rect 2823 648 2852 694
rect 2898 648 2927 694
rect 2823 635 2927 648
rect 3027 898 3115 911
rect 3027 758 3056 898
rect 3102 758 3115 898
rect 3027 635 3115 758
rect 3219 726 3307 939
rect 1600 573 1688 620
rect 3219 586 3232 726
rect 3278 586 3307 726
rect 3219 573 3307 586
rect 3407 926 3495 939
rect 3407 786 3436 926
rect 3482 786 3495 926
rect 3407 573 3495 786
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 641 188 687 234
rect 865 256 911 302
rect 1089 256 1135 302
rect 1649 188 1695 234
rect 1927 256 1973 302
rect 2156 256 2202 302
rect 2380 256 2426 302
rect 2604 188 2650 234
rect 3088 274 3134 320
rect 3232 180 3278 320
rect 3456 82 3502 222
<< mvpdiffc >>
rect 57 599 103 739
rect 261 696 307 836
rect 2648 852 2694 898
rect 465 586 511 726
rect 609 714 655 760
rect 813 586 859 726
rect 1017 586 1063 726
rect 1221 620 1267 760
rect 1425 714 1471 760
rect 1629 620 1675 760
rect 1773 682 1819 822
rect 1977 648 2023 788
rect 2181 648 2227 788
rect 2385 648 2431 694
rect 2852 648 2898 694
rect 3056 758 3102 898
rect 3232 586 3278 726
rect 3436 786 3482 926
<< polysilicon >>
rect 336 909 988 949
rect 132 849 232 893
rect 336 849 436 909
rect 684 773 784 817
rect 888 773 988 909
rect 1092 927 2152 967
rect 1092 852 1192 927
rect 1092 806 1105 852
rect 1151 806 1192 852
rect 1848 835 1948 879
rect 2052 835 2152 927
rect 2723 911 2823 955
rect 2927 911 3027 955
rect 3307 939 3407 983
rect 2256 835 2356 879
rect 2475 835 2575 879
rect 1092 773 1192 806
rect 1296 773 1396 817
rect 1500 773 1600 817
rect 132 504 232 573
rect 132 458 145 504
rect 191 458 232 504
rect 132 377 232 458
rect 336 412 436 573
rect 336 393 361 412
rect 124 333 244 377
rect 348 366 361 393
rect 407 393 436 412
rect 684 508 784 573
rect 888 529 988 573
rect 1092 529 1192 573
rect 684 462 697 508
rect 743 462 784 508
rect 407 366 468 393
rect 684 375 784 462
rect 1092 435 1132 529
rect 1296 513 1396 573
rect 940 395 1132 435
rect 1332 436 1404 513
rect 348 333 468 366
rect 716 315 836 375
rect 940 315 1060 395
rect 1212 394 1284 407
rect 1212 359 1225 394
rect 1164 348 1225 359
rect 1271 348 1284 394
rect 1164 315 1284 348
rect 1332 390 1345 436
rect 1391 390 1404 436
rect 1332 359 1404 390
rect 1500 359 1600 573
rect 1848 563 1948 635
rect 1848 522 1861 563
rect 1844 517 1861 522
rect 1907 517 1948 563
rect 1844 504 1948 517
rect 1844 359 1884 504
rect 2052 495 2152 635
rect 2256 602 2356 635
rect 2256 556 2269 602
rect 2315 556 2356 602
rect 2256 543 2356 556
rect 2475 602 2575 635
rect 2475 556 2516 602
rect 2562 556 2575 602
rect 2052 455 2351 495
rect 1332 315 1452 359
rect 1500 315 1620 359
rect 1764 315 1884 359
rect 2003 394 2123 407
rect 2003 348 2064 394
rect 2110 348 2123 394
rect 2003 315 2123 348
rect 2231 315 2351 455
rect 2475 359 2575 556
rect 2723 394 2823 635
rect 2723 381 2736 394
rect 2455 315 2575 359
rect 2679 348 2736 381
rect 2782 381 2823 394
rect 2927 602 3027 635
rect 2927 556 2944 602
rect 2990 556 3027 602
rect 2927 393 3027 556
rect 3307 465 3407 573
rect 3127 452 3407 465
rect 3127 406 3140 452
rect 3186 406 3407 452
rect 3127 393 3407 406
rect 2782 348 2799 381
rect 2679 315 2799 348
rect 2939 333 3059 393
rect 3307 377 3407 393
rect 3307 333 3427 377
rect 124 131 244 175
rect 348 83 468 175
rect 716 131 836 175
rect 940 131 1060 175
rect 1164 83 1284 175
rect 1332 131 1452 175
rect 348 43 1284 83
rect 1500 83 1620 175
rect 1764 131 1884 175
rect 2003 131 2123 175
rect 2231 131 2351 175
rect 2455 131 2575 175
rect 2679 131 2799 175
rect 2939 131 3059 175
rect 2723 83 2799 131
rect 1500 43 2823 83
rect 3307 25 3427 69
<< polycontact >>
rect 1105 806 1151 852
rect 145 458 191 504
rect 361 366 407 412
rect 697 462 743 508
rect 1225 348 1271 394
rect 1345 390 1391 436
rect 1861 517 1907 563
rect 2269 556 2315 602
rect 2516 556 2562 602
rect 2064 348 2110 394
rect 2736 348 2782 394
rect 2944 556 2990 602
rect 3140 406 3186 452
<< metal1 >>
rect 0 926 3584 1098
rect 0 918 3436 926
rect 261 836 307 918
rect 57 739 103 750
rect 609 760 655 918
rect 261 685 307 696
rect 465 726 511 737
rect 103 599 407 634
rect 57 588 407 599
rect 133 504 315 542
rect 133 458 145 504
rect 191 458 315 504
rect 133 447 315 458
rect 361 412 407 588
rect 361 348 407 366
rect 49 320 407 348
rect 95 302 407 320
rect 609 703 655 714
rect 701 852 1151 863
rect 701 806 1105 852
rect 701 795 1151 806
rect 701 657 747 795
rect 1221 760 1267 771
rect 511 611 747 657
rect 813 726 859 737
rect 511 586 543 611
rect 465 320 543 586
rect 589 508 754 542
rect 589 462 697 508
rect 743 462 754 508
rect 49 263 95 274
rect 465 274 497 320
rect 465 263 543 274
rect 813 302 859 586
rect 1017 726 1063 737
rect 1425 760 1471 918
rect 1773 822 1819 918
rect 2637 898 2705 918
rect 2637 852 2648 898
rect 2694 852 2705 898
rect 3056 898 3102 918
rect 1425 703 1471 714
rect 1629 760 1675 771
rect 1267 620 1629 655
rect 1773 671 1819 682
rect 1977 788 2023 799
rect 1221 609 1675 620
rect 1063 586 1134 599
rect 1017 563 1134 586
rect 1017 553 1861 563
rect 1089 517 1861 553
rect 1907 517 1918 563
rect 1089 302 1135 517
rect 1977 472 2023 648
rect 1928 436 2023 472
rect 813 256 865 302
rect 911 256 922 302
rect 1225 394 1271 405
rect 1334 390 1345 436
rect 1391 426 2023 436
rect 2156 788 2990 799
rect 2156 648 2181 788
rect 2227 753 2990 788
rect 2156 637 2227 648
rect 2380 694 2431 705
rect 2380 648 2385 694
rect 1391 390 1973 426
rect 1225 337 1271 348
rect 1225 291 1881 337
rect 1089 245 1135 256
rect 273 234 319 245
rect 273 90 319 188
rect 641 234 687 245
rect 641 90 687 188
rect 1649 234 1695 245
rect 1649 90 1695 188
rect 1835 199 1881 291
rect 1927 302 1973 390
rect 1927 245 1973 256
rect 2064 394 2110 405
rect 2064 199 2110 348
rect 2156 302 2202 637
rect 2156 245 2202 256
rect 2269 602 2315 613
rect 2269 199 2315 556
rect 2380 302 2431 648
rect 2516 694 2898 705
rect 2516 659 2852 694
rect 2516 602 2562 659
rect 2516 545 2562 556
rect 2852 499 2898 648
rect 2944 602 2990 753
rect 3482 918 3584 926
rect 3436 775 3482 786
rect 3056 747 3102 758
rect 3166 726 3278 766
rect 3166 690 3232 726
rect 2944 545 2990 556
rect 2852 453 3186 499
rect 3088 452 3186 453
rect 3088 406 3140 452
rect 2426 256 2431 302
rect 2380 245 2431 256
rect 2718 394 2782 405
rect 2718 348 2736 394
rect 1835 153 2315 199
rect 2604 234 2650 245
rect 2718 242 2782 348
rect 3088 395 3186 406
rect 3088 320 3134 395
rect 3088 263 3134 274
rect 3232 320 3278 586
rect 2604 90 2650 188
rect 3232 169 3278 180
rect 3456 222 3502 233
rect 0 82 3456 90
rect 3502 82 3584 90
rect 0 -90 3584 82
<< labels >>
flabel metal1 s 133 447 315 542 0 FreeSans 200 0 0 0 CLKN
port 3 nsew clock input
flabel metal1 s 589 462 754 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3166 690 3278 766 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2718 242 2782 405 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 0 918 3584 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 2604 233 2650 245 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 6 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 3232 169 3278 690 1 Q
port 4 nsew default output
rlabel metal1 s 3436 852 3482 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3056 852 3102 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2637 852 2705 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1773 852 1819 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1425 852 1471 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 609 852 655 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 261 852 307 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3436 775 3482 852 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3056 775 3102 852 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1773 775 1819 852 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1425 775 1471 852 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 609 775 655 852 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 261 775 307 852 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3056 747 3102 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1773 747 1819 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1425 747 1471 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 609 747 655 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 261 747 307 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1773 703 1819 747 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1425 703 1471 747 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 609 703 655 747 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 261 703 307 747 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1773 685 1819 703 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 261 685 307 703 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1773 671 1819 685 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1649 233 1695 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 641 233 687 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 245 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 3456 90 3502 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2604 90 2650 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1649 90 1695 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3584 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3584 1008
string GDS_END 1518830
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1509914
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
