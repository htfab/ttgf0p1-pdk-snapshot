magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 352 1206 870
<< pwell >>
rect -86 -86 1206 352
<< metal1 >>
rect 0 724 1120 844
rect 242 657 310 724
rect 108 354 314 430
rect 250 224 314 354
rect 360 224 424 483
rect 472 224 582 483
rect 749 506 795 724
rect 729 60 775 218
rect 914 130 1002 676
rect 0 -60 1120 60
<< obsm1 >>
rect 38 611 106 668
rect 446 611 514 668
rect 38 565 683 611
rect 637 360 683 565
rect 637 292 863 360
rect 38 161 106 207
rect 637 161 683 292
rect 38 115 683 161
<< labels >>
rlabel metal1 s 250 224 314 354 6 A1
port 1 nsew default input
rlabel metal1 s 108 354 314 430 6 A1
port 1 nsew default input
rlabel metal1 s 360 224 424 483 6 A2
port 2 nsew default input
rlabel metal1 s 472 224 582 483 6 A3
port 3 nsew default input
rlabel metal1 s 914 130 1002 676 6 Z
port 4 nsew default output
rlabel metal1 s 749 506 795 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 242 657 310 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 724 1120 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel nwell s -86 352 1206 870 6 VNW
port 6 nsew power bidirectional
rlabel pwell s -86 -86 1206 352 6 VPW
port 7 nsew ground bidirectional
rlabel metal1 s 0 -60 1120 60 8 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 729 60 775 218 6 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1223666
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1220322
<< end >>
