* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__fill_8.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__fill_8 VDD VNW VPW VSS
.ends

