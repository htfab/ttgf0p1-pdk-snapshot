magic
tech gf180mcuD
magscale 1 10
timestamp 1755615451
<< nwell >>
rect -86 680 770 1486
<< nmos >>
rect 120 209 176 584
rect 280 209 336 584
rect 440 209 496 584
<< pmos >>
rect 120 776 176 1191
rect 280 776 336 1191
rect 440 776 496 1191
<< ndiff >>
rect 32 268 120 584
rect 32 222 45 268
rect 91 222 120 268
rect 32 209 120 222
rect 176 209 280 584
rect 336 571 440 584
rect 336 325 365 571
rect 411 325 440 571
rect 336 209 440 325
rect 496 268 620 584
rect 496 222 561 268
rect 607 222 620 268
rect 496 209 620 222
<< pdiff >>
rect 32 1055 120 1191
rect 32 809 45 1055
rect 91 809 120 1055
rect 32 776 120 809
rect 176 1178 280 1191
rect 176 1132 205 1178
rect 251 1132 280 1178
rect 176 776 280 1132
rect 336 1055 440 1191
rect 336 809 365 1055
rect 411 809 440 1055
rect 336 776 440 809
rect 496 1055 620 1191
rect 496 809 561 1055
rect 607 809 620 1055
rect 496 776 620 809
<< ndiffc >>
rect 45 222 91 268
rect 365 325 411 571
rect 561 222 607 268
<< pdiffc >>
rect 45 809 91 1055
rect 205 1132 251 1178
rect 365 809 411 1055
rect 561 809 607 1055
<< psubdiff >>
rect 28 87 656 100
rect 28 41 69 87
rect 615 41 656 87
rect 28 28 656 41
<< nsubdiff >>
rect 28 1359 656 1372
rect 28 1313 69 1359
rect 615 1313 656 1359
rect 28 1300 656 1313
<< psubdiffcont >>
rect 69 41 615 87
<< nsubdiffcont >>
rect 69 1313 615 1359
<< polysilicon >>
rect 120 1191 176 1235
rect 280 1191 336 1235
rect 440 1191 496 1235
rect 120 716 176 776
rect 280 716 336 776
rect 32 703 176 716
rect 32 657 45 703
rect 91 657 176 703
rect 32 644 176 657
rect 224 703 336 716
rect 224 657 237 703
rect 283 657 336 703
rect 224 644 336 657
rect 120 584 176 644
rect 280 584 336 644
rect 440 716 496 776
rect 440 703 522 716
rect 440 657 463 703
rect 509 657 522 703
rect 440 644 522 657
rect 440 584 496 644
rect 120 165 176 209
rect 280 165 336 209
rect 440 165 496 209
<< polycontact >>
rect 45 657 91 703
rect 237 657 283 703
rect 463 657 509 703
<< metal1 >>
rect 0 1359 684 1400
rect 0 1313 69 1359
rect 615 1313 684 1359
rect 0 1178 684 1313
rect 0 1132 205 1178
rect 251 1132 684 1178
rect 45 1055 411 1086
rect 91 809 365 1055
rect 45 798 411 809
rect 42 703 94 752
rect 42 657 45 703
rect 91 657 94 703
rect 42 314 94 657
rect 234 703 286 752
rect 234 657 237 703
rect 283 657 286 703
rect 234 314 286 657
rect 460 703 512 1086
rect 460 657 463 703
rect 509 657 512 703
rect 460 628 512 657
rect 558 1055 610 1086
rect 558 809 561 1055
rect 607 809 610 1055
rect 558 582 610 809
rect 365 571 610 582
rect 411 325 610 571
rect 365 314 610 325
rect 0 222 45 268
rect 91 222 561 268
rect 607 222 684 268
rect 0 87 684 222
rect 0 41 69 87
rect 615 41 684 87
rect 0 0 684 41
<< labels >>
rlabel metal1 s 0 0 684 268 4 vss
port 3 nsew
rlabel metal1 s 0 1132 684 1400 4 vdd
port 5 nsew
rlabel metal1 s 42 314 94 752 4 i0
port 7 nsew
rlabel metal1 s 558 314 610 1086 4 nq
port 9 nsew
rlabel metal1 s 234 314 286 752 4 i1
port 11 nsew
rlabel metal1 s 460 628 512 1086 4 i2
port 13 nsew
<< end >>
