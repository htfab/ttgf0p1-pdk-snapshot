VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO and4_x1
  CLASS BLOCK ;
  FOREIGN and4_x1 ;
  ORIGIN 0.430 0.000 ;
  SIZE 6.560 BY 7.430 ;
  PIN vdd
    ANTENNADIFFAREA 3.973000 ;
    PORT
      LAYER Nwell ;
        RECT -0.430 3.400 6.130 7.430 ;
      LAYER Metal1 ;
        RECT 0.000 5.660 5.700 7.000 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 3.040200 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 5.700 1.340 ;
    END
  END vss
  PIN i0
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 0.210 2.140 0.470 5.430 ;
    END
  END i0
  PIN i1
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.170 2.140 1.430 4.860 ;
    END
  END i1
  PIN i2
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.970 2.140 2.230 4.860 ;
    END
  END i2
  PIN i3
    ANTENNAGATEAREA 0.492800 ;
    PORT
      LAYER Metal1 ;
        RECT 2.770 2.140 3.030 4.860 ;
    END
  END i3
  PIN q
    ANTENNADIFFAREA 1.738000 ;
    PORT
      LAYER Metal1 ;
        RECT 4.430 1.570 4.690 5.430 ;
    END
  END q
  OBS
      LAYER Metal1 ;
        RECT 1.025 5.090 3.830 5.430 ;
        RECT 3.570 1.910 3.830 5.090 ;
        RECT 0.225 1.570 3.830 1.910 ;
  END
END and4_x1
END LIBRARY

