* NGSPICE file created from gf180mcu_as_sc_mcu7t3v3__maj3_2.ext - technology: gf180mcuD

.subckt gf180mcu_as_sc_mcu7t3v3__maj3_2 VDD VNW VPW VSS Y A B C
X0 a_436_68# B VSS VPW nfet_03v3 ad=0.12p pd=1.24u as=0.26p ps=1.52u w=1u l=0.28u
X1 VSS A a_700_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.28u
X2 Y a_28_68# VDD VNW pfet_03v3 ad=0.4485p pd=2.03u as=0.3588p ps=1.9u w=1.38u l=0.28u
X3 a_172_68# A a_28_68# VPW nfet_03v3 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.28u
X4 VSS a_28_68# Y VPW nfet_03v3 ad=0.83p pd=3.66u as=0.325p ps=1.65u w=1u l=0.28u
X5 VSS B a_172_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.28u
X6 VDD B a_172_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.1656p ps=1.62u w=1.38u l=0.28u
X7 a_700_440# C a_28_68# VNW pfet_03v3 ad=0.1656p pd=1.62u as=0.3588p ps=1.9u w=1.38u l=0.28u
X8 a_700_68# C a_28_68# VPW nfet_03v3 ad=0.12p pd=1.24u as=0.26p ps=1.52u w=1u l=0.28u
X9 a_436_440# B VDD VNW pfet_03v3 ad=0.1656p pd=1.62u as=0.3588p ps=1.9u w=1.38u l=0.28u
X10 a_28_68# C a_436_68# VPW nfet_03v3 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.28u
X11 VDD A a_700_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.1656p ps=1.62u w=1.38u l=0.28u
X12 Y a_28_68# VSS VPW nfet_03v3 ad=0.325p pd=1.65u as=0.26p ps=1.52u w=1u l=0.28u
X13 a_28_68# C a_436_440# VNW pfet_03v3 ad=0.3588p pd=1.9u as=0.1656p ps=1.62u w=1.38u l=0.28u
X14 a_172_440# A a_28_68# VNW pfet_03v3 ad=0.1656p pd=1.62u as=0.6072p ps=3.64u w=1.38u l=0.28u
X15 VDD a_28_68# Y VNW pfet_03v3 ad=1.1454p pd=4.42u as=0.4485p ps=2.03u w=1.38u l=0.28u
.ends

