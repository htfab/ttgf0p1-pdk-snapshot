magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< metal1 >>
rect 14757 50970 14833 50982
rect 14757 50918 14769 50970
rect 14821 50918 14833 50970
rect 14757 50862 14833 50918
rect 14757 50810 14769 50862
rect 14821 50810 14833 50862
rect 14757 50754 14833 50810
rect 14757 50702 14769 50754
rect 14821 50702 14833 50754
rect 14757 50646 14833 50702
rect 14757 50594 14769 50646
rect 14821 50594 14833 50646
rect 14757 50538 14833 50594
rect 14757 50486 14769 50538
rect 14821 50486 14833 50538
rect 14757 50430 14833 50486
rect 14757 50378 14769 50430
rect 14821 50378 14833 50430
rect 14757 50322 14833 50378
rect 14757 50270 14769 50322
rect 14821 50270 14833 50322
rect 14757 50214 14833 50270
rect 14757 50162 14769 50214
rect 14821 50162 14833 50214
rect 14757 50106 14833 50162
rect 14757 50054 14769 50106
rect 14821 50054 14833 50106
rect 14757 49998 14833 50054
rect 14757 49946 14769 49998
rect 14821 49946 14833 49998
rect 14757 49890 14833 49946
rect 14757 49838 14769 49890
rect 14821 49838 14833 49890
rect 14757 49782 14833 49838
rect 14757 49730 14769 49782
rect 14821 49730 14833 49782
rect 14757 49674 14833 49730
rect 14757 49622 14769 49674
rect 14821 49622 14833 49674
rect 14757 49610 14833 49622
rect 14757 36570 14833 36582
rect 14757 36518 14769 36570
rect 14821 36518 14833 36570
rect 14757 36462 14833 36518
rect 14757 36410 14769 36462
rect 14821 36410 14833 36462
rect 14757 36354 14833 36410
rect 14757 36302 14769 36354
rect 14821 36302 14833 36354
rect 14757 36246 14833 36302
rect 14757 36194 14769 36246
rect 14821 36194 14833 36246
rect 14757 36138 14833 36194
rect 14757 36086 14769 36138
rect 14821 36086 14833 36138
rect 14757 36030 14833 36086
rect 14757 35978 14769 36030
rect 14821 35978 14833 36030
rect 14757 35922 14833 35978
rect 14757 35870 14769 35922
rect 14821 35870 14833 35922
rect 14757 35814 14833 35870
rect 14757 35762 14769 35814
rect 14821 35762 14833 35814
rect 14757 35706 14833 35762
rect 14757 35654 14769 35706
rect 14821 35654 14833 35706
rect 14757 35598 14833 35654
rect 14757 35546 14769 35598
rect 14821 35546 14833 35598
rect 14757 35490 14833 35546
rect 14757 35438 14769 35490
rect 14821 35438 14833 35490
rect 14757 35382 14833 35438
rect 14757 35330 14769 35382
rect 14821 35330 14833 35382
rect 14757 35274 14833 35330
rect 14757 35222 14769 35274
rect 14821 35222 14833 35274
rect 14757 35210 14833 35222
<< via1 >>
rect 14769 50918 14821 50970
rect 14769 50810 14821 50862
rect 14769 50702 14821 50754
rect 14769 50594 14821 50646
rect 14769 50486 14821 50538
rect 14769 50378 14821 50430
rect 14769 50270 14821 50322
rect 14769 50162 14821 50214
rect 14769 50054 14821 50106
rect 14769 49946 14821 49998
rect 14769 49838 14821 49890
rect 14769 49730 14821 49782
rect 14769 49622 14821 49674
rect 14769 36518 14821 36570
rect 14769 36410 14821 36462
rect 14769 36302 14821 36354
rect 14769 36194 14821 36246
rect 14769 36086 14821 36138
rect 14769 35978 14821 36030
rect 14769 35870 14821 35922
rect 14769 35762 14821 35814
rect 14769 35654 14821 35706
rect 14769 35546 14821 35598
rect 14769 35438 14821 35490
rect 14769 35330 14821 35382
rect 14769 35222 14821 35274
<< metal2 >>
rect 14757 50972 14833 50982
rect 14757 49620 14767 50972
rect 14823 49620 14833 50972
rect 14757 49610 14833 49620
rect 6384 46670 6460 46680
rect 6384 46614 6394 46670
rect 6450 46614 6460 46670
rect 6384 46546 6460 46614
rect 6384 46490 6394 46546
rect 6450 46490 6460 46546
rect 6384 46422 6460 46490
rect 6384 46366 6394 46422
rect 6450 46366 6460 46422
rect 4460 46323 4536 46333
rect 4460 46267 4470 46323
rect 4526 46267 4536 46323
rect 4460 46199 4536 46267
rect 6384 46298 6460 46366
rect 6384 46242 6394 46298
rect 6450 46242 6460 46298
rect 4460 46143 4470 46199
rect 4526 46143 4536 46199
rect 4460 46075 4536 46143
rect 4460 46019 4470 46075
rect 4526 46019 4536 46075
rect 4460 45951 4536 46019
rect 4460 45895 4470 45951
rect 4526 45895 4536 45951
rect 4460 45827 4536 45895
rect 4460 45771 4470 45827
rect 4526 45771 4536 45827
rect 4460 45703 4536 45771
rect 4460 45647 4470 45703
rect 4526 45647 4536 45703
rect 4460 45579 4536 45647
rect 4460 45523 4470 45579
rect 4526 45523 4536 45579
rect 4460 45455 4536 45523
rect 4460 45399 4470 45455
rect 4526 45399 4536 45455
rect 4460 45331 4536 45399
rect 4460 45275 4470 45331
rect 4526 45275 4536 45331
rect 1094 45255 1170 45265
rect 1094 45199 1104 45255
rect 1160 45199 1170 45255
rect 1094 45131 1170 45199
rect 4460 45207 4536 45275
rect 4460 45151 4470 45207
rect 4526 45151 4536 45207
rect 1094 45075 1104 45131
rect 1160 45075 1170 45131
rect 1094 45007 1170 45075
rect 1094 44951 1104 45007
rect 1160 44951 1170 45007
rect 1094 44883 1170 44951
rect 1094 44827 1104 44883
rect 1160 44827 1170 44883
rect 1094 44759 1170 44827
rect 1094 44703 1104 44759
rect 1160 44703 1170 44759
rect 1094 44635 1170 44703
rect 1094 44579 1104 44635
rect 1160 44579 1170 44635
rect 1094 44511 1170 44579
rect 1094 44455 1104 44511
rect 1160 44455 1170 44511
rect 1094 44387 1170 44455
rect 1094 44331 1104 44387
rect 1160 44331 1170 44387
rect 1094 44263 1170 44331
rect 1094 44207 1104 44263
rect 1160 44207 1170 44263
rect 1094 44139 1170 44207
rect 1094 44083 1104 44139
rect 1160 44083 1170 44139
rect 1094 44015 1170 44083
rect 1094 43959 1104 44015
rect 1160 43959 1170 44015
rect 1094 43891 1170 43959
rect 1094 43835 1104 43891
rect 1160 43835 1170 43891
rect 1094 43767 1170 43835
rect 1094 43711 1104 43767
rect 1160 43711 1170 43767
rect 1094 43643 1170 43711
rect 1094 43587 1104 43643
rect 1160 43587 1170 43643
rect 1094 43519 1170 43587
rect 1094 43463 1104 43519
rect 1160 43463 1170 43519
rect 1094 43453 1170 43463
rect 1218 45131 1294 45141
rect 1218 45075 1228 45131
rect 1284 45075 1294 45131
rect 1218 45007 1294 45075
rect 4460 45083 4536 45151
rect 4460 45027 4470 45083
rect 4526 45027 4536 45083
rect 1218 44951 1228 45007
rect 1284 44951 1294 45007
rect 1218 44883 1294 44951
rect 1218 44827 1228 44883
rect 1284 44827 1294 44883
rect 1218 44759 1294 44827
rect 1218 44703 1228 44759
rect 1284 44703 1294 44759
rect 1218 44635 1294 44703
rect 1218 44579 1228 44635
rect 1284 44579 1294 44635
rect 1218 44511 1294 44579
rect 1218 44455 1228 44511
rect 1284 44455 1294 44511
rect 1218 44387 1294 44455
rect 1218 44331 1228 44387
rect 1284 44331 1294 44387
rect 1218 44263 1294 44331
rect 1218 44207 1228 44263
rect 1284 44207 1294 44263
rect 1218 44139 1294 44207
rect 1218 44083 1228 44139
rect 1284 44083 1294 44139
rect 1218 44015 1294 44083
rect 1218 43959 1228 44015
rect 1284 43959 1294 44015
rect 1218 43891 1294 43959
rect 1218 43835 1228 43891
rect 1284 43835 1294 43891
rect 1218 43767 1294 43835
rect 1218 43711 1228 43767
rect 1284 43711 1294 43767
rect 1218 43643 1294 43711
rect 1218 43587 1228 43643
rect 1284 43587 1294 43643
rect 1218 43519 1294 43587
rect 1218 43463 1228 43519
rect 1284 43463 1294 43519
rect 1218 43395 1294 43463
rect 1218 43339 1228 43395
rect 1284 43339 1294 43395
rect 1218 43329 1294 43339
rect 1342 45007 1418 45017
rect 1342 44951 1352 45007
rect 1408 44951 1418 45007
rect 1342 44883 1418 44951
rect 4460 44959 4536 45027
rect 4460 44903 4470 44959
rect 4526 44903 4536 44959
rect 1342 44827 1352 44883
rect 1408 44827 1418 44883
rect 1342 44759 1418 44827
rect 1342 44703 1352 44759
rect 1408 44703 1418 44759
rect 1342 44635 1418 44703
rect 1342 44579 1352 44635
rect 1408 44579 1418 44635
rect 1342 44511 1418 44579
rect 1342 44455 1352 44511
rect 1408 44455 1418 44511
rect 1342 44387 1418 44455
rect 1342 44331 1352 44387
rect 1408 44331 1418 44387
rect 1342 44263 1418 44331
rect 1342 44207 1352 44263
rect 1408 44207 1418 44263
rect 1342 44139 1418 44207
rect 1342 44083 1352 44139
rect 1408 44083 1418 44139
rect 1342 44015 1418 44083
rect 1342 43959 1352 44015
rect 1408 43959 1418 44015
rect 1342 43891 1418 43959
rect 1342 43835 1352 43891
rect 1408 43835 1418 43891
rect 1342 43767 1418 43835
rect 1342 43711 1352 43767
rect 1408 43711 1418 43767
rect 1342 43643 1418 43711
rect 1342 43587 1352 43643
rect 1408 43587 1418 43643
rect 1342 43519 1418 43587
rect 1342 43463 1352 43519
rect 1408 43463 1418 43519
rect 1342 43395 1418 43463
rect 1342 43339 1352 43395
rect 1408 43339 1418 43395
rect 1342 43271 1418 43339
rect 1342 43215 1352 43271
rect 1408 43215 1418 43271
rect 1342 43205 1418 43215
rect 1466 44883 1542 44893
rect 1466 44827 1476 44883
rect 1532 44827 1542 44883
rect 1466 44759 1542 44827
rect 4460 44835 4536 44903
rect 4460 44779 4470 44835
rect 4526 44779 4536 44835
rect 1466 44703 1476 44759
rect 1532 44703 1542 44759
rect 1466 44635 1542 44703
rect 1466 44579 1476 44635
rect 1532 44579 1542 44635
rect 1466 44511 1542 44579
rect 1466 44455 1476 44511
rect 1532 44455 1542 44511
rect 1466 44387 1542 44455
rect 1466 44331 1476 44387
rect 1532 44331 1542 44387
rect 1466 44263 1542 44331
rect 1466 44207 1476 44263
rect 1532 44207 1542 44263
rect 1466 44139 1542 44207
rect 1466 44083 1476 44139
rect 1532 44083 1542 44139
rect 1466 44015 1542 44083
rect 1466 43959 1476 44015
rect 1532 43959 1542 44015
rect 1466 43891 1542 43959
rect 1466 43835 1476 43891
rect 1532 43835 1542 43891
rect 1466 43767 1542 43835
rect 1466 43711 1476 43767
rect 1532 43711 1542 43767
rect 1466 43643 1542 43711
rect 1466 43587 1476 43643
rect 1532 43587 1542 43643
rect 1466 43519 1542 43587
rect 1466 43463 1476 43519
rect 1532 43463 1542 43519
rect 1466 43395 1542 43463
rect 1466 43339 1476 43395
rect 1532 43339 1542 43395
rect 1466 43271 1542 43339
rect 1466 43215 1476 43271
rect 1532 43215 1542 43271
rect 1466 43147 1542 43215
rect 1466 43091 1476 43147
rect 1532 43091 1542 43147
rect 1466 43081 1542 43091
rect 1590 44759 1666 44769
rect 1590 44703 1600 44759
rect 1656 44703 1666 44759
rect 1590 44635 1666 44703
rect 4460 44711 4536 44779
rect 4460 44655 4470 44711
rect 4526 44655 4536 44711
rect 4460 44645 4536 44655
rect 4584 46199 4660 46209
rect 4584 46143 4594 46199
rect 4650 46143 4660 46199
rect 4584 46075 4660 46143
rect 6384 46174 6460 46242
rect 6384 46118 6394 46174
rect 6450 46118 6460 46174
rect 4584 46019 4594 46075
rect 4650 46019 4660 46075
rect 4584 45951 4660 46019
rect 4584 45895 4594 45951
rect 4650 45895 4660 45951
rect 4584 45827 4660 45895
rect 4584 45771 4594 45827
rect 4650 45771 4660 45827
rect 4584 45703 4660 45771
rect 4584 45647 4594 45703
rect 4650 45647 4660 45703
rect 4584 45579 4660 45647
rect 4584 45523 4594 45579
rect 4650 45523 4660 45579
rect 4584 45455 4660 45523
rect 4584 45399 4594 45455
rect 4650 45399 4660 45455
rect 4584 45331 4660 45399
rect 4584 45275 4594 45331
rect 4650 45275 4660 45331
rect 4584 45207 4660 45275
rect 4584 45151 4594 45207
rect 4650 45151 4660 45207
rect 4584 45083 4660 45151
rect 4584 45027 4594 45083
rect 4650 45027 4660 45083
rect 4584 44959 4660 45027
rect 4584 44903 4594 44959
rect 4650 44903 4660 44959
rect 4584 44835 4660 44903
rect 4584 44779 4594 44835
rect 4650 44779 4660 44835
rect 4584 44711 4660 44779
rect 4584 44655 4594 44711
rect 4650 44655 4660 44711
rect 1590 44579 1600 44635
rect 1656 44579 1666 44635
rect 1590 44511 1666 44579
rect 1590 44455 1600 44511
rect 1656 44455 1666 44511
rect 1590 44387 1666 44455
rect 1590 44331 1600 44387
rect 1656 44331 1666 44387
rect 1590 44263 1666 44331
rect 1590 44207 1600 44263
rect 1656 44207 1666 44263
rect 1590 44139 1666 44207
rect 1590 44083 1600 44139
rect 1656 44083 1666 44139
rect 1590 44015 1666 44083
rect 1590 43959 1600 44015
rect 1656 43959 1666 44015
rect 1590 43891 1666 43959
rect 1590 43835 1600 43891
rect 1656 43835 1666 43891
rect 1590 43767 1666 43835
rect 1590 43711 1600 43767
rect 1656 43711 1666 43767
rect 1590 43643 1666 43711
rect 1590 43587 1600 43643
rect 1656 43587 1666 43643
rect 1590 43519 1666 43587
rect 1590 43463 1600 43519
rect 1656 43463 1666 43519
rect 1590 43395 1666 43463
rect 1590 43339 1600 43395
rect 1656 43339 1666 43395
rect 1590 43271 1666 43339
rect 1590 43215 1600 43271
rect 1656 43215 1666 43271
rect 1590 43147 1666 43215
rect 1590 43091 1600 43147
rect 1656 43091 1666 43147
rect 1590 43023 1666 43091
rect 1590 42967 1600 43023
rect 1656 42967 1666 43023
rect 1590 42957 1666 42967
rect 1714 44635 1790 44645
rect 1714 44579 1724 44635
rect 1780 44579 1790 44635
rect 1714 44511 1790 44579
rect 4584 44587 4660 44655
rect 4584 44531 4594 44587
rect 4650 44531 4660 44587
rect 4584 44521 4660 44531
rect 4708 46075 4784 46085
rect 4708 46019 4718 46075
rect 4774 46019 4784 46075
rect 4708 45951 4784 46019
rect 6384 46050 6460 46118
rect 6384 45994 6394 46050
rect 6450 45994 6460 46050
rect 4708 45895 4718 45951
rect 4774 45895 4784 45951
rect 4708 45827 4784 45895
rect 4708 45771 4718 45827
rect 4774 45771 4784 45827
rect 4708 45703 4784 45771
rect 4708 45647 4718 45703
rect 4774 45647 4784 45703
rect 4708 45579 4784 45647
rect 4708 45523 4718 45579
rect 4774 45523 4784 45579
rect 4708 45455 4784 45523
rect 4708 45399 4718 45455
rect 4774 45399 4784 45455
rect 4708 45331 4784 45399
rect 4708 45275 4718 45331
rect 4774 45275 4784 45331
rect 4708 45207 4784 45275
rect 4708 45151 4718 45207
rect 4774 45151 4784 45207
rect 4708 45083 4784 45151
rect 4708 45027 4718 45083
rect 4774 45027 4784 45083
rect 4708 44959 4784 45027
rect 4708 44903 4718 44959
rect 4774 44903 4784 44959
rect 4708 44835 4784 44903
rect 4708 44779 4718 44835
rect 4774 44779 4784 44835
rect 4708 44711 4784 44779
rect 4708 44655 4718 44711
rect 4774 44655 4784 44711
rect 4708 44587 4784 44655
rect 4708 44531 4718 44587
rect 4774 44531 4784 44587
rect 1714 44455 1724 44511
rect 1780 44455 1790 44511
rect 1714 44387 1790 44455
rect 1714 44331 1724 44387
rect 1780 44331 1790 44387
rect 1714 44263 1790 44331
rect 1714 44207 1724 44263
rect 1780 44207 1790 44263
rect 1714 44139 1790 44207
rect 1714 44083 1724 44139
rect 1780 44083 1790 44139
rect 1714 44015 1790 44083
rect 1714 43959 1724 44015
rect 1780 43959 1790 44015
rect 1714 43891 1790 43959
rect 1714 43835 1724 43891
rect 1780 43835 1790 43891
rect 1714 43767 1790 43835
rect 1714 43711 1724 43767
rect 1780 43711 1790 43767
rect 1714 43643 1790 43711
rect 1714 43587 1724 43643
rect 1780 43587 1790 43643
rect 1714 43519 1790 43587
rect 1714 43463 1724 43519
rect 1780 43463 1790 43519
rect 1714 43395 1790 43463
rect 1714 43339 1724 43395
rect 1780 43339 1790 43395
rect 1714 43271 1790 43339
rect 1714 43215 1724 43271
rect 1780 43215 1790 43271
rect 1714 43147 1790 43215
rect 1714 43091 1724 43147
rect 1780 43091 1790 43147
rect 1714 43023 1790 43091
rect 1714 42967 1724 43023
rect 1780 42967 1790 43023
rect 1714 42899 1790 42967
rect 1714 42843 1724 42899
rect 1780 42843 1790 42899
rect 1714 42833 1790 42843
rect 1838 44511 1914 44521
rect 1838 44455 1848 44511
rect 1904 44455 1914 44511
rect 1838 44387 1914 44455
rect 4708 44463 4784 44531
rect 4708 44407 4718 44463
rect 4774 44407 4784 44463
rect 4708 44397 4784 44407
rect 4832 45951 4908 45961
rect 4832 45895 4842 45951
rect 4898 45895 4908 45951
rect 4832 45827 4908 45895
rect 6384 45926 6460 45994
rect 6384 45870 6394 45926
rect 6450 45870 6460 45926
rect 4832 45771 4842 45827
rect 4898 45771 4908 45827
rect 4832 45703 4908 45771
rect 4832 45647 4842 45703
rect 4898 45647 4908 45703
rect 4832 45579 4908 45647
rect 4832 45523 4842 45579
rect 4898 45523 4908 45579
rect 4832 45455 4908 45523
rect 4832 45399 4842 45455
rect 4898 45399 4908 45455
rect 4832 45331 4908 45399
rect 4832 45275 4842 45331
rect 4898 45275 4908 45331
rect 4832 45207 4908 45275
rect 4832 45151 4842 45207
rect 4898 45151 4908 45207
rect 4832 45083 4908 45151
rect 4832 45027 4842 45083
rect 4898 45027 4908 45083
rect 4832 44959 4908 45027
rect 4832 44903 4842 44959
rect 4898 44903 4908 44959
rect 4832 44835 4908 44903
rect 4832 44779 4842 44835
rect 4898 44779 4908 44835
rect 4832 44711 4908 44779
rect 4832 44655 4842 44711
rect 4898 44655 4908 44711
rect 4832 44587 4908 44655
rect 4832 44531 4842 44587
rect 4898 44531 4908 44587
rect 4832 44463 4908 44531
rect 4832 44407 4842 44463
rect 4898 44407 4908 44463
rect 1838 44331 1848 44387
rect 1904 44331 1914 44387
rect 1838 44263 1914 44331
rect 1838 44207 1848 44263
rect 1904 44207 1914 44263
rect 1838 44139 1914 44207
rect 1838 44083 1848 44139
rect 1904 44083 1914 44139
rect 1838 44015 1914 44083
rect 1838 43959 1848 44015
rect 1904 43959 1914 44015
rect 1838 43891 1914 43959
rect 1838 43835 1848 43891
rect 1904 43835 1914 43891
rect 1838 43767 1914 43835
rect 1838 43711 1848 43767
rect 1904 43711 1914 43767
rect 1838 43643 1914 43711
rect 1838 43587 1848 43643
rect 1904 43587 1914 43643
rect 1838 43519 1914 43587
rect 1838 43463 1848 43519
rect 1904 43463 1914 43519
rect 1838 43395 1914 43463
rect 1838 43339 1848 43395
rect 1904 43339 1914 43395
rect 1838 43271 1914 43339
rect 1838 43215 1848 43271
rect 1904 43215 1914 43271
rect 1838 43147 1914 43215
rect 1838 43091 1848 43147
rect 1904 43091 1914 43147
rect 1838 43023 1914 43091
rect 1838 42967 1848 43023
rect 1904 42967 1914 43023
rect 1838 42899 1914 42967
rect 1838 42843 1848 42899
rect 1904 42843 1914 42899
rect 1838 42775 1914 42843
rect 1838 42719 1848 42775
rect 1904 42719 1914 42775
rect 1838 42709 1914 42719
rect 1962 44387 2038 44397
rect 1962 44331 1972 44387
rect 2028 44331 2038 44387
rect 1962 44263 2038 44331
rect 4832 44339 4908 44407
rect 4832 44283 4842 44339
rect 4898 44283 4908 44339
rect 4832 44273 4908 44283
rect 4956 45827 5032 45837
rect 4956 45771 4966 45827
rect 5022 45771 5032 45827
rect 4956 45703 5032 45771
rect 6384 45802 6460 45870
rect 6384 45746 6394 45802
rect 6450 45746 6460 45802
rect 4956 45647 4966 45703
rect 5022 45647 5032 45703
rect 4956 45579 5032 45647
rect 4956 45523 4966 45579
rect 5022 45523 5032 45579
rect 4956 45455 5032 45523
rect 4956 45399 4966 45455
rect 5022 45399 5032 45455
rect 4956 45331 5032 45399
rect 4956 45275 4966 45331
rect 5022 45275 5032 45331
rect 4956 45207 5032 45275
rect 4956 45151 4966 45207
rect 5022 45151 5032 45207
rect 4956 45083 5032 45151
rect 4956 45027 4966 45083
rect 5022 45027 5032 45083
rect 4956 44959 5032 45027
rect 4956 44903 4966 44959
rect 5022 44903 5032 44959
rect 4956 44835 5032 44903
rect 4956 44779 4966 44835
rect 5022 44779 5032 44835
rect 4956 44711 5032 44779
rect 4956 44655 4966 44711
rect 5022 44655 5032 44711
rect 4956 44587 5032 44655
rect 4956 44531 4966 44587
rect 5022 44531 5032 44587
rect 4956 44463 5032 44531
rect 4956 44407 4966 44463
rect 5022 44407 5032 44463
rect 4956 44339 5032 44407
rect 4956 44283 4966 44339
rect 5022 44283 5032 44339
rect 1962 44207 1972 44263
rect 2028 44207 2038 44263
rect 1962 44139 2038 44207
rect 4956 44215 5032 44283
rect 4956 44159 4966 44215
rect 5022 44159 5032 44215
rect 4956 44149 5032 44159
rect 5080 45703 5156 45713
rect 5080 45647 5090 45703
rect 5146 45647 5156 45703
rect 5080 45579 5156 45647
rect 6384 45678 6460 45746
rect 6384 45622 6394 45678
rect 6450 45622 6460 45678
rect 5080 45523 5090 45579
rect 5146 45523 5156 45579
rect 5080 45455 5156 45523
rect 5080 45399 5090 45455
rect 5146 45399 5156 45455
rect 5080 45331 5156 45399
rect 5080 45275 5090 45331
rect 5146 45275 5156 45331
rect 5080 45207 5156 45275
rect 5080 45151 5090 45207
rect 5146 45151 5156 45207
rect 5080 45083 5156 45151
rect 5080 45027 5090 45083
rect 5146 45027 5156 45083
rect 5080 44959 5156 45027
rect 5080 44903 5090 44959
rect 5146 44903 5156 44959
rect 5080 44835 5156 44903
rect 5080 44779 5090 44835
rect 5146 44779 5156 44835
rect 5080 44711 5156 44779
rect 5080 44655 5090 44711
rect 5146 44655 5156 44711
rect 5080 44587 5156 44655
rect 5080 44531 5090 44587
rect 5146 44531 5156 44587
rect 5080 44463 5156 44531
rect 5080 44407 5090 44463
rect 5146 44407 5156 44463
rect 5080 44339 5156 44407
rect 5080 44283 5090 44339
rect 5146 44283 5156 44339
rect 5080 44215 5156 44283
rect 5080 44159 5090 44215
rect 5146 44159 5156 44215
rect 1962 44083 1972 44139
rect 2028 44083 2038 44139
rect 1962 44015 2038 44083
rect 5080 44091 5156 44159
rect 5080 44035 5090 44091
rect 5146 44035 5156 44091
rect 1962 43959 1972 44015
rect 2028 43959 2038 44015
rect 1962 43891 2038 43959
rect 1962 43835 1972 43891
rect 2028 43835 2038 43891
rect 1962 43767 2038 43835
rect 1962 43711 1972 43767
rect 2028 43711 2038 43767
rect 1962 43643 2038 43711
rect 1962 43587 1972 43643
rect 2028 43587 2038 43643
rect 1962 43519 2038 43587
rect 1962 43463 1972 43519
rect 2028 43463 2038 43519
rect 1962 43395 2038 43463
rect 1962 43339 1972 43395
rect 2028 43339 2038 43395
rect 1962 43271 2038 43339
rect 1962 43215 1972 43271
rect 2028 43215 2038 43271
rect 1962 43147 2038 43215
rect 1962 43091 1972 43147
rect 2028 43091 2038 43147
rect 1962 43023 2038 43091
rect 1962 42967 1972 43023
rect 2028 42967 2038 43023
rect 1962 42899 2038 42967
rect 1962 42843 1972 42899
rect 2028 42843 2038 42899
rect 1962 42775 2038 42843
rect 1962 42719 1972 42775
rect 2028 42719 2038 42775
rect 1962 42651 2038 42719
rect 1962 42595 1972 42651
rect 2028 42595 2038 42651
rect 1962 42585 2038 42595
rect 4460 44024 4536 44034
rect 5080 44025 5156 44035
rect 5204 45579 5280 45589
rect 5204 45523 5214 45579
rect 5270 45523 5280 45579
rect 5204 45455 5280 45523
rect 6384 45554 6460 45622
rect 6384 45498 6394 45554
rect 6450 45498 6460 45554
rect 5204 45399 5214 45455
rect 5270 45399 5280 45455
rect 5204 45331 5280 45399
rect 5204 45275 5214 45331
rect 5270 45275 5280 45331
rect 5204 45207 5280 45275
rect 5204 45151 5214 45207
rect 5270 45151 5280 45207
rect 5204 45083 5280 45151
rect 5204 45027 5214 45083
rect 5270 45027 5280 45083
rect 5204 44959 5280 45027
rect 5204 44903 5214 44959
rect 5270 44903 5280 44959
rect 5204 44835 5280 44903
rect 5204 44779 5214 44835
rect 5270 44779 5280 44835
rect 5204 44711 5280 44779
rect 5204 44655 5214 44711
rect 5270 44655 5280 44711
rect 5204 44587 5280 44655
rect 5204 44531 5214 44587
rect 5270 44531 5280 44587
rect 5204 44463 5280 44531
rect 5204 44407 5214 44463
rect 5270 44407 5280 44463
rect 5204 44339 5280 44407
rect 5204 44283 5214 44339
rect 5270 44283 5280 44339
rect 5204 44215 5280 44283
rect 5204 44159 5214 44215
rect 5270 44159 5280 44215
rect 5204 44091 5280 44159
rect 5204 44035 5214 44091
rect 5270 44035 5280 44091
rect 4460 43968 4470 44024
rect 4526 43968 4536 44024
rect 4460 43900 4536 43968
rect 5204 43967 5280 44035
rect 5204 43911 5214 43967
rect 5270 43911 5280 43967
rect 4460 43844 4470 43900
rect 4526 43844 4536 43900
rect 4460 43776 4536 43844
rect 4460 43720 4470 43776
rect 4526 43720 4536 43776
rect 4460 43652 4536 43720
rect 4460 43596 4470 43652
rect 4526 43596 4536 43652
rect 4460 43528 4536 43596
rect 4460 43472 4470 43528
rect 4526 43472 4536 43528
rect 4460 43404 4536 43472
rect 4460 43348 4470 43404
rect 4526 43348 4536 43404
rect 4460 43280 4536 43348
rect 4460 43224 4470 43280
rect 4526 43224 4536 43280
rect 4460 43156 4536 43224
rect 4460 43100 4470 43156
rect 4526 43100 4536 43156
rect 4460 43032 4536 43100
rect 4460 42976 4470 43032
rect 4526 42976 4536 43032
rect 4460 42908 4536 42976
rect 4460 42852 4470 42908
rect 4526 42852 4536 42908
rect 4460 42784 4536 42852
rect 4460 42728 4470 42784
rect 4526 42728 4536 42784
rect 4460 42660 4536 42728
rect 4460 42604 4470 42660
rect 4526 42604 4536 42660
rect 4460 42536 4536 42604
rect 4460 42480 4470 42536
rect 4526 42480 4536 42536
rect 4460 42412 4536 42480
rect 4460 42356 4470 42412
rect 4526 42356 4536 42412
rect 4460 42346 4536 42356
rect 4584 43900 4660 43910
rect 5204 43901 5280 43911
rect 5328 45455 5404 45465
rect 5328 45399 5338 45455
rect 5394 45399 5404 45455
rect 5328 45331 5404 45399
rect 6384 45430 6460 45498
rect 6384 45374 6394 45430
rect 6450 45374 6460 45430
rect 5328 45275 5338 45331
rect 5394 45275 5404 45331
rect 5328 45207 5404 45275
rect 5328 45151 5338 45207
rect 5394 45151 5404 45207
rect 5328 45083 5404 45151
rect 5328 45027 5338 45083
rect 5394 45027 5404 45083
rect 5328 44959 5404 45027
rect 5328 44903 5338 44959
rect 5394 44903 5404 44959
rect 5328 44835 5404 44903
rect 5328 44779 5338 44835
rect 5394 44779 5404 44835
rect 5328 44711 5404 44779
rect 5328 44655 5338 44711
rect 5394 44655 5404 44711
rect 5328 44587 5404 44655
rect 5328 44531 5338 44587
rect 5394 44531 5404 44587
rect 5328 44463 5404 44531
rect 5328 44407 5338 44463
rect 5394 44407 5404 44463
rect 5328 44339 5404 44407
rect 5328 44283 5338 44339
rect 5394 44283 5404 44339
rect 5328 44215 5404 44283
rect 5328 44159 5338 44215
rect 5394 44159 5404 44215
rect 5328 44091 5404 44159
rect 5328 44035 5338 44091
rect 5394 44035 5404 44091
rect 5328 43967 5404 44035
rect 5328 43911 5338 43967
rect 5394 43911 5404 43967
rect 4584 43844 4594 43900
rect 4650 43844 4660 43900
rect 4584 43776 4660 43844
rect 5328 43843 5404 43911
rect 5328 43787 5338 43843
rect 5394 43787 5404 43843
rect 4584 43720 4594 43776
rect 4650 43720 4660 43776
rect 4584 43652 4660 43720
rect 4584 43596 4594 43652
rect 4650 43596 4660 43652
rect 4584 43528 4660 43596
rect 4584 43472 4594 43528
rect 4650 43472 4660 43528
rect 4584 43404 4660 43472
rect 4584 43348 4594 43404
rect 4650 43348 4660 43404
rect 4584 43280 4660 43348
rect 4584 43224 4594 43280
rect 4650 43224 4660 43280
rect 4584 43156 4660 43224
rect 4584 43100 4594 43156
rect 4650 43100 4660 43156
rect 4584 43032 4660 43100
rect 4584 42976 4594 43032
rect 4650 42976 4660 43032
rect 4584 42908 4660 42976
rect 4584 42852 4594 42908
rect 4650 42852 4660 42908
rect 4584 42784 4660 42852
rect 4584 42728 4594 42784
rect 4650 42728 4660 42784
rect 4584 42660 4660 42728
rect 4584 42604 4594 42660
rect 4650 42604 4660 42660
rect 4584 42536 4660 42604
rect 4584 42480 4594 42536
rect 4650 42480 4660 42536
rect 4584 42412 4660 42480
rect 4584 42356 4594 42412
rect 4650 42356 4660 42412
rect 4584 42288 4660 42356
rect 4584 42232 4594 42288
rect 4650 42232 4660 42288
rect 4584 42222 4660 42232
rect 4708 43776 4784 43786
rect 5328 43777 5404 43787
rect 5452 45331 5528 45341
rect 5452 45275 5462 45331
rect 5518 45275 5528 45331
rect 5452 45207 5528 45275
rect 6384 45306 6460 45374
rect 6384 45250 6394 45306
rect 6450 45250 6460 45306
rect 5452 45151 5462 45207
rect 5518 45151 5528 45207
rect 5452 45083 5528 45151
rect 5452 45027 5462 45083
rect 5518 45027 5528 45083
rect 5452 44959 5528 45027
rect 5452 44903 5462 44959
rect 5518 44903 5528 44959
rect 5452 44835 5528 44903
rect 5452 44779 5462 44835
rect 5518 44779 5528 44835
rect 5452 44711 5528 44779
rect 5452 44655 5462 44711
rect 5518 44655 5528 44711
rect 5452 44587 5528 44655
rect 5452 44531 5462 44587
rect 5518 44531 5528 44587
rect 5452 44463 5528 44531
rect 5452 44407 5462 44463
rect 5518 44407 5528 44463
rect 5452 44339 5528 44407
rect 5452 44283 5462 44339
rect 5518 44283 5528 44339
rect 5452 44215 5528 44283
rect 5452 44159 5462 44215
rect 5518 44159 5528 44215
rect 5452 44091 5528 44159
rect 5452 44035 5462 44091
rect 5518 44035 5528 44091
rect 5452 43967 5528 44035
rect 5452 43911 5462 43967
rect 5518 43911 5528 43967
rect 5452 43843 5528 43911
rect 5452 43787 5462 43843
rect 5518 43787 5528 43843
rect 4708 43720 4718 43776
rect 4774 43720 4784 43776
rect 4708 43652 4784 43720
rect 5452 43719 5528 43787
rect 5452 43663 5462 43719
rect 5518 43663 5528 43719
rect 4708 43596 4718 43652
rect 4774 43596 4784 43652
rect 4708 43528 4784 43596
rect 4708 43472 4718 43528
rect 4774 43472 4784 43528
rect 4708 43404 4784 43472
rect 4708 43348 4718 43404
rect 4774 43348 4784 43404
rect 4708 43280 4784 43348
rect 4708 43224 4718 43280
rect 4774 43224 4784 43280
rect 4708 43156 4784 43224
rect 4708 43100 4718 43156
rect 4774 43100 4784 43156
rect 4708 43032 4784 43100
rect 4708 42976 4718 43032
rect 4774 42976 4784 43032
rect 4708 42908 4784 42976
rect 4708 42852 4718 42908
rect 4774 42852 4784 42908
rect 4708 42784 4784 42852
rect 4708 42728 4718 42784
rect 4774 42728 4784 42784
rect 4708 42660 4784 42728
rect 4708 42604 4718 42660
rect 4774 42604 4784 42660
rect 4708 42536 4784 42604
rect 4708 42480 4718 42536
rect 4774 42480 4784 42536
rect 4708 42412 4784 42480
rect 4708 42356 4718 42412
rect 4774 42356 4784 42412
rect 4708 42288 4784 42356
rect 4708 42232 4718 42288
rect 4774 42232 4784 42288
rect 4708 42164 4784 42232
rect 4708 42108 4718 42164
rect 4774 42108 4784 42164
rect 4708 42098 4784 42108
rect 4832 43652 4908 43662
rect 5452 43653 5528 43663
rect 5576 45207 5652 45217
rect 5576 45151 5586 45207
rect 5642 45151 5652 45207
rect 5576 45083 5652 45151
rect 6384 45182 6460 45250
rect 6384 45126 6394 45182
rect 6450 45126 6460 45182
rect 5576 45027 5586 45083
rect 5642 45027 5652 45083
rect 5576 44959 5652 45027
rect 5576 44903 5586 44959
rect 5642 44903 5652 44959
rect 5576 44835 5652 44903
rect 5576 44779 5586 44835
rect 5642 44779 5652 44835
rect 5576 44711 5652 44779
rect 5576 44655 5586 44711
rect 5642 44655 5652 44711
rect 5576 44587 5652 44655
rect 5576 44531 5586 44587
rect 5642 44531 5652 44587
rect 5576 44463 5652 44531
rect 5576 44407 5586 44463
rect 5642 44407 5652 44463
rect 5576 44339 5652 44407
rect 5576 44283 5586 44339
rect 5642 44283 5652 44339
rect 5576 44215 5652 44283
rect 5576 44159 5586 44215
rect 5642 44159 5652 44215
rect 5576 44091 5652 44159
rect 5576 44035 5586 44091
rect 5642 44035 5652 44091
rect 5576 43967 5652 44035
rect 5576 43911 5586 43967
rect 5642 43911 5652 43967
rect 5576 43843 5652 43911
rect 5576 43787 5586 43843
rect 5642 43787 5652 43843
rect 5576 43719 5652 43787
rect 5576 43663 5586 43719
rect 5642 43663 5652 43719
rect 4832 43596 4842 43652
rect 4898 43596 4908 43652
rect 4832 43528 4908 43596
rect 5576 43595 5652 43663
rect 5576 43539 5586 43595
rect 5642 43539 5652 43595
rect 4832 43472 4842 43528
rect 4898 43472 4908 43528
rect 4832 43404 4908 43472
rect 4832 43348 4842 43404
rect 4898 43348 4908 43404
rect 4832 43280 4908 43348
rect 4832 43224 4842 43280
rect 4898 43224 4908 43280
rect 4832 43156 4908 43224
rect 4832 43100 4842 43156
rect 4898 43100 4908 43156
rect 4832 43032 4908 43100
rect 4832 42976 4842 43032
rect 4898 42976 4908 43032
rect 4832 42908 4908 42976
rect 4832 42852 4842 42908
rect 4898 42852 4908 42908
rect 4832 42784 4908 42852
rect 4832 42728 4842 42784
rect 4898 42728 4908 42784
rect 4832 42660 4908 42728
rect 4832 42604 4842 42660
rect 4898 42604 4908 42660
rect 4832 42536 4908 42604
rect 4832 42480 4842 42536
rect 4898 42480 4908 42536
rect 4832 42412 4908 42480
rect 4832 42356 4842 42412
rect 4898 42356 4908 42412
rect 4832 42288 4908 42356
rect 4832 42232 4842 42288
rect 4898 42232 4908 42288
rect 4832 42164 4908 42232
rect 4832 42108 4842 42164
rect 4898 42108 4908 42164
rect 4832 42040 4908 42108
rect 4832 41984 4842 42040
rect 4898 41984 4908 42040
rect 4832 41974 4908 41984
rect 4956 43528 5032 43538
rect 5576 43529 5652 43539
rect 5700 45083 5776 45093
rect 5700 45027 5710 45083
rect 5766 45027 5776 45083
rect 5700 44959 5776 45027
rect 6384 45058 6460 45126
rect 6384 45002 6394 45058
rect 6450 45002 6460 45058
rect 6384 44992 6460 45002
rect 6508 46546 6584 46556
rect 6508 46490 6518 46546
rect 6574 46490 6584 46546
rect 6508 46422 6584 46490
rect 6508 46366 6518 46422
rect 6574 46366 6584 46422
rect 6508 46298 6584 46366
rect 6508 46242 6518 46298
rect 6574 46242 6584 46298
rect 6508 46174 6584 46242
rect 6508 46118 6518 46174
rect 6574 46118 6584 46174
rect 6508 46050 6584 46118
rect 6508 45994 6518 46050
rect 6574 45994 6584 46050
rect 6508 45926 6584 45994
rect 6508 45870 6518 45926
rect 6574 45870 6584 45926
rect 6508 45802 6584 45870
rect 6508 45746 6518 45802
rect 6574 45746 6584 45802
rect 6508 45678 6584 45746
rect 6508 45622 6518 45678
rect 6574 45622 6584 45678
rect 6508 45554 6584 45622
rect 6508 45498 6518 45554
rect 6574 45498 6584 45554
rect 6508 45430 6584 45498
rect 6508 45374 6518 45430
rect 6574 45374 6584 45430
rect 6508 45306 6584 45374
rect 6508 45250 6518 45306
rect 6574 45250 6584 45306
rect 6508 45182 6584 45250
rect 6508 45126 6518 45182
rect 6574 45126 6584 45182
rect 6508 45058 6584 45126
rect 6508 45002 6518 45058
rect 6574 45002 6584 45058
rect 5700 44903 5710 44959
rect 5766 44903 5776 44959
rect 5700 44835 5776 44903
rect 5700 44779 5710 44835
rect 5766 44779 5776 44835
rect 5700 44711 5776 44779
rect 5700 44655 5710 44711
rect 5766 44655 5776 44711
rect 5700 44587 5776 44655
rect 5700 44531 5710 44587
rect 5766 44531 5776 44587
rect 5700 44463 5776 44531
rect 5700 44407 5710 44463
rect 5766 44407 5776 44463
rect 5700 44339 5776 44407
rect 5700 44283 5710 44339
rect 5766 44283 5776 44339
rect 5700 44215 5776 44283
rect 5700 44159 5710 44215
rect 5766 44159 5776 44215
rect 5700 44091 5776 44159
rect 5700 44035 5710 44091
rect 5766 44035 5776 44091
rect 5700 43967 5776 44035
rect 5700 43911 5710 43967
rect 5766 43911 5776 43967
rect 5700 43843 5776 43911
rect 5700 43787 5710 43843
rect 5766 43787 5776 43843
rect 5700 43719 5776 43787
rect 5700 43663 5710 43719
rect 5766 43663 5776 43719
rect 5700 43595 5776 43663
rect 5700 43539 5710 43595
rect 5766 43539 5776 43595
rect 4956 43472 4966 43528
rect 5022 43472 5032 43528
rect 4956 43404 5032 43472
rect 5700 43471 5776 43539
rect 5700 43415 5710 43471
rect 5766 43415 5776 43471
rect 4956 43348 4966 43404
rect 5022 43348 5032 43404
rect 4956 43280 5032 43348
rect 4956 43224 4966 43280
rect 5022 43224 5032 43280
rect 4956 43156 5032 43224
rect 4956 43100 4966 43156
rect 5022 43100 5032 43156
rect 4956 43032 5032 43100
rect 4956 42976 4966 43032
rect 5022 42976 5032 43032
rect 4956 42908 5032 42976
rect 4956 42852 4966 42908
rect 5022 42852 5032 42908
rect 4956 42784 5032 42852
rect 4956 42728 4966 42784
rect 5022 42728 5032 42784
rect 4956 42660 5032 42728
rect 4956 42604 4966 42660
rect 5022 42604 5032 42660
rect 4956 42536 5032 42604
rect 4956 42480 4966 42536
rect 5022 42480 5032 42536
rect 4956 42412 5032 42480
rect 4956 42356 4966 42412
rect 5022 42356 5032 42412
rect 4956 42288 5032 42356
rect 4956 42232 4966 42288
rect 5022 42232 5032 42288
rect 4956 42164 5032 42232
rect 4956 42108 4966 42164
rect 5022 42108 5032 42164
rect 4956 42040 5032 42108
rect 4956 41984 4966 42040
rect 5022 41984 5032 42040
rect 4956 41916 5032 41984
rect 4956 41860 4966 41916
rect 5022 41860 5032 41916
rect 4956 41850 5032 41860
rect 5080 43404 5156 43414
rect 5700 43405 5776 43415
rect 5824 44959 5900 44969
rect 5824 44903 5834 44959
rect 5890 44903 5900 44959
rect 5824 44835 5900 44903
rect 6508 44934 6584 45002
rect 6508 44878 6518 44934
rect 6574 44878 6584 44934
rect 6508 44868 6584 44878
rect 6632 46422 6708 46432
rect 6632 46366 6642 46422
rect 6698 46366 6708 46422
rect 6632 46298 6708 46366
rect 6632 46242 6642 46298
rect 6698 46242 6708 46298
rect 6632 46174 6708 46242
rect 6632 46118 6642 46174
rect 6698 46118 6708 46174
rect 6632 46050 6708 46118
rect 6632 45994 6642 46050
rect 6698 45994 6708 46050
rect 6632 45926 6708 45994
rect 6632 45870 6642 45926
rect 6698 45870 6708 45926
rect 6632 45802 6708 45870
rect 6632 45746 6642 45802
rect 6698 45746 6708 45802
rect 6632 45678 6708 45746
rect 6632 45622 6642 45678
rect 6698 45622 6708 45678
rect 6632 45554 6708 45622
rect 6632 45498 6642 45554
rect 6698 45498 6708 45554
rect 6632 45430 6708 45498
rect 6632 45374 6642 45430
rect 6698 45374 6708 45430
rect 6632 45306 6708 45374
rect 6632 45250 6642 45306
rect 6698 45250 6708 45306
rect 6632 45182 6708 45250
rect 6632 45126 6642 45182
rect 6698 45126 6708 45182
rect 6632 45058 6708 45126
rect 6632 45002 6642 45058
rect 6698 45002 6708 45058
rect 6632 44934 6708 45002
rect 6632 44878 6642 44934
rect 6698 44878 6708 44934
rect 5824 44779 5834 44835
rect 5890 44779 5900 44835
rect 5824 44711 5900 44779
rect 5824 44655 5834 44711
rect 5890 44655 5900 44711
rect 5824 44587 5900 44655
rect 5824 44531 5834 44587
rect 5890 44531 5900 44587
rect 5824 44463 5900 44531
rect 5824 44407 5834 44463
rect 5890 44407 5900 44463
rect 5824 44339 5900 44407
rect 5824 44283 5834 44339
rect 5890 44283 5900 44339
rect 5824 44215 5900 44283
rect 5824 44159 5834 44215
rect 5890 44159 5900 44215
rect 5824 44091 5900 44159
rect 5824 44035 5834 44091
rect 5890 44035 5900 44091
rect 5824 43967 5900 44035
rect 5824 43911 5834 43967
rect 5890 43911 5900 43967
rect 5824 43843 5900 43911
rect 5824 43787 5834 43843
rect 5890 43787 5900 43843
rect 5824 43719 5900 43787
rect 5824 43663 5834 43719
rect 5890 43663 5900 43719
rect 5824 43595 5900 43663
rect 5824 43539 5834 43595
rect 5890 43539 5900 43595
rect 5824 43471 5900 43539
rect 5824 43415 5834 43471
rect 5890 43415 5900 43471
rect 5080 43348 5090 43404
rect 5146 43348 5156 43404
rect 5080 43280 5156 43348
rect 5824 43347 5900 43415
rect 5824 43291 5834 43347
rect 5890 43291 5900 43347
rect 5080 43224 5090 43280
rect 5146 43224 5156 43280
rect 5080 43156 5156 43224
rect 5080 43100 5090 43156
rect 5146 43100 5156 43156
rect 5080 43032 5156 43100
rect 5080 42976 5090 43032
rect 5146 42976 5156 43032
rect 5080 42908 5156 42976
rect 5080 42852 5090 42908
rect 5146 42852 5156 42908
rect 5080 42784 5156 42852
rect 5080 42728 5090 42784
rect 5146 42728 5156 42784
rect 5080 42660 5156 42728
rect 5080 42604 5090 42660
rect 5146 42604 5156 42660
rect 5080 42536 5156 42604
rect 5080 42480 5090 42536
rect 5146 42480 5156 42536
rect 5080 42412 5156 42480
rect 5080 42356 5090 42412
rect 5146 42356 5156 42412
rect 5080 42288 5156 42356
rect 5080 42232 5090 42288
rect 5146 42232 5156 42288
rect 5080 42164 5156 42232
rect 5080 42108 5090 42164
rect 5146 42108 5156 42164
rect 5080 42040 5156 42108
rect 5080 41984 5090 42040
rect 5146 41984 5156 42040
rect 5080 41916 5156 41984
rect 5080 41860 5090 41916
rect 5146 41860 5156 41916
rect 4460 41789 4536 41799
rect 4460 41733 4470 41789
rect 4526 41733 4536 41789
rect 4460 41665 4536 41733
rect 5080 41792 5156 41860
rect 5080 41736 5090 41792
rect 5146 41736 5156 41792
rect 5080 41726 5156 41736
rect 5204 43280 5280 43290
rect 5824 43281 5900 43291
rect 5948 44835 6024 44845
rect 5948 44779 5958 44835
rect 6014 44779 6024 44835
rect 5948 44711 6024 44779
rect 6632 44810 6708 44878
rect 6632 44754 6642 44810
rect 6698 44754 6708 44810
rect 6632 44744 6708 44754
rect 6756 46298 6832 46308
rect 6756 46242 6766 46298
rect 6822 46242 6832 46298
rect 6756 46174 6832 46242
rect 6756 46118 6766 46174
rect 6822 46118 6832 46174
rect 6756 46050 6832 46118
rect 6756 45994 6766 46050
rect 6822 45994 6832 46050
rect 6756 45926 6832 45994
rect 6756 45870 6766 45926
rect 6822 45870 6832 45926
rect 6756 45802 6832 45870
rect 6756 45746 6766 45802
rect 6822 45746 6832 45802
rect 6756 45678 6832 45746
rect 6756 45622 6766 45678
rect 6822 45622 6832 45678
rect 6756 45554 6832 45622
rect 6756 45498 6766 45554
rect 6822 45498 6832 45554
rect 6756 45430 6832 45498
rect 6756 45374 6766 45430
rect 6822 45374 6832 45430
rect 6756 45306 6832 45374
rect 6756 45250 6766 45306
rect 6822 45250 6832 45306
rect 6756 45182 6832 45250
rect 6756 45126 6766 45182
rect 6822 45126 6832 45182
rect 6756 45058 6832 45126
rect 6756 45002 6766 45058
rect 6822 45002 6832 45058
rect 6756 44934 6832 45002
rect 6756 44878 6766 44934
rect 6822 44878 6832 44934
rect 6756 44810 6832 44878
rect 6756 44754 6766 44810
rect 6822 44754 6832 44810
rect 5948 44655 5958 44711
rect 6014 44655 6024 44711
rect 5948 44587 6024 44655
rect 5948 44531 5958 44587
rect 6014 44531 6024 44587
rect 5948 44463 6024 44531
rect 5948 44407 5958 44463
rect 6014 44407 6024 44463
rect 5948 44339 6024 44407
rect 5948 44283 5958 44339
rect 6014 44283 6024 44339
rect 5948 44215 6024 44283
rect 5948 44159 5958 44215
rect 6014 44159 6024 44215
rect 5948 44091 6024 44159
rect 5948 44035 5958 44091
rect 6014 44035 6024 44091
rect 5948 43967 6024 44035
rect 5948 43911 5958 43967
rect 6014 43911 6024 43967
rect 5948 43843 6024 43911
rect 5948 43787 5958 43843
rect 6014 43787 6024 43843
rect 5948 43719 6024 43787
rect 5948 43663 5958 43719
rect 6014 43663 6024 43719
rect 5948 43595 6024 43663
rect 5948 43539 5958 43595
rect 6014 43539 6024 43595
rect 5948 43471 6024 43539
rect 5948 43415 5958 43471
rect 6014 43415 6024 43471
rect 5948 43347 6024 43415
rect 5948 43291 5958 43347
rect 6014 43291 6024 43347
rect 5204 43224 5214 43280
rect 5270 43224 5280 43280
rect 5204 43156 5280 43224
rect 5948 43223 6024 43291
rect 5948 43167 5958 43223
rect 6014 43167 6024 43223
rect 5204 43100 5214 43156
rect 5270 43100 5280 43156
rect 5204 43032 5280 43100
rect 5204 42976 5214 43032
rect 5270 42976 5280 43032
rect 5204 42908 5280 42976
rect 5204 42852 5214 42908
rect 5270 42852 5280 42908
rect 5204 42784 5280 42852
rect 5204 42728 5214 42784
rect 5270 42728 5280 42784
rect 5204 42660 5280 42728
rect 5204 42604 5214 42660
rect 5270 42604 5280 42660
rect 5204 42536 5280 42604
rect 5204 42480 5214 42536
rect 5270 42480 5280 42536
rect 5204 42412 5280 42480
rect 5204 42356 5214 42412
rect 5270 42356 5280 42412
rect 5204 42288 5280 42356
rect 5204 42232 5214 42288
rect 5270 42232 5280 42288
rect 5204 42164 5280 42232
rect 5204 42108 5214 42164
rect 5270 42108 5280 42164
rect 5204 42040 5280 42108
rect 5204 41984 5214 42040
rect 5270 41984 5280 42040
rect 5204 41916 5280 41984
rect 5204 41860 5214 41916
rect 5270 41860 5280 41916
rect 5204 41792 5280 41860
rect 5204 41736 5214 41792
rect 5270 41736 5280 41792
rect 4460 41609 4470 41665
rect 4526 41609 4536 41665
rect 4460 41541 4536 41609
rect 4460 41485 4470 41541
rect 4526 41485 4536 41541
rect 4460 41417 4536 41485
rect 4460 41361 4470 41417
rect 4526 41361 4536 41417
rect 4460 41293 4536 41361
rect 4460 41237 4470 41293
rect 4526 41237 4536 41293
rect 4460 41169 4536 41237
rect 4460 41113 4470 41169
rect 4526 41113 4536 41169
rect 4460 41045 4536 41113
rect 4460 40989 4470 41045
rect 4526 40989 4536 41045
rect 4460 40921 4536 40989
rect 4460 40865 4470 40921
rect 4526 40865 4536 40921
rect 4460 40797 4536 40865
rect 4460 40741 4470 40797
rect 4526 40741 4536 40797
rect 4460 40673 4536 40741
rect 4460 40617 4470 40673
rect 4526 40617 4536 40673
rect 4460 40549 4536 40617
rect 4460 40493 4470 40549
rect 4526 40493 4536 40549
rect 4460 40425 4536 40493
rect 4460 40369 4470 40425
rect 4526 40369 4536 40425
rect 4460 40301 4536 40369
rect 4460 40245 4470 40301
rect 4526 40245 4536 40301
rect 4460 40177 4536 40245
rect 4460 40121 4470 40177
rect 4526 40121 4536 40177
rect 4460 40111 4536 40121
rect 4584 41665 4660 41675
rect 4584 41609 4594 41665
rect 4650 41609 4660 41665
rect 4584 41541 4660 41609
rect 5204 41668 5280 41736
rect 5204 41612 5214 41668
rect 5270 41612 5280 41668
rect 5204 41602 5280 41612
rect 5328 43156 5404 43166
rect 5948 43157 6024 43167
rect 6072 44711 6148 44721
rect 6072 44655 6082 44711
rect 6138 44655 6148 44711
rect 6072 44587 6148 44655
rect 6756 44686 6832 44754
rect 6756 44630 6766 44686
rect 6822 44630 6832 44686
rect 6756 44620 6832 44630
rect 6880 46174 6956 46184
rect 6880 46118 6890 46174
rect 6946 46118 6956 46174
rect 6880 46050 6956 46118
rect 6880 45994 6890 46050
rect 6946 45994 6956 46050
rect 6880 45926 6956 45994
rect 6880 45870 6890 45926
rect 6946 45870 6956 45926
rect 6880 45802 6956 45870
rect 6880 45746 6890 45802
rect 6946 45746 6956 45802
rect 6880 45678 6956 45746
rect 6880 45622 6890 45678
rect 6946 45622 6956 45678
rect 6880 45554 6956 45622
rect 6880 45498 6890 45554
rect 6946 45498 6956 45554
rect 6880 45430 6956 45498
rect 6880 45374 6890 45430
rect 6946 45374 6956 45430
rect 6880 45306 6956 45374
rect 6880 45250 6890 45306
rect 6946 45250 6956 45306
rect 6880 45182 6956 45250
rect 6880 45126 6890 45182
rect 6946 45126 6956 45182
rect 6880 45058 6956 45126
rect 6880 45002 6890 45058
rect 6946 45002 6956 45058
rect 6880 44934 6956 45002
rect 6880 44878 6890 44934
rect 6946 44878 6956 44934
rect 6880 44810 6956 44878
rect 6880 44754 6890 44810
rect 6946 44754 6956 44810
rect 6880 44686 6956 44754
rect 6880 44630 6890 44686
rect 6946 44630 6956 44686
rect 6072 44531 6082 44587
rect 6138 44531 6148 44587
rect 6072 44463 6148 44531
rect 6880 44562 6956 44630
rect 6880 44506 6890 44562
rect 6946 44506 6956 44562
rect 6880 44496 6956 44506
rect 7004 46050 7080 46060
rect 7004 45994 7014 46050
rect 7070 45994 7080 46050
rect 7004 45926 7080 45994
rect 7004 45870 7014 45926
rect 7070 45870 7080 45926
rect 7004 45802 7080 45870
rect 7004 45746 7014 45802
rect 7070 45746 7080 45802
rect 7004 45678 7080 45746
rect 7004 45622 7014 45678
rect 7070 45622 7080 45678
rect 7004 45554 7080 45622
rect 7004 45498 7014 45554
rect 7070 45498 7080 45554
rect 7004 45430 7080 45498
rect 7004 45374 7014 45430
rect 7070 45374 7080 45430
rect 7004 45306 7080 45374
rect 7004 45250 7014 45306
rect 7070 45250 7080 45306
rect 7004 45182 7080 45250
rect 7004 45126 7014 45182
rect 7070 45126 7080 45182
rect 7004 45058 7080 45126
rect 7004 45002 7014 45058
rect 7070 45002 7080 45058
rect 7004 44934 7080 45002
rect 7004 44878 7014 44934
rect 7070 44878 7080 44934
rect 7004 44810 7080 44878
rect 7004 44754 7014 44810
rect 7070 44754 7080 44810
rect 7004 44686 7080 44754
rect 7004 44630 7014 44686
rect 7070 44630 7080 44686
rect 7004 44562 7080 44630
rect 7004 44506 7014 44562
rect 7070 44506 7080 44562
rect 6072 44407 6082 44463
rect 6138 44407 6148 44463
rect 6072 44339 6148 44407
rect 7004 44438 7080 44506
rect 7004 44382 7014 44438
rect 7070 44382 7080 44438
rect 7004 44372 7080 44382
rect 7128 45926 7204 45936
rect 7128 45870 7138 45926
rect 7194 45870 7204 45926
rect 7128 45802 7204 45870
rect 7128 45746 7138 45802
rect 7194 45746 7204 45802
rect 7128 45678 7204 45746
rect 7128 45622 7138 45678
rect 7194 45622 7204 45678
rect 7128 45554 7204 45622
rect 7128 45498 7138 45554
rect 7194 45498 7204 45554
rect 7128 45430 7204 45498
rect 7128 45374 7138 45430
rect 7194 45374 7204 45430
rect 7128 45306 7204 45374
rect 7128 45250 7138 45306
rect 7194 45250 7204 45306
rect 7128 45182 7204 45250
rect 7128 45126 7138 45182
rect 7194 45126 7204 45182
rect 7128 45058 7204 45126
rect 7128 45002 7138 45058
rect 7194 45002 7204 45058
rect 7128 44934 7204 45002
rect 7128 44878 7138 44934
rect 7194 44878 7204 44934
rect 7128 44810 7204 44878
rect 7128 44754 7138 44810
rect 7194 44754 7204 44810
rect 7128 44686 7204 44754
rect 7128 44630 7138 44686
rect 7194 44630 7204 44686
rect 7128 44562 7204 44630
rect 7128 44506 7138 44562
rect 7194 44506 7204 44562
rect 7128 44438 7204 44506
rect 7128 44382 7138 44438
rect 7194 44382 7204 44438
rect 6072 44283 6082 44339
rect 6138 44283 6148 44339
rect 6072 44215 6148 44283
rect 7128 44314 7204 44382
rect 7128 44258 7138 44314
rect 7194 44258 7204 44314
rect 7128 44248 7204 44258
rect 7252 45802 7328 45812
rect 7252 45746 7262 45802
rect 7318 45746 7328 45802
rect 7252 45678 7328 45746
rect 7252 45622 7262 45678
rect 7318 45622 7328 45678
rect 7252 45554 7328 45622
rect 7252 45498 7262 45554
rect 7318 45498 7328 45554
rect 7252 45430 7328 45498
rect 7252 45374 7262 45430
rect 7318 45374 7328 45430
rect 7252 45306 7328 45374
rect 7252 45250 7262 45306
rect 7318 45250 7328 45306
rect 7252 45182 7328 45250
rect 7252 45126 7262 45182
rect 7318 45126 7328 45182
rect 7252 45058 7328 45126
rect 7252 45002 7262 45058
rect 7318 45002 7328 45058
rect 7252 44934 7328 45002
rect 7252 44878 7262 44934
rect 7318 44878 7328 44934
rect 7252 44810 7328 44878
rect 7252 44754 7262 44810
rect 7318 44754 7328 44810
rect 7252 44686 7328 44754
rect 7252 44630 7262 44686
rect 7318 44630 7328 44686
rect 7252 44562 7328 44630
rect 7252 44506 7262 44562
rect 7318 44506 7328 44562
rect 7252 44438 7328 44506
rect 7252 44382 7262 44438
rect 7318 44382 7328 44438
rect 7252 44314 7328 44382
rect 7252 44258 7262 44314
rect 7318 44258 7328 44314
rect 6072 44159 6082 44215
rect 6138 44159 6148 44215
rect 6072 44091 6148 44159
rect 7252 44190 7328 44258
rect 7252 44134 7262 44190
rect 7318 44134 7328 44190
rect 7252 44124 7328 44134
rect 8741 44544 10553 44554
rect 8741 44488 8751 44544
rect 8807 44488 8875 44544
rect 8931 44488 8999 44544
rect 9055 44488 9123 44544
rect 9179 44488 9247 44544
rect 9303 44488 9371 44544
rect 9427 44488 9495 44544
rect 9551 44488 9619 44544
rect 9675 44488 9743 44544
rect 9799 44488 9867 44544
rect 9923 44488 9991 44544
rect 10047 44488 10115 44544
rect 10171 44488 10239 44544
rect 10295 44488 10363 44544
rect 10419 44488 10487 44544
rect 10543 44488 10553 44544
rect 8741 44420 10553 44488
rect 8741 44364 8751 44420
rect 8807 44364 8875 44420
rect 8931 44364 8999 44420
rect 9055 44364 9123 44420
rect 9179 44364 9247 44420
rect 9303 44364 9371 44420
rect 9427 44364 9495 44420
rect 9551 44364 9619 44420
rect 9675 44364 9743 44420
rect 9799 44364 9867 44420
rect 9923 44364 9991 44420
rect 10047 44364 10115 44420
rect 10171 44364 10239 44420
rect 10295 44364 10363 44420
rect 10419 44364 10487 44420
rect 10543 44364 10553 44420
rect 8741 44296 10553 44364
rect 8741 44240 8751 44296
rect 8807 44240 8875 44296
rect 8931 44240 8999 44296
rect 9055 44240 9123 44296
rect 9179 44240 9247 44296
rect 9303 44240 9371 44296
rect 9427 44240 9495 44296
rect 9551 44240 9619 44296
rect 9675 44240 9743 44296
rect 9799 44240 9867 44296
rect 9923 44240 9991 44296
rect 10047 44240 10115 44296
rect 10171 44240 10239 44296
rect 10295 44240 10363 44296
rect 10419 44240 10487 44296
rect 10543 44240 10553 44296
rect 8741 44172 10553 44240
rect 6072 44035 6082 44091
rect 6138 44035 6148 44091
rect 6072 43967 6148 44035
rect 6072 43911 6082 43967
rect 6138 43911 6148 43967
rect 6072 43843 6148 43911
rect 6072 43787 6082 43843
rect 6138 43787 6148 43843
rect 6072 43719 6148 43787
rect 6072 43663 6082 43719
rect 6138 43663 6148 43719
rect 6072 43595 6148 43663
rect 6072 43539 6082 43595
rect 6138 43539 6148 43595
rect 6072 43471 6148 43539
rect 6072 43415 6082 43471
rect 6138 43415 6148 43471
rect 6072 43347 6148 43415
rect 6072 43291 6082 43347
rect 6138 43291 6148 43347
rect 6072 43223 6148 43291
rect 8741 44116 8751 44172
rect 8807 44116 8875 44172
rect 8931 44116 8999 44172
rect 9055 44116 9123 44172
rect 9179 44116 9247 44172
rect 9303 44116 9371 44172
rect 9427 44116 9495 44172
rect 9551 44116 9619 44172
rect 9675 44116 9743 44172
rect 9799 44116 9867 44172
rect 9923 44116 9991 44172
rect 10047 44116 10115 44172
rect 10171 44116 10239 44172
rect 10295 44116 10363 44172
rect 10419 44116 10487 44172
rect 10543 44116 10553 44172
rect 8741 44048 10553 44116
rect 8741 43992 8751 44048
rect 8807 43992 8875 44048
rect 8931 43992 8999 44048
rect 9055 43992 9123 44048
rect 9179 43992 9247 44048
rect 9303 43992 9371 44048
rect 9427 43992 9495 44048
rect 9551 43992 9619 44048
rect 9675 43992 9743 44048
rect 9799 43992 9867 44048
rect 9923 43992 9991 44048
rect 10047 43992 10115 44048
rect 10171 43992 10239 44048
rect 10295 43992 10363 44048
rect 10419 43992 10487 44048
rect 10543 43992 10553 44048
rect 8741 43924 10553 43992
rect 8741 43868 8751 43924
rect 8807 43868 8875 43924
rect 8931 43868 8999 43924
rect 9055 43868 9123 43924
rect 9179 43868 9247 43924
rect 9303 43868 9371 43924
rect 9427 43868 9495 43924
rect 9551 43868 9619 43924
rect 9675 43868 9743 43924
rect 9799 43868 9867 43924
rect 9923 43868 9991 43924
rect 10047 43868 10115 43924
rect 10171 43868 10239 43924
rect 10295 43868 10363 43924
rect 10419 43868 10487 43924
rect 10543 43868 10553 43924
rect 8741 43800 10553 43868
rect 8741 43744 8751 43800
rect 8807 43744 8875 43800
rect 8931 43744 8999 43800
rect 9055 43744 9123 43800
rect 9179 43744 9247 43800
rect 9303 43744 9371 43800
rect 9427 43744 9495 43800
rect 9551 43744 9619 43800
rect 9675 43744 9743 43800
rect 9799 43744 9867 43800
rect 9923 43744 9991 43800
rect 10047 43744 10115 43800
rect 10171 43744 10239 43800
rect 10295 43744 10363 43800
rect 10419 43744 10487 43800
rect 10543 43744 10553 43800
rect 8741 43676 10553 43744
rect 8741 43620 8751 43676
rect 8807 43620 8875 43676
rect 8931 43620 8999 43676
rect 9055 43620 9123 43676
rect 9179 43620 9247 43676
rect 9303 43620 9371 43676
rect 9427 43620 9495 43676
rect 9551 43620 9619 43676
rect 9675 43620 9743 43676
rect 9799 43620 9867 43676
rect 9923 43620 9991 43676
rect 10047 43620 10115 43676
rect 10171 43620 10239 43676
rect 10295 43620 10363 43676
rect 10419 43620 10487 43676
rect 10543 43620 10553 43676
rect 8741 43552 10553 43620
rect 8741 43496 8751 43552
rect 8807 43496 8875 43552
rect 8931 43496 8999 43552
rect 9055 43496 9123 43552
rect 9179 43496 9247 43552
rect 9303 43496 9371 43552
rect 9427 43496 9495 43552
rect 9551 43496 9619 43552
rect 9675 43496 9743 43552
rect 9799 43496 9867 43552
rect 9923 43496 9991 43552
rect 10047 43496 10115 43552
rect 10171 43496 10239 43552
rect 10295 43496 10363 43552
rect 10419 43496 10487 43552
rect 10543 43496 10553 43552
rect 8741 43428 10553 43496
rect 8741 43372 8751 43428
rect 8807 43372 8875 43428
rect 8931 43372 8999 43428
rect 9055 43372 9123 43428
rect 9179 43372 9247 43428
rect 9303 43372 9371 43428
rect 9427 43372 9495 43428
rect 9551 43372 9619 43428
rect 9675 43372 9743 43428
rect 9799 43372 9867 43428
rect 9923 43372 9991 43428
rect 10047 43372 10115 43428
rect 10171 43372 10239 43428
rect 10295 43372 10363 43428
rect 10419 43372 10487 43428
rect 10543 43372 10553 43428
rect 8741 43304 10553 43372
rect 8741 43248 8751 43304
rect 8807 43248 8875 43304
rect 8931 43248 8999 43304
rect 9055 43248 9123 43304
rect 9179 43248 9247 43304
rect 9303 43248 9371 43304
rect 9427 43248 9495 43304
rect 9551 43248 9619 43304
rect 9675 43248 9743 43304
rect 9799 43248 9867 43304
rect 9923 43248 9991 43304
rect 10047 43248 10115 43304
rect 10171 43248 10239 43304
rect 10295 43248 10363 43304
rect 10419 43248 10487 43304
rect 10543 43248 10553 43304
rect 8741 43238 10553 43248
rect 12842 44544 13910 44554
rect 12842 44488 12852 44544
rect 12908 44488 12976 44544
rect 13032 44488 13100 44544
rect 13156 44488 13224 44544
rect 13280 44488 13348 44544
rect 13404 44488 13472 44544
rect 13528 44488 13596 44544
rect 13652 44488 13720 44544
rect 13776 44488 13844 44544
rect 13900 44488 13910 44544
rect 12842 44420 13910 44488
rect 12842 44364 12852 44420
rect 12908 44364 12976 44420
rect 13032 44364 13100 44420
rect 13156 44364 13224 44420
rect 13280 44364 13348 44420
rect 13404 44364 13472 44420
rect 13528 44364 13596 44420
rect 13652 44364 13720 44420
rect 13776 44364 13844 44420
rect 13900 44364 13910 44420
rect 12842 44296 13910 44364
rect 12842 44240 12852 44296
rect 12908 44240 12976 44296
rect 13032 44240 13100 44296
rect 13156 44240 13224 44296
rect 13280 44240 13348 44296
rect 13404 44240 13472 44296
rect 13528 44240 13596 44296
rect 13652 44240 13720 44296
rect 13776 44240 13844 44296
rect 13900 44240 13910 44296
rect 12842 44172 13910 44240
rect 12842 44116 12852 44172
rect 12908 44116 12976 44172
rect 13032 44116 13100 44172
rect 13156 44116 13224 44172
rect 13280 44116 13348 44172
rect 13404 44116 13472 44172
rect 13528 44116 13596 44172
rect 13652 44116 13720 44172
rect 13776 44116 13844 44172
rect 13900 44116 13910 44172
rect 12842 44048 13910 44116
rect 12842 43992 12852 44048
rect 12908 43992 12976 44048
rect 13032 43992 13100 44048
rect 13156 43992 13224 44048
rect 13280 43992 13348 44048
rect 13404 43992 13472 44048
rect 13528 43992 13596 44048
rect 13652 43992 13720 44048
rect 13776 43992 13844 44048
rect 13900 43992 13910 44048
rect 12842 43924 13910 43992
rect 12842 43868 12852 43924
rect 12908 43868 12976 43924
rect 13032 43868 13100 43924
rect 13156 43868 13224 43924
rect 13280 43868 13348 43924
rect 13404 43868 13472 43924
rect 13528 43868 13596 43924
rect 13652 43868 13720 43924
rect 13776 43868 13844 43924
rect 13900 43868 13910 43924
rect 12842 43800 13910 43868
rect 12842 43744 12852 43800
rect 12908 43744 12976 43800
rect 13032 43744 13100 43800
rect 13156 43744 13224 43800
rect 13280 43744 13348 43800
rect 13404 43744 13472 43800
rect 13528 43744 13596 43800
rect 13652 43744 13720 43800
rect 13776 43744 13844 43800
rect 13900 43744 13910 43800
rect 12842 43676 13910 43744
rect 12842 43620 12852 43676
rect 12908 43620 12976 43676
rect 13032 43620 13100 43676
rect 13156 43620 13224 43676
rect 13280 43620 13348 43676
rect 13404 43620 13472 43676
rect 13528 43620 13596 43676
rect 13652 43620 13720 43676
rect 13776 43620 13844 43676
rect 13900 43620 13910 43676
rect 12842 43552 13910 43620
rect 12842 43496 12852 43552
rect 12908 43496 12976 43552
rect 13032 43496 13100 43552
rect 13156 43496 13224 43552
rect 13280 43496 13348 43552
rect 13404 43496 13472 43552
rect 13528 43496 13596 43552
rect 13652 43496 13720 43552
rect 13776 43496 13844 43552
rect 13900 43496 13910 43552
rect 12842 43428 13910 43496
rect 12842 43372 12852 43428
rect 12908 43372 12976 43428
rect 13032 43372 13100 43428
rect 13156 43372 13224 43428
rect 13280 43372 13348 43428
rect 13404 43372 13472 43428
rect 13528 43372 13596 43428
rect 13652 43372 13720 43428
rect 13776 43372 13844 43428
rect 13900 43372 13910 43428
rect 12842 43304 13910 43372
rect 12842 43248 12852 43304
rect 12908 43248 12976 43304
rect 13032 43248 13100 43304
rect 13156 43248 13224 43304
rect 13280 43248 13348 43304
rect 13404 43248 13472 43304
rect 13528 43248 13596 43304
rect 13652 43248 13720 43304
rect 13776 43248 13844 43304
rect 13900 43248 13910 43304
rect 12842 43238 13910 43248
rect 6072 43167 6082 43223
rect 6138 43167 6148 43223
rect 5328 43100 5338 43156
rect 5394 43100 5404 43156
rect 5328 43032 5404 43100
rect 6072 43099 6148 43167
rect 6072 43043 6082 43099
rect 6138 43043 6148 43099
rect 5328 42976 5338 43032
rect 5394 42976 5404 43032
rect 5328 42908 5404 42976
rect 5328 42852 5338 42908
rect 5394 42852 5404 42908
rect 5328 42784 5404 42852
rect 5328 42728 5338 42784
rect 5394 42728 5404 42784
rect 5328 42660 5404 42728
rect 5328 42604 5338 42660
rect 5394 42604 5404 42660
rect 5328 42536 5404 42604
rect 5328 42480 5338 42536
rect 5394 42480 5404 42536
rect 5328 42412 5404 42480
rect 5328 42356 5338 42412
rect 5394 42356 5404 42412
rect 5328 42288 5404 42356
rect 5328 42232 5338 42288
rect 5394 42232 5404 42288
rect 5328 42164 5404 42232
rect 5328 42108 5338 42164
rect 5394 42108 5404 42164
rect 5328 42040 5404 42108
rect 5328 41984 5338 42040
rect 5394 41984 5404 42040
rect 5328 41916 5404 41984
rect 5328 41860 5338 41916
rect 5394 41860 5404 41916
rect 5328 41792 5404 41860
rect 5328 41736 5338 41792
rect 5394 41736 5404 41792
rect 5328 41668 5404 41736
rect 5328 41612 5338 41668
rect 5394 41612 5404 41668
rect 4584 41485 4594 41541
rect 4650 41485 4660 41541
rect 4584 41417 4660 41485
rect 4584 41361 4594 41417
rect 4650 41361 4660 41417
rect 4584 41293 4660 41361
rect 4584 41237 4594 41293
rect 4650 41237 4660 41293
rect 4584 41169 4660 41237
rect 4584 41113 4594 41169
rect 4650 41113 4660 41169
rect 4584 41045 4660 41113
rect 4584 40989 4594 41045
rect 4650 40989 4660 41045
rect 4584 40921 4660 40989
rect 4584 40865 4594 40921
rect 4650 40865 4660 40921
rect 4584 40797 4660 40865
rect 4584 40741 4594 40797
rect 4650 40741 4660 40797
rect 4584 40673 4660 40741
rect 4584 40617 4594 40673
rect 4650 40617 4660 40673
rect 4584 40549 4660 40617
rect 4584 40493 4594 40549
rect 4650 40493 4660 40549
rect 4584 40425 4660 40493
rect 4584 40369 4594 40425
rect 4650 40369 4660 40425
rect 4584 40301 4660 40369
rect 4584 40245 4594 40301
rect 4650 40245 4660 40301
rect 4584 40177 4660 40245
rect 4584 40121 4594 40177
rect 4650 40121 4660 40177
rect 4584 40053 4660 40121
rect 4584 39997 4594 40053
rect 4650 39997 4660 40053
rect 4584 39987 4660 39997
rect 4708 41541 4784 41551
rect 4708 41485 4718 41541
rect 4774 41485 4784 41541
rect 4708 41417 4784 41485
rect 5328 41544 5404 41612
rect 5328 41488 5338 41544
rect 5394 41488 5404 41544
rect 5328 41478 5404 41488
rect 5452 43032 5528 43042
rect 6072 43033 6148 43043
rect 5452 42976 5462 43032
rect 5518 42976 5528 43032
rect 5452 42908 5528 42976
rect 7552 42944 8620 42954
rect 5452 42852 5462 42908
rect 5518 42852 5528 42908
rect 5452 42784 5528 42852
rect 5452 42728 5462 42784
rect 5518 42728 5528 42784
rect 5452 42660 5528 42728
rect 5452 42604 5462 42660
rect 5518 42604 5528 42660
rect 5452 42536 5528 42604
rect 5452 42480 5462 42536
rect 5518 42480 5528 42536
rect 5452 42412 5528 42480
rect 5452 42356 5462 42412
rect 5518 42356 5528 42412
rect 5452 42288 5528 42356
rect 5452 42232 5462 42288
rect 5518 42232 5528 42288
rect 5452 42164 5528 42232
rect 5452 42108 5462 42164
rect 5518 42108 5528 42164
rect 5452 42040 5528 42108
rect 5452 41984 5462 42040
rect 5518 41984 5528 42040
rect 5452 41916 5528 41984
rect 5452 41860 5462 41916
rect 5518 41860 5528 41916
rect 5452 41792 5528 41860
rect 5452 41736 5462 41792
rect 5518 41736 5528 41792
rect 5452 41668 5528 41736
rect 5452 41612 5462 41668
rect 5518 41612 5528 41668
rect 5452 41544 5528 41612
rect 5452 41488 5462 41544
rect 5518 41488 5528 41544
rect 4708 41361 4718 41417
rect 4774 41361 4784 41417
rect 4708 41293 4784 41361
rect 4708 41237 4718 41293
rect 4774 41237 4784 41293
rect 4708 41169 4784 41237
rect 4708 41113 4718 41169
rect 4774 41113 4784 41169
rect 4708 41045 4784 41113
rect 4708 40989 4718 41045
rect 4774 40989 4784 41045
rect 4708 40921 4784 40989
rect 4708 40865 4718 40921
rect 4774 40865 4784 40921
rect 4708 40797 4784 40865
rect 4708 40741 4718 40797
rect 4774 40741 4784 40797
rect 4708 40673 4784 40741
rect 4708 40617 4718 40673
rect 4774 40617 4784 40673
rect 4708 40549 4784 40617
rect 4708 40493 4718 40549
rect 4774 40493 4784 40549
rect 4708 40425 4784 40493
rect 4708 40369 4718 40425
rect 4774 40369 4784 40425
rect 4708 40301 4784 40369
rect 4708 40245 4718 40301
rect 4774 40245 4784 40301
rect 4708 40177 4784 40245
rect 4708 40121 4718 40177
rect 4774 40121 4784 40177
rect 4708 40053 4784 40121
rect 4708 39997 4718 40053
rect 4774 39997 4784 40053
rect 4708 39929 4784 39997
rect 4708 39873 4718 39929
rect 4774 39873 4784 39929
rect 4708 39863 4784 39873
rect 4832 41417 4908 41427
rect 4832 41361 4842 41417
rect 4898 41361 4908 41417
rect 4832 41293 4908 41361
rect 5452 41420 5528 41488
rect 5452 41364 5462 41420
rect 5518 41364 5528 41420
rect 5452 41354 5528 41364
rect 5576 42908 5652 42918
rect 5576 42852 5586 42908
rect 5642 42852 5652 42908
rect 5576 42784 5652 42852
rect 7552 42888 7562 42944
rect 7618 42888 7686 42944
rect 7742 42888 7810 42944
rect 7866 42888 7934 42944
rect 7990 42888 8058 42944
rect 8114 42888 8182 42944
rect 8238 42888 8306 42944
rect 8362 42888 8430 42944
rect 8486 42888 8554 42944
rect 8610 42888 8620 42944
rect 7552 42820 8620 42888
rect 5576 42728 5586 42784
rect 5642 42728 5652 42784
rect 5576 42660 5652 42728
rect 5576 42604 5586 42660
rect 5642 42604 5652 42660
rect 5576 42536 5652 42604
rect 5576 42480 5586 42536
rect 5642 42480 5652 42536
rect 5576 42412 5652 42480
rect 5576 42356 5586 42412
rect 5642 42356 5652 42412
rect 5576 42288 5652 42356
rect 5576 42232 5586 42288
rect 5642 42232 5652 42288
rect 5576 42164 5652 42232
rect 5576 42108 5586 42164
rect 5642 42108 5652 42164
rect 5576 42040 5652 42108
rect 5576 41984 5586 42040
rect 5642 41984 5652 42040
rect 5576 41916 5652 41984
rect 5576 41860 5586 41916
rect 5642 41860 5652 41916
rect 5576 41792 5652 41860
rect 5576 41736 5586 41792
rect 5642 41736 5652 41792
rect 5576 41668 5652 41736
rect 5576 41612 5586 41668
rect 5642 41612 5652 41668
rect 5576 41544 5652 41612
rect 5576 41488 5586 41544
rect 5642 41488 5652 41544
rect 5576 41420 5652 41488
rect 5576 41364 5586 41420
rect 5642 41364 5652 41420
rect 4832 41237 4842 41293
rect 4898 41237 4908 41293
rect 4832 41169 4908 41237
rect 4832 41113 4842 41169
rect 4898 41113 4908 41169
rect 4832 41045 4908 41113
rect 4832 40989 4842 41045
rect 4898 40989 4908 41045
rect 4832 40921 4908 40989
rect 4832 40865 4842 40921
rect 4898 40865 4908 40921
rect 4832 40797 4908 40865
rect 4832 40741 4842 40797
rect 4898 40741 4908 40797
rect 4832 40673 4908 40741
rect 4832 40617 4842 40673
rect 4898 40617 4908 40673
rect 4832 40549 4908 40617
rect 4832 40493 4842 40549
rect 4898 40493 4908 40549
rect 4832 40425 4908 40493
rect 4832 40369 4842 40425
rect 4898 40369 4908 40425
rect 4832 40301 4908 40369
rect 4832 40245 4842 40301
rect 4898 40245 4908 40301
rect 4832 40177 4908 40245
rect 4832 40121 4842 40177
rect 4898 40121 4908 40177
rect 4832 40053 4908 40121
rect 4832 39997 4842 40053
rect 4898 39997 4908 40053
rect 4832 39929 4908 39997
rect 4832 39873 4842 39929
rect 4898 39873 4908 39929
rect 4832 39805 4908 39873
rect 4832 39749 4842 39805
rect 4898 39749 4908 39805
rect 4832 39739 4908 39749
rect 4956 41293 5032 41303
rect 4956 41237 4966 41293
rect 5022 41237 5032 41293
rect 4956 41169 5032 41237
rect 5576 41296 5652 41364
rect 5576 41240 5586 41296
rect 5642 41240 5652 41296
rect 5576 41230 5652 41240
rect 5700 42784 5776 42794
rect 5700 42728 5710 42784
rect 5766 42728 5776 42784
rect 5700 42660 5776 42728
rect 7552 42764 7562 42820
rect 7618 42764 7686 42820
rect 7742 42764 7810 42820
rect 7866 42764 7934 42820
rect 7990 42764 8058 42820
rect 8114 42764 8182 42820
rect 8238 42764 8306 42820
rect 8362 42764 8430 42820
rect 8486 42764 8554 42820
rect 8610 42764 8620 42820
rect 7552 42696 8620 42764
rect 5700 42604 5710 42660
rect 5766 42604 5776 42660
rect 5700 42536 5776 42604
rect 5700 42480 5710 42536
rect 5766 42480 5776 42536
rect 5700 42412 5776 42480
rect 5700 42356 5710 42412
rect 5766 42356 5776 42412
rect 5700 42288 5776 42356
rect 5700 42232 5710 42288
rect 5766 42232 5776 42288
rect 5700 42164 5776 42232
rect 5700 42108 5710 42164
rect 5766 42108 5776 42164
rect 5700 42040 5776 42108
rect 5700 41984 5710 42040
rect 5766 41984 5776 42040
rect 5700 41916 5776 41984
rect 5700 41860 5710 41916
rect 5766 41860 5776 41916
rect 5700 41792 5776 41860
rect 5700 41736 5710 41792
rect 5766 41736 5776 41792
rect 5700 41668 5776 41736
rect 5700 41612 5710 41668
rect 5766 41612 5776 41668
rect 5700 41544 5776 41612
rect 5700 41488 5710 41544
rect 5766 41488 5776 41544
rect 5700 41420 5776 41488
rect 5700 41364 5710 41420
rect 5766 41364 5776 41420
rect 5700 41296 5776 41364
rect 5700 41240 5710 41296
rect 5766 41240 5776 41296
rect 4956 41113 4966 41169
rect 5022 41113 5032 41169
rect 4956 41045 5032 41113
rect 4956 40989 4966 41045
rect 5022 40989 5032 41045
rect 4956 40921 5032 40989
rect 4956 40865 4966 40921
rect 5022 40865 5032 40921
rect 4956 40797 5032 40865
rect 4956 40741 4966 40797
rect 5022 40741 5032 40797
rect 4956 40673 5032 40741
rect 4956 40617 4966 40673
rect 5022 40617 5032 40673
rect 4956 40549 5032 40617
rect 4956 40493 4966 40549
rect 5022 40493 5032 40549
rect 4956 40425 5032 40493
rect 4956 40369 4966 40425
rect 5022 40369 5032 40425
rect 4956 40301 5032 40369
rect 4956 40245 4966 40301
rect 5022 40245 5032 40301
rect 4956 40177 5032 40245
rect 4956 40121 4966 40177
rect 5022 40121 5032 40177
rect 4956 40053 5032 40121
rect 4956 39997 4966 40053
rect 5022 39997 5032 40053
rect 4956 39929 5032 39997
rect 4956 39873 4966 39929
rect 5022 39873 5032 39929
rect 4956 39805 5032 39873
rect 4956 39749 4966 39805
rect 5022 39749 5032 39805
rect 4956 39681 5032 39749
rect 4956 39625 4966 39681
rect 5022 39625 5032 39681
rect 4956 39615 5032 39625
rect 5080 41169 5156 41179
rect 5080 41113 5090 41169
rect 5146 41113 5156 41169
rect 5080 41045 5156 41113
rect 5700 41172 5776 41240
rect 5700 41116 5710 41172
rect 5766 41116 5776 41172
rect 5700 41106 5776 41116
rect 5824 42660 5900 42670
rect 5824 42604 5834 42660
rect 5890 42604 5900 42660
rect 5824 42536 5900 42604
rect 7552 42640 7562 42696
rect 7618 42640 7686 42696
rect 7742 42640 7810 42696
rect 7866 42640 7934 42696
rect 7990 42640 8058 42696
rect 8114 42640 8182 42696
rect 8238 42640 8306 42696
rect 8362 42640 8430 42696
rect 8486 42640 8554 42696
rect 8610 42640 8620 42696
rect 7552 42572 8620 42640
rect 5824 42480 5834 42536
rect 5890 42480 5900 42536
rect 5824 42412 5900 42480
rect 5824 42356 5834 42412
rect 5890 42356 5900 42412
rect 5824 42288 5900 42356
rect 5824 42232 5834 42288
rect 5890 42232 5900 42288
rect 5824 42164 5900 42232
rect 5824 42108 5834 42164
rect 5890 42108 5900 42164
rect 5824 42040 5900 42108
rect 5824 41984 5834 42040
rect 5890 41984 5900 42040
rect 5824 41916 5900 41984
rect 5824 41860 5834 41916
rect 5890 41860 5900 41916
rect 5824 41792 5900 41860
rect 5824 41736 5834 41792
rect 5890 41736 5900 41792
rect 5824 41668 5900 41736
rect 5824 41612 5834 41668
rect 5890 41612 5900 41668
rect 5824 41544 5900 41612
rect 5824 41488 5834 41544
rect 5890 41488 5900 41544
rect 5824 41420 5900 41488
rect 5824 41364 5834 41420
rect 5890 41364 5900 41420
rect 5824 41296 5900 41364
rect 5824 41240 5834 41296
rect 5890 41240 5900 41296
rect 5824 41172 5900 41240
rect 5824 41116 5834 41172
rect 5890 41116 5900 41172
rect 5080 40989 5090 41045
rect 5146 40989 5156 41045
rect 5080 40921 5156 40989
rect 5080 40865 5090 40921
rect 5146 40865 5156 40921
rect 5080 40797 5156 40865
rect 5080 40741 5090 40797
rect 5146 40741 5156 40797
rect 5080 40673 5156 40741
rect 5080 40617 5090 40673
rect 5146 40617 5156 40673
rect 5080 40549 5156 40617
rect 5080 40493 5090 40549
rect 5146 40493 5156 40549
rect 5080 40425 5156 40493
rect 5080 40369 5090 40425
rect 5146 40369 5156 40425
rect 5080 40301 5156 40369
rect 5080 40245 5090 40301
rect 5146 40245 5156 40301
rect 5080 40177 5156 40245
rect 5080 40121 5090 40177
rect 5146 40121 5156 40177
rect 5080 40053 5156 40121
rect 5080 39997 5090 40053
rect 5146 39997 5156 40053
rect 5080 39929 5156 39997
rect 5080 39873 5090 39929
rect 5146 39873 5156 39929
rect 5080 39805 5156 39873
rect 5080 39749 5090 39805
rect 5146 39749 5156 39805
rect 5080 39681 5156 39749
rect 5080 39625 5090 39681
rect 5146 39625 5156 39681
rect 5080 39557 5156 39625
rect 5080 39501 5090 39557
rect 5146 39501 5156 39557
rect 5080 39491 5156 39501
rect 5204 41045 5280 41055
rect 5204 40989 5214 41045
rect 5270 40989 5280 41045
rect 5204 40921 5280 40989
rect 5824 41048 5900 41116
rect 5824 40992 5834 41048
rect 5890 40992 5900 41048
rect 5824 40982 5900 40992
rect 5948 42536 6024 42546
rect 5948 42480 5958 42536
rect 6014 42480 6024 42536
rect 5948 42412 6024 42480
rect 7552 42516 7562 42572
rect 7618 42516 7686 42572
rect 7742 42516 7810 42572
rect 7866 42516 7934 42572
rect 7990 42516 8058 42572
rect 8114 42516 8182 42572
rect 8238 42516 8306 42572
rect 8362 42516 8430 42572
rect 8486 42516 8554 42572
rect 8610 42516 8620 42572
rect 7552 42448 8620 42516
rect 5948 42356 5958 42412
rect 6014 42356 6024 42412
rect 5948 42288 6024 42356
rect 5948 42232 5958 42288
rect 6014 42232 6024 42288
rect 5948 42164 6024 42232
rect 5948 42108 5958 42164
rect 6014 42108 6024 42164
rect 5948 42040 6024 42108
rect 5948 41984 5958 42040
rect 6014 41984 6024 42040
rect 5948 41916 6024 41984
rect 5948 41860 5958 41916
rect 6014 41860 6024 41916
rect 5948 41792 6024 41860
rect 5948 41736 5958 41792
rect 6014 41736 6024 41792
rect 5948 41668 6024 41736
rect 5948 41612 5958 41668
rect 6014 41612 6024 41668
rect 5948 41544 6024 41612
rect 5948 41488 5958 41544
rect 6014 41488 6024 41544
rect 5948 41420 6024 41488
rect 5948 41364 5958 41420
rect 6014 41364 6024 41420
rect 5948 41296 6024 41364
rect 5948 41240 5958 41296
rect 6014 41240 6024 41296
rect 5948 41172 6024 41240
rect 5948 41116 5958 41172
rect 6014 41116 6024 41172
rect 5948 41048 6024 41116
rect 5948 40992 5958 41048
rect 6014 40992 6024 41048
rect 5204 40865 5214 40921
rect 5270 40865 5280 40921
rect 5204 40797 5280 40865
rect 5204 40741 5214 40797
rect 5270 40741 5280 40797
rect 5204 40673 5280 40741
rect 5204 40617 5214 40673
rect 5270 40617 5280 40673
rect 5204 40549 5280 40617
rect 5204 40493 5214 40549
rect 5270 40493 5280 40549
rect 5204 40425 5280 40493
rect 5204 40369 5214 40425
rect 5270 40369 5280 40425
rect 5204 40301 5280 40369
rect 5204 40245 5214 40301
rect 5270 40245 5280 40301
rect 5204 40177 5280 40245
rect 5204 40121 5214 40177
rect 5270 40121 5280 40177
rect 5204 40053 5280 40121
rect 5204 39997 5214 40053
rect 5270 39997 5280 40053
rect 5204 39929 5280 39997
rect 5204 39873 5214 39929
rect 5270 39873 5280 39929
rect 5204 39805 5280 39873
rect 5204 39749 5214 39805
rect 5270 39749 5280 39805
rect 5204 39681 5280 39749
rect 5204 39625 5214 39681
rect 5270 39625 5280 39681
rect 5204 39557 5280 39625
rect 5204 39501 5214 39557
rect 5270 39501 5280 39557
rect 5204 39433 5280 39501
rect 5204 39377 5214 39433
rect 5270 39377 5280 39433
rect 5204 39367 5280 39377
rect 5328 40921 5404 40931
rect 5328 40865 5338 40921
rect 5394 40865 5404 40921
rect 5328 40797 5404 40865
rect 5948 40924 6024 40992
rect 5948 40868 5958 40924
rect 6014 40868 6024 40924
rect 5948 40858 6024 40868
rect 6072 42412 6148 42422
rect 6072 42356 6082 42412
rect 6138 42356 6148 42412
rect 6072 42288 6148 42356
rect 6072 42232 6082 42288
rect 6138 42232 6148 42288
rect 6072 42164 6148 42232
rect 6072 42108 6082 42164
rect 6138 42108 6148 42164
rect 6072 42040 6148 42108
rect 6072 41984 6082 42040
rect 6138 41984 6148 42040
rect 6072 41916 6148 41984
rect 6072 41860 6082 41916
rect 6138 41860 6148 41916
rect 6072 41792 6148 41860
rect 6072 41736 6082 41792
rect 6138 41736 6148 41792
rect 6072 41668 6148 41736
rect 6072 41612 6082 41668
rect 6138 41612 6148 41668
rect 7552 42392 7562 42448
rect 7618 42392 7686 42448
rect 7742 42392 7810 42448
rect 7866 42392 7934 42448
rect 7990 42392 8058 42448
rect 8114 42392 8182 42448
rect 8238 42392 8306 42448
rect 8362 42392 8430 42448
rect 8486 42392 8554 42448
rect 8610 42392 8620 42448
rect 7552 42324 8620 42392
rect 7552 42268 7562 42324
rect 7618 42268 7686 42324
rect 7742 42268 7810 42324
rect 7866 42268 7934 42324
rect 7990 42268 8058 42324
rect 8114 42268 8182 42324
rect 8238 42268 8306 42324
rect 8362 42268 8430 42324
rect 8486 42268 8554 42324
rect 8610 42268 8620 42324
rect 7552 42200 8620 42268
rect 7552 42144 7562 42200
rect 7618 42144 7686 42200
rect 7742 42144 7810 42200
rect 7866 42144 7934 42200
rect 7990 42144 8058 42200
rect 8114 42144 8182 42200
rect 8238 42144 8306 42200
rect 8362 42144 8430 42200
rect 8486 42144 8554 42200
rect 8610 42144 8620 42200
rect 7552 42076 8620 42144
rect 7552 42020 7562 42076
rect 7618 42020 7686 42076
rect 7742 42020 7810 42076
rect 7866 42020 7934 42076
rect 7990 42020 8058 42076
rect 8114 42020 8182 42076
rect 8238 42020 8306 42076
rect 8362 42020 8430 42076
rect 8486 42020 8554 42076
rect 8610 42020 8620 42076
rect 7552 41952 8620 42020
rect 7552 41896 7562 41952
rect 7618 41896 7686 41952
rect 7742 41896 7810 41952
rect 7866 41896 7934 41952
rect 7990 41896 8058 41952
rect 8114 41896 8182 41952
rect 8238 41896 8306 41952
rect 8362 41896 8430 41952
rect 8486 41896 8554 41952
rect 8610 41896 8620 41952
rect 7552 41828 8620 41896
rect 7552 41772 7562 41828
rect 7618 41772 7686 41828
rect 7742 41772 7810 41828
rect 7866 41772 7934 41828
rect 7990 41772 8058 41828
rect 8114 41772 8182 41828
rect 8238 41772 8306 41828
rect 8362 41772 8430 41828
rect 8486 41772 8554 41828
rect 8610 41772 8620 41828
rect 7552 41704 8620 41772
rect 7552 41648 7562 41704
rect 7618 41648 7686 41704
rect 7742 41648 7810 41704
rect 7866 41648 7934 41704
rect 7990 41648 8058 41704
rect 8114 41648 8182 41704
rect 8238 41648 8306 41704
rect 8362 41648 8430 41704
rect 8486 41648 8554 41704
rect 8610 41648 8620 41704
rect 7552 41638 8620 41648
rect 10669 42944 12481 42954
rect 10669 42888 10679 42944
rect 10735 42888 10803 42944
rect 10859 42888 10927 42944
rect 10983 42888 11051 42944
rect 11107 42888 11175 42944
rect 11231 42888 11299 42944
rect 11355 42888 11423 42944
rect 11479 42888 11547 42944
rect 11603 42888 11671 42944
rect 11727 42888 11795 42944
rect 11851 42888 11919 42944
rect 11975 42888 12043 42944
rect 12099 42888 12167 42944
rect 12223 42888 12291 42944
rect 12347 42888 12415 42944
rect 12471 42888 12481 42944
rect 10669 42820 12481 42888
rect 10669 42764 10679 42820
rect 10735 42764 10803 42820
rect 10859 42764 10927 42820
rect 10983 42764 11051 42820
rect 11107 42764 11175 42820
rect 11231 42764 11299 42820
rect 11355 42764 11423 42820
rect 11479 42764 11547 42820
rect 11603 42764 11671 42820
rect 11727 42764 11795 42820
rect 11851 42764 11919 42820
rect 11975 42764 12043 42820
rect 12099 42764 12167 42820
rect 12223 42764 12291 42820
rect 12347 42764 12415 42820
rect 12471 42764 12481 42820
rect 10669 42696 12481 42764
rect 10669 42640 10679 42696
rect 10735 42640 10803 42696
rect 10859 42640 10927 42696
rect 10983 42640 11051 42696
rect 11107 42640 11175 42696
rect 11231 42640 11299 42696
rect 11355 42640 11423 42696
rect 11479 42640 11547 42696
rect 11603 42640 11671 42696
rect 11727 42640 11795 42696
rect 11851 42640 11919 42696
rect 11975 42640 12043 42696
rect 12099 42640 12167 42696
rect 12223 42640 12291 42696
rect 12347 42640 12415 42696
rect 12471 42640 12481 42696
rect 10669 42572 12481 42640
rect 10669 42516 10679 42572
rect 10735 42516 10803 42572
rect 10859 42516 10927 42572
rect 10983 42516 11051 42572
rect 11107 42516 11175 42572
rect 11231 42516 11299 42572
rect 11355 42516 11423 42572
rect 11479 42516 11547 42572
rect 11603 42516 11671 42572
rect 11727 42516 11795 42572
rect 11851 42516 11919 42572
rect 11975 42516 12043 42572
rect 12099 42516 12167 42572
rect 12223 42516 12291 42572
rect 12347 42516 12415 42572
rect 12471 42516 12481 42572
rect 10669 42448 12481 42516
rect 10669 42392 10679 42448
rect 10735 42392 10803 42448
rect 10859 42392 10927 42448
rect 10983 42392 11051 42448
rect 11107 42392 11175 42448
rect 11231 42392 11299 42448
rect 11355 42392 11423 42448
rect 11479 42392 11547 42448
rect 11603 42392 11671 42448
rect 11727 42392 11795 42448
rect 11851 42392 11919 42448
rect 11975 42392 12043 42448
rect 12099 42392 12167 42448
rect 12223 42392 12291 42448
rect 12347 42392 12415 42448
rect 12471 42392 12481 42448
rect 10669 42324 12481 42392
rect 10669 42268 10679 42324
rect 10735 42268 10803 42324
rect 10859 42268 10927 42324
rect 10983 42268 11051 42324
rect 11107 42268 11175 42324
rect 11231 42268 11299 42324
rect 11355 42268 11423 42324
rect 11479 42268 11547 42324
rect 11603 42268 11671 42324
rect 11727 42268 11795 42324
rect 11851 42268 11919 42324
rect 11975 42268 12043 42324
rect 12099 42268 12167 42324
rect 12223 42268 12291 42324
rect 12347 42268 12415 42324
rect 12471 42268 12481 42324
rect 10669 42200 12481 42268
rect 10669 42144 10679 42200
rect 10735 42144 10803 42200
rect 10859 42144 10927 42200
rect 10983 42144 11051 42200
rect 11107 42144 11175 42200
rect 11231 42144 11299 42200
rect 11355 42144 11423 42200
rect 11479 42144 11547 42200
rect 11603 42144 11671 42200
rect 11727 42144 11795 42200
rect 11851 42144 11919 42200
rect 11975 42144 12043 42200
rect 12099 42144 12167 42200
rect 12223 42144 12291 42200
rect 12347 42144 12415 42200
rect 12471 42144 12481 42200
rect 10669 42076 12481 42144
rect 10669 42020 10679 42076
rect 10735 42020 10803 42076
rect 10859 42020 10927 42076
rect 10983 42020 11051 42076
rect 11107 42020 11175 42076
rect 11231 42020 11299 42076
rect 11355 42020 11423 42076
rect 11479 42020 11547 42076
rect 11603 42020 11671 42076
rect 11727 42020 11795 42076
rect 11851 42020 11919 42076
rect 11975 42020 12043 42076
rect 12099 42020 12167 42076
rect 12223 42020 12291 42076
rect 12347 42020 12415 42076
rect 12471 42020 12481 42076
rect 10669 41952 12481 42020
rect 10669 41896 10679 41952
rect 10735 41896 10803 41952
rect 10859 41896 10927 41952
rect 10983 41896 11051 41952
rect 11107 41896 11175 41952
rect 11231 41896 11299 41952
rect 11355 41896 11423 41952
rect 11479 41896 11547 41952
rect 11603 41896 11671 41952
rect 11727 41896 11795 41952
rect 11851 41896 11919 41952
rect 11975 41896 12043 41952
rect 12099 41896 12167 41952
rect 12223 41896 12291 41952
rect 12347 41896 12415 41952
rect 12471 41896 12481 41952
rect 10669 41828 12481 41896
rect 10669 41772 10679 41828
rect 10735 41772 10803 41828
rect 10859 41772 10927 41828
rect 10983 41772 11051 41828
rect 11107 41772 11175 41828
rect 11231 41772 11299 41828
rect 11355 41772 11423 41828
rect 11479 41772 11547 41828
rect 11603 41772 11671 41828
rect 11727 41772 11795 41828
rect 11851 41772 11919 41828
rect 11975 41772 12043 41828
rect 12099 41772 12167 41828
rect 12223 41772 12291 41828
rect 12347 41772 12415 41828
rect 12471 41772 12481 41828
rect 10669 41704 12481 41772
rect 10669 41648 10679 41704
rect 10735 41648 10803 41704
rect 10859 41648 10927 41704
rect 10983 41648 11051 41704
rect 11107 41648 11175 41704
rect 11231 41648 11299 41704
rect 11355 41648 11423 41704
rect 11479 41648 11547 41704
rect 11603 41648 11671 41704
rect 11727 41648 11795 41704
rect 11851 41648 11919 41704
rect 11975 41648 12043 41704
rect 12099 41648 12167 41704
rect 12223 41648 12291 41704
rect 12347 41648 12415 41704
rect 12471 41648 12481 41704
rect 10669 41638 12481 41648
rect 6072 41544 6148 41612
rect 6072 41488 6082 41544
rect 6138 41488 6148 41544
rect 6072 41420 6148 41488
rect 6072 41364 6082 41420
rect 6138 41364 6148 41420
rect 6072 41296 6148 41364
rect 6072 41240 6082 41296
rect 6138 41240 6148 41296
rect 6072 41172 6148 41240
rect 6072 41116 6082 41172
rect 6138 41116 6148 41172
rect 6072 41048 6148 41116
rect 6072 40992 6082 41048
rect 6138 40992 6148 41048
rect 6072 40924 6148 40992
rect 6072 40868 6082 40924
rect 6138 40868 6148 40924
rect 5328 40741 5338 40797
rect 5394 40741 5404 40797
rect 5328 40673 5404 40741
rect 5328 40617 5338 40673
rect 5394 40617 5404 40673
rect 5328 40549 5404 40617
rect 5328 40493 5338 40549
rect 5394 40493 5404 40549
rect 5328 40425 5404 40493
rect 5328 40369 5338 40425
rect 5394 40369 5404 40425
rect 5328 40301 5404 40369
rect 5328 40245 5338 40301
rect 5394 40245 5404 40301
rect 5328 40177 5404 40245
rect 5328 40121 5338 40177
rect 5394 40121 5404 40177
rect 5328 40053 5404 40121
rect 5328 39997 5338 40053
rect 5394 39997 5404 40053
rect 5328 39929 5404 39997
rect 5328 39873 5338 39929
rect 5394 39873 5404 39929
rect 5328 39805 5404 39873
rect 5328 39749 5338 39805
rect 5394 39749 5404 39805
rect 5328 39681 5404 39749
rect 5328 39625 5338 39681
rect 5394 39625 5404 39681
rect 5328 39557 5404 39625
rect 5328 39501 5338 39557
rect 5394 39501 5404 39557
rect 5328 39433 5404 39501
rect 5328 39377 5338 39433
rect 5394 39377 5404 39433
rect 5328 39309 5404 39377
rect 5328 39253 5338 39309
rect 5394 39253 5404 39309
rect 5328 39243 5404 39253
rect 5452 40797 5528 40807
rect 5452 40741 5462 40797
rect 5518 40741 5528 40797
rect 5452 40673 5528 40741
rect 6072 40800 6148 40868
rect 6072 40744 6082 40800
rect 6138 40744 6148 40800
rect 6072 40734 6148 40744
rect 7552 41344 8620 41354
rect 7552 41288 7562 41344
rect 7618 41288 7686 41344
rect 7742 41288 7810 41344
rect 7866 41288 7934 41344
rect 7990 41288 8058 41344
rect 8114 41288 8182 41344
rect 8238 41288 8306 41344
rect 8362 41288 8430 41344
rect 8486 41288 8554 41344
rect 8610 41288 8620 41344
rect 7552 41220 8620 41288
rect 7552 41164 7562 41220
rect 7618 41164 7686 41220
rect 7742 41164 7810 41220
rect 7866 41164 7934 41220
rect 7990 41164 8058 41220
rect 8114 41164 8182 41220
rect 8238 41164 8306 41220
rect 8362 41164 8430 41220
rect 8486 41164 8554 41220
rect 8610 41164 8620 41220
rect 7552 41096 8620 41164
rect 7552 41040 7562 41096
rect 7618 41040 7686 41096
rect 7742 41040 7810 41096
rect 7866 41040 7934 41096
rect 7990 41040 8058 41096
rect 8114 41040 8182 41096
rect 8238 41040 8306 41096
rect 8362 41040 8430 41096
rect 8486 41040 8554 41096
rect 8610 41040 8620 41096
rect 7552 40972 8620 41040
rect 7552 40916 7562 40972
rect 7618 40916 7686 40972
rect 7742 40916 7810 40972
rect 7866 40916 7934 40972
rect 7990 40916 8058 40972
rect 8114 40916 8182 40972
rect 8238 40916 8306 40972
rect 8362 40916 8430 40972
rect 8486 40916 8554 40972
rect 8610 40916 8620 40972
rect 7552 40848 8620 40916
rect 7552 40792 7562 40848
rect 7618 40792 7686 40848
rect 7742 40792 7810 40848
rect 7866 40792 7934 40848
rect 7990 40792 8058 40848
rect 8114 40792 8182 40848
rect 8238 40792 8306 40848
rect 8362 40792 8430 40848
rect 8486 40792 8554 40848
rect 8610 40792 8620 40848
rect 7552 40724 8620 40792
rect 5452 40617 5462 40673
rect 5518 40617 5528 40673
rect 5452 40549 5528 40617
rect 5452 40493 5462 40549
rect 5518 40493 5528 40549
rect 5452 40425 5528 40493
rect 5452 40369 5462 40425
rect 5518 40369 5528 40425
rect 5452 40301 5528 40369
rect 5452 40245 5462 40301
rect 5518 40245 5528 40301
rect 5452 40177 5528 40245
rect 5452 40121 5462 40177
rect 5518 40121 5528 40177
rect 5452 40053 5528 40121
rect 5452 39997 5462 40053
rect 5518 39997 5528 40053
rect 5452 39929 5528 39997
rect 5452 39873 5462 39929
rect 5518 39873 5528 39929
rect 5452 39805 5528 39873
rect 5452 39749 5462 39805
rect 5518 39749 5528 39805
rect 5452 39681 5528 39749
rect 5452 39625 5462 39681
rect 5518 39625 5528 39681
rect 5452 39557 5528 39625
rect 5452 39501 5462 39557
rect 5518 39501 5528 39557
rect 5452 39433 5528 39501
rect 5452 39377 5462 39433
rect 5518 39377 5528 39433
rect 5452 39309 5528 39377
rect 5452 39253 5462 39309
rect 5518 39253 5528 39309
rect 5452 39185 5528 39253
rect 5452 39129 5462 39185
rect 5518 39129 5528 39185
rect 5452 39119 5528 39129
rect 5576 40673 5652 40683
rect 5576 40617 5586 40673
rect 5642 40617 5652 40673
rect 5576 40549 5652 40617
rect 7552 40668 7562 40724
rect 7618 40668 7686 40724
rect 7742 40668 7810 40724
rect 7866 40668 7934 40724
rect 7990 40668 8058 40724
rect 8114 40668 8182 40724
rect 8238 40668 8306 40724
rect 8362 40668 8430 40724
rect 8486 40668 8554 40724
rect 8610 40668 8620 40724
rect 7552 40600 8620 40668
rect 5576 40493 5586 40549
rect 5642 40493 5652 40549
rect 5576 40425 5652 40493
rect 5576 40369 5586 40425
rect 5642 40369 5652 40425
rect 5576 40301 5652 40369
rect 5576 40245 5586 40301
rect 5642 40245 5652 40301
rect 5576 40177 5652 40245
rect 5576 40121 5586 40177
rect 5642 40121 5652 40177
rect 5576 40053 5652 40121
rect 5576 39997 5586 40053
rect 5642 39997 5652 40053
rect 5576 39929 5652 39997
rect 5576 39873 5586 39929
rect 5642 39873 5652 39929
rect 5576 39805 5652 39873
rect 5576 39749 5586 39805
rect 5642 39749 5652 39805
rect 5576 39681 5652 39749
rect 5576 39625 5586 39681
rect 5642 39625 5652 39681
rect 5576 39557 5652 39625
rect 5576 39501 5586 39557
rect 5642 39501 5652 39557
rect 5576 39433 5652 39501
rect 5576 39377 5586 39433
rect 5642 39377 5652 39433
rect 5576 39309 5652 39377
rect 5576 39253 5586 39309
rect 5642 39253 5652 39309
rect 5576 39185 5652 39253
rect 5576 39129 5586 39185
rect 5642 39129 5652 39185
rect 5576 39061 5652 39129
rect 5576 39005 5586 39061
rect 5642 39005 5652 39061
rect 5576 38995 5652 39005
rect 5700 40549 5776 40559
rect 5700 40493 5710 40549
rect 5766 40493 5776 40549
rect 5700 40425 5776 40493
rect 7552 40544 7562 40600
rect 7618 40544 7686 40600
rect 7742 40544 7810 40600
rect 7866 40544 7934 40600
rect 7990 40544 8058 40600
rect 8114 40544 8182 40600
rect 8238 40544 8306 40600
rect 8362 40544 8430 40600
rect 8486 40544 8554 40600
rect 8610 40544 8620 40600
rect 7552 40476 8620 40544
rect 5700 40369 5710 40425
rect 5766 40369 5776 40425
rect 5700 40301 5776 40369
rect 5700 40245 5710 40301
rect 5766 40245 5776 40301
rect 5700 40177 5776 40245
rect 5700 40121 5710 40177
rect 5766 40121 5776 40177
rect 5700 40053 5776 40121
rect 5700 39997 5710 40053
rect 5766 39997 5776 40053
rect 5700 39929 5776 39997
rect 5700 39873 5710 39929
rect 5766 39873 5776 39929
rect 5700 39805 5776 39873
rect 5700 39749 5710 39805
rect 5766 39749 5776 39805
rect 5700 39681 5776 39749
rect 5700 39625 5710 39681
rect 5766 39625 5776 39681
rect 5700 39557 5776 39625
rect 5700 39501 5710 39557
rect 5766 39501 5776 39557
rect 5700 39433 5776 39501
rect 5700 39377 5710 39433
rect 5766 39377 5776 39433
rect 5700 39309 5776 39377
rect 5700 39253 5710 39309
rect 5766 39253 5776 39309
rect 5700 39185 5776 39253
rect 5700 39129 5710 39185
rect 5766 39129 5776 39185
rect 5700 39061 5776 39129
rect 5700 39005 5710 39061
rect 5766 39005 5776 39061
rect 5700 38937 5776 39005
rect 5700 38881 5710 38937
rect 5766 38881 5776 38937
rect 5700 38871 5776 38881
rect 5824 40425 5900 40435
rect 5824 40369 5834 40425
rect 5890 40369 5900 40425
rect 5824 40301 5900 40369
rect 7552 40420 7562 40476
rect 7618 40420 7686 40476
rect 7742 40420 7810 40476
rect 7866 40420 7934 40476
rect 7990 40420 8058 40476
rect 8114 40420 8182 40476
rect 8238 40420 8306 40476
rect 8362 40420 8430 40476
rect 8486 40420 8554 40476
rect 8610 40420 8620 40476
rect 7552 40352 8620 40420
rect 5824 40245 5834 40301
rect 5890 40245 5900 40301
rect 5824 40177 5900 40245
rect 5824 40121 5834 40177
rect 5890 40121 5900 40177
rect 5824 40053 5900 40121
rect 5824 39997 5834 40053
rect 5890 39997 5900 40053
rect 5824 39929 5900 39997
rect 5824 39873 5834 39929
rect 5890 39873 5900 39929
rect 5824 39805 5900 39873
rect 5824 39749 5834 39805
rect 5890 39749 5900 39805
rect 5824 39681 5900 39749
rect 5824 39625 5834 39681
rect 5890 39625 5900 39681
rect 5824 39557 5900 39625
rect 5824 39501 5834 39557
rect 5890 39501 5900 39557
rect 5824 39433 5900 39501
rect 5824 39377 5834 39433
rect 5890 39377 5900 39433
rect 5824 39309 5900 39377
rect 5824 39253 5834 39309
rect 5890 39253 5900 39309
rect 5824 39185 5900 39253
rect 5824 39129 5834 39185
rect 5890 39129 5900 39185
rect 5824 39061 5900 39129
rect 5824 39005 5834 39061
rect 5890 39005 5900 39061
rect 5824 38937 5900 39005
rect 5824 38881 5834 38937
rect 5890 38881 5900 38937
rect 5824 38813 5900 38881
rect 5824 38757 5834 38813
rect 5890 38757 5900 38813
rect 5824 38747 5900 38757
rect 5948 40301 6024 40311
rect 5948 40245 5958 40301
rect 6014 40245 6024 40301
rect 5948 40177 6024 40245
rect 7552 40296 7562 40352
rect 7618 40296 7686 40352
rect 7742 40296 7810 40352
rect 7866 40296 7934 40352
rect 7990 40296 8058 40352
rect 8114 40296 8182 40352
rect 8238 40296 8306 40352
rect 8362 40296 8430 40352
rect 8486 40296 8554 40352
rect 8610 40296 8620 40352
rect 7552 40228 8620 40296
rect 5948 40121 5958 40177
rect 6014 40121 6024 40177
rect 5948 40053 6024 40121
rect 5948 39997 5958 40053
rect 6014 39997 6024 40053
rect 5948 39929 6024 39997
rect 5948 39873 5958 39929
rect 6014 39873 6024 39929
rect 5948 39805 6024 39873
rect 5948 39749 5958 39805
rect 6014 39749 6024 39805
rect 5948 39681 6024 39749
rect 5948 39625 5958 39681
rect 6014 39625 6024 39681
rect 5948 39557 6024 39625
rect 5948 39501 5958 39557
rect 6014 39501 6024 39557
rect 5948 39433 6024 39501
rect 5948 39377 5958 39433
rect 6014 39377 6024 39433
rect 5948 39309 6024 39377
rect 5948 39253 5958 39309
rect 6014 39253 6024 39309
rect 5948 39185 6024 39253
rect 5948 39129 5958 39185
rect 6014 39129 6024 39185
rect 5948 39061 6024 39129
rect 5948 39005 5958 39061
rect 6014 39005 6024 39061
rect 5948 38937 6024 39005
rect 5948 38881 5958 38937
rect 6014 38881 6024 38937
rect 5948 38813 6024 38881
rect 5948 38757 5958 38813
rect 6014 38757 6024 38813
rect 5948 38689 6024 38757
rect 5948 38633 5958 38689
rect 6014 38633 6024 38689
rect 5948 38623 6024 38633
rect 6072 40177 6148 40187
rect 6072 40121 6082 40177
rect 6138 40121 6148 40177
rect 6072 40053 6148 40121
rect 6072 39997 6082 40053
rect 6138 39997 6148 40053
rect 7552 40172 7562 40228
rect 7618 40172 7686 40228
rect 7742 40172 7810 40228
rect 7866 40172 7934 40228
rect 7990 40172 8058 40228
rect 8114 40172 8182 40228
rect 8238 40172 8306 40228
rect 8362 40172 8430 40228
rect 8486 40172 8554 40228
rect 8610 40172 8620 40228
rect 7552 40104 8620 40172
rect 7552 40048 7562 40104
rect 7618 40048 7686 40104
rect 7742 40048 7810 40104
rect 7866 40048 7934 40104
rect 7990 40048 8058 40104
rect 8114 40048 8182 40104
rect 8238 40048 8306 40104
rect 8362 40048 8430 40104
rect 8486 40048 8554 40104
rect 8610 40048 8620 40104
rect 7552 40038 8620 40048
rect 10669 41344 12481 41354
rect 10669 41288 10679 41344
rect 10735 41288 10803 41344
rect 10859 41288 10927 41344
rect 10983 41288 11051 41344
rect 11107 41288 11175 41344
rect 11231 41288 11299 41344
rect 11355 41288 11423 41344
rect 11479 41288 11547 41344
rect 11603 41288 11671 41344
rect 11727 41288 11795 41344
rect 11851 41288 11919 41344
rect 11975 41288 12043 41344
rect 12099 41288 12167 41344
rect 12223 41288 12291 41344
rect 12347 41288 12415 41344
rect 12471 41288 12481 41344
rect 10669 41220 12481 41288
rect 10669 41164 10679 41220
rect 10735 41164 10803 41220
rect 10859 41164 10927 41220
rect 10983 41164 11051 41220
rect 11107 41164 11175 41220
rect 11231 41164 11299 41220
rect 11355 41164 11423 41220
rect 11479 41164 11547 41220
rect 11603 41164 11671 41220
rect 11727 41164 11795 41220
rect 11851 41164 11919 41220
rect 11975 41164 12043 41220
rect 12099 41164 12167 41220
rect 12223 41164 12291 41220
rect 12347 41164 12415 41220
rect 12471 41164 12481 41220
rect 10669 41096 12481 41164
rect 10669 41040 10679 41096
rect 10735 41040 10803 41096
rect 10859 41040 10927 41096
rect 10983 41040 11051 41096
rect 11107 41040 11175 41096
rect 11231 41040 11299 41096
rect 11355 41040 11423 41096
rect 11479 41040 11547 41096
rect 11603 41040 11671 41096
rect 11727 41040 11795 41096
rect 11851 41040 11919 41096
rect 11975 41040 12043 41096
rect 12099 41040 12167 41096
rect 12223 41040 12291 41096
rect 12347 41040 12415 41096
rect 12471 41040 12481 41096
rect 10669 40972 12481 41040
rect 10669 40916 10679 40972
rect 10735 40916 10803 40972
rect 10859 40916 10927 40972
rect 10983 40916 11051 40972
rect 11107 40916 11175 40972
rect 11231 40916 11299 40972
rect 11355 40916 11423 40972
rect 11479 40916 11547 40972
rect 11603 40916 11671 40972
rect 11727 40916 11795 40972
rect 11851 40916 11919 40972
rect 11975 40916 12043 40972
rect 12099 40916 12167 40972
rect 12223 40916 12291 40972
rect 12347 40916 12415 40972
rect 12471 40916 12481 40972
rect 10669 40848 12481 40916
rect 10669 40792 10679 40848
rect 10735 40792 10803 40848
rect 10859 40792 10927 40848
rect 10983 40792 11051 40848
rect 11107 40792 11175 40848
rect 11231 40792 11299 40848
rect 11355 40792 11423 40848
rect 11479 40792 11547 40848
rect 11603 40792 11671 40848
rect 11727 40792 11795 40848
rect 11851 40792 11919 40848
rect 11975 40792 12043 40848
rect 12099 40792 12167 40848
rect 12223 40792 12291 40848
rect 12347 40792 12415 40848
rect 12471 40792 12481 40848
rect 10669 40724 12481 40792
rect 10669 40668 10679 40724
rect 10735 40668 10803 40724
rect 10859 40668 10927 40724
rect 10983 40668 11051 40724
rect 11107 40668 11175 40724
rect 11231 40668 11299 40724
rect 11355 40668 11423 40724
rect 11479 40668 11547 40724
rect 11603 40668 11671 40724
rect 11727 40668 11795 40724
rect 11851 40668 11919 40724
rect 11975 40668 12043 40724
rect 12099 40668 12167 40724
rect 12223 40668 12291 40724
rect 12347 40668 12415 40724
rect 12471 40668 12481 40724
rect 10669 40600 12481 40668
rect 10669 40544 10679 40600
rect 10735 40544 10803 40600
rect 10859 40544 10927 40600
rect 10983 40544 11051 40600
rect 11107 40544 11175 40600
rect 11231 40544 11299 40600
rect 11355 40544 11423 40600
rect 11479 40544 11547 40600
rect 11603 40544 11671 40600
rect 11727 40544 11795 40600
rect 11851 40544 11919 40600
rect 11975 40544 12043 40600
rect 12099 40544 12167 40600
rect 12223 40544 12291 40600
rect 12347 40544 12415 40600
rect 12471 40544 12481 40600
rect 10669 40476 12481 40544
rect 10669 40420 10679 40476
rect 10735 40420 10803 40476
rect 10859 40420 10927 40476
rect 10983 40420 11051 40476
rect 11107 40420 11175 40476
rect 11231 40420 11299 40476
rect 11355 40420 11423 40476
rect 11479 40420 11547 40476
rect 11603 40420 11671 40476
rect 11727 40420 11795 40476
rect 11851 40420 11919 40476
rect 11975 40420 12043 40476
rect 12099 40420 12167 40476
rect 12223 40420 12291 40476
rect 12347 40420 12415 40476
rect 12471 40420 12481 40476
rect 10669 40352 12481 40420
rect 10669 40296 10679 40352
rect 10735 40296 10803 40352
rect 10859 40296 10927 40352
rect 10983 40296 11051 40352
rect 11107 40296 11175 40352
rect 11231 40296 11299 40352
rect 11355 40296 11423 40352
rect 11479 40296 11547 40352
rect 11603 40296 11671 40352
rect 11727 40296 11795 40352
rect 11851 40296 11919 40352
rect 11975 40296 12043 40352
rect 12099 40296 12167 40352
rect 12223 40296 12291 40352
rect 12347 40296 12415 40352
rect 12471 40296 12481 40352
rect 10669 40228 12481 40296
rect 10669 40172 10679 40228
rect 10735 40172 10803 40228
rect 10859 40172 10927 40228
rect 10983 40172 11051 40228
rect 11107 40172 11175 40228
rect 11231 40172 11299 40228
rect 11355 40172 11423 40228
rect 11479 40172 11547 40228
rect 11603 40172 11671 40228
rect 11727 40172 11795 40228
rect 11851 40172 11919 40228
rect 11975 40172 12043 40228
rect 12099 40172 12167 40228
rect 12223 40172 12291 40228
rect 12347 40172 12415 40228
rect 12471 40172 12481 40228
rect 10669 40104 12481 40172
rect 10669 40048 10679 40104
rect 10735 40048 10803 40104
rect 10859 40048 10927 40104
rect 10983 40048 11051 40104
rect 11107 40048 11175 40104
rect 11231 40048 11299 40104
rect 11355 40048 11423 40104
rect 11479 40048 11547 40104
rect 11603 40048 11671 40104
rect 11727 40048 11795 40104
rect 11851 40048 11919 40104
rect 11975 40048 12043 40104
rect 12099 40048 12167 40104
rect 12223 40048 12291 40104
rect 12347 40048 12415 40104
rect 12471 40048 12481 40104
rect 10669 40038 12481 40048
rect 6072 39929 6148 39997
rect 6072 39873 6082 39929
rect 6138 39873 6148 39929
rect 6072 39805 6148 39873
rect 6072 39749 6082 39805
rect 6138 39749 6148 39805
rect 6072 39681 6148 39749
rect 6072 39625 6082 39681
rect 6138 39625 6148 39681
rect 6072 39557 6148 39625
rect 6072 39501 6082 39557
rect 6138 39501 6148 39557
rect 6072 39433 6148 39501
rect 6072 39377 6082 39433
rect 6138 39377 6148 39433
rect 6072 39309 6148 39377
rect 6072 39253 6082 39309
rect 6138 39253 6148 39309
rect 6072 39185 6148 39253
rect 6072 39129 6082 39185
rect 6138 39129 6148 39185
rect 6072 39061 6148 39129
rect 6072 39005 6082 39061
rect 6138 39005 6148 39061
rect 6072 38937 6148 39005
rect 6072 38881 6082 38937
rect 6138 38881 6148 38937
rect 6072 38813 6148 38881
rect 6072 38757 6082 38813
rect 6138 38757 6148 38813
rect 6072 38689 6148 38757
rect 6072 38633 6082 38689
rect 6138 38633 6148 38689
rect 6072 38565 6148 38633
rect 6072 38509 6082 38565
rect 6138 38509 6148 38565
rect 6072 38499 6148 38509
rect 7552 39744 8620 39754
rect 7552 39688 7562 39744
rect 7618 39688 7686 39744
rect 7742 39688 7810 39744
rect 7866 39688 7934 39744
rect 7990 39688 8058 39744
rect 8114 39688 8182 39744
rect 8238 39688 8306 39744
rect 8362 39688 8430 39744
rect 8486 39688 8554 39744
rect 8610 39688 8620 39744
rect 7552 39620 8620 39688
rect 7552 39564 7562 39620
rect 7618 39564 7686 39620
rect 7742 39564 7810 39620
rect 7866 39564 7934 39620
rect 7990 39564 8058 39620
rect 8114 39564 8182 39620
rect 8238 39564 8306 39620
rect 8362 39564 8430 39620
rect 8486 39564 8554 39620
rect 8610 39564 8620 39620
rect 7552 39496 8620 39564
rect 7552 39440 7562 39496
rect 7618 39440 7686 39496
rect 7742 39440 7810 39496
rect 7866 39440 7934 39496
rect 7990 39440 8058 39496
rect 8114 39440 8182 39496
rect 8238 39440 8306 39496
rect 8362 39440 8430 39496
rect 8486 39440 8554 39496
rect 8610 39440 8620 39496
rect 7552 39372 8620 39440
rect 7552 39316 7562 39372
rect 7618 39316 7686 39372
rect 7742 39316 7810 39372
rect 7866 39316 7934 39372
rect 7990 39316 8058 39372
rect 8114 39316 8182 39372
rect 8238 39316 8306 39372
rect 8362 39316 8430 39372
rect 8486 39316 8554 39372
rect 8610 39316 8620 39372
rect 7552 39248 8620 39316
rect 7552 39192 7562 39248
rect 7618 39192 7686 39248
rect 7742 39192 7810 39248
rect 7866 39192 7934 39248
rect 7990 39192 8058 39248
rect 8114 39192 8182 39248
rect 8238 39192 8306 39248
rect 8362 39192 8430 39248
rect 8486 39192 8554 39248
rect 8610 39192 8620 39248
rect 7552 39124 8620 39192
rect 7552 39068 7562 39124
rect 7618 39068 7686 39124
rect 7742 39068 7810 39124
rect 7866 39068 7934 39124
rect 7990 39068 8058 39124
rect 8114 39068 8182 39124
rect 8238 39068 8306 39124
rect 8362 39068 8430 39124
rect 8486 39068 8554 39124
rect 8610 39068 8620 39124
rect 7552 39000 8620 39068
rect 7552 38944 7562 39000
rect 7618 38944 7686 39000
rect 7742 38944 7810 39000
rect 7866 38944 7934 39000
rect 7990 38944 8058 39000
rect 8114 38944 8182 39000
rect 8238 38944 8306 39000
rect 8362 38944 8430 39000
rect 8486 38944 8554 39000
rect 8610 38944 8620 39000
rect 7552 38876 8620 38944
rect 7552 38820 7562 38876
rect 7618 38820 7686 38876
rect 7742 38820 7810 38876
rect 7866 38820 7934 38876
rect 7990 38820 8058 38876
rect 8114 38820 8182 38876
rect 8238 38820 8306 38876
rect 8362 38820 8430 38876
rect 8486 38820 8554 38876
rect 8610 38820 8620 38876
rect 7552 38752 8620 38820
rect 7552 38696 7562 38752
rect 7618 38696 7686 38752
rect 7742 38696 7810 38752
rect 7866 38696 7934 38752
rect 7990 38696 8058 38752
rect 8114 38696 8182 38752
rect 8238 38696 8306 38752
rect 8362 38696 8430 38752
rect 8486 38696 8554 38752
rect 8610 38696 8620 38752
rect 7552 38628 8620 38696
rect 7552 38572 7562 38628
rect 7618 38572 7686 38628
rect 7742 38572 7810 38628
rect 7866 38572 7934 38628
rect 7990 38572 8058 38628
rect 8114 38572 8182 38628
rect 8238 38572 8306 38628
rect 8362 38572 8430 38628
rect 8486 38572 8554 38628
rect 8610 38572 8620 38628
rect 7552 38504 8620 38572
rect 7552 38448 7562 38504
rect 7618 38448 7686 38504
rect 7742 38448 7810 38504
rect 7866 38448 7934 38504
rect 7990 38448 8058 38504
rect 8114 38448 8182 38504
rect 8238 38448 8306 38504
rect 8362 38448 8430 38504
rect 8486 38448 8554 38504
rect 8610 38448 8620 38504
rect 7552 38438 8620 38448
rect 10669 39744 12481 39754
rect 10669 39688 10679 39744
rect 10735 39688 10803 39744
rect 10859 39688 10927 39744
rect 10983 39688 11051 39744
rect 11107 39688 11175 39744
rect 11231 39688 11299 39744
rect 11355 39688 11423 39744
rect 11479 39688 11547 39744
rect 11603 39688 11671 39744
rect 11727 39688 11795 39744
rect 11851 39688 11919 39744
rect 11975 39688 12043 39744
rect 12099 39688 12167 39744
rect 12223 39688 12291 39744
rect 12347 39688 12415 39744
rect 12471 39688 12481 39744
rect 10669 39620 12481 39688
rect 10669 39564 10679 39620
rect 10735 39564 10803 39620
rect 10859 39564 10927 39620
rect 10983 39564 11051 39620
rect 11107 39564 11175 39620
rect 11231 39564 11299 39620
rect 11355 39564 11423 39620
rect 11479 39564 11547 39620
rect 11603 39564 11671 39620
rect 11727 39564 11795 39620
rect 11851 39564 11919 39620
rect 11975 39564 12043 39620
rect 12099 39564 12167 39620
rect 12223 39564 12291 39620
rect 12347 39564 12415 39620
rect 12471 39564 12481 39620
rect 10669 39496 12481 39564
rect 10669 39440 10679 39496
rect 10735 39440 10803 39496
rect 10859 39440 10927 39496
rect 10983 39440 11051 39496
rect 11107 39440 11175 39496
rect 11231 39440 11299 39496
rect 11355 39440 11423 39496
rect 11479 39440 11547 39496
rect 11603 39440 11671 39496
rect 11727 39440 11795 39496
rect 11851 39440 11919 39496
rect 11975 39440 12043 39496
rect 12099 39440 12167 39496
rect 12223 39440 12291 39496
rect 12347 39440 12415 39496
rect 12471 39440 12481 39496
rect 10669 39372 12481 39440
rect 10669 39316 10679 39372
rect 10735 39316 10803 39372
rect 10859 39316 10927 39372
rect 10983 39316 11051 39372
rect 11107 39316 11175 39372
rect 11231 39316 11299 39372
rect 11355 39316 11423 39372
rect 11479 39316 11547 39372
rect 11603 39316 11671 39372
rect 11727 39316 11795 39372
rect 11851 39316 11919 39372
rect 11975 39316 12043 39372
rect 12099 39316 12167 39372
rect 12223 39316 12291 39372
rect 12347 39316 12415 39372
rect 12471 39316 12481 39372
rect 10669 39248 12481 39316
rect 10669 39192 10679 39248
rect 10735 39192 10803 39248
rect 10859 39192 10927 39248
rect 10983 39192 11051 39248
rect 11107 39192 11175 39248
rect 11231 39192 11299 39248
rect 11355 39192 11423 39248
rect 11479 39192 11547 39248
rect 11603 39192 11671 39248
rect 11727 39192 11795 39248
rect 11851 39192 11919 39248
rect 11975 39192 12043 39248
rect 12099 39192 12167 39248
rect 12223 39192 12291 39248
rect 12347 39192 12415 39248
rect 12471 39192 12481 39248
rect 10669 39124 12481 39192
rect 10669 39068 10679 39124
rect 10735 39068 10803 39124
rect 10859 39068 10927 39124
rect 10983 39068 11051 39124
rect 11107 39068 11175 39124
rect 11231 39068 11299 39124
rect 11355 39068 11423 39124
rect 11479 39068 11547 39124
rect 11603 39068 11671 39124
rect 11727 39068 11795 39124
rect 11851 39068 11919 39124
rect 11975 39068 12043 39124
rect 12099 39068 12167 39124
rect 12223 39068 12291 39124
rect 12347 39068 12415 39124
rect 12471 39068 12481 39124
rect 10669 39000 12481 39068
rect 10669 38944 10679 39000
rect 10735 38944 10803 39000
rect 10859 38944 10927 39000
rect 10983 38944 11051 39000
rect 11107 38944 11175 39000
rect 11231 38944 11299 39000
rect 11355 38944 11423 39000
rect 11479 38944 11547 39000
rect 11603 38944 11671 39000
rect 11727 38944 11795 39000
rect 11851 38944 11919 39000
rect 11975 38944 12043 39000
rect 12099 38944 12167 39000
rect 12223 38944 12291 39000
rect 12347 38944 12415 39000
rect 12471 38944 12481 39000
rect 10669 38876 12481 38944
rect 10669 38820 10679 38876
rect 10735 38820 10803 38876
rect 10859 38820 10927 38876
rect 10983 38820 11051 38876
rect 11107 38820 11175 38876
rect 11231 38820 11299 38876
rect 11355 38820 11423 38876
rect 11479 38820 11547 38876
rect 11603 38820 11671 38876
rect 11727 38820 11795 38876
rect 11851 38820 11919 38876
rect 11975 38820 12043 38876
rect 12099 38820 12167 38876
rect 12223 38820 12291 38876
rect 12347 38820 12415 38876
rect 12471 38820 12481 38876
rect 10669 38752 12481 38820
rect 10669 38696 10679 38752
rect 10735 38696 10803 38752
rect 10859 38696 10927 38752
rect 10983 38696 11051 38752
rect 11107 38696 11175 38752
rect 11231 38696 11299 38752
rect 11355 38696 11423 38752
rect 11479 38696 11547 38752
rect 11603 38696 11671 38752
rect 11727 38696 11795 38752
rect 11851 38696 11919 38752
rect 11975 38696 12043 38752
rect 12099 38696 12167 38752
rect 12223 38696 12291 38752
rect 12347 38696 12415 38752
rect 12471 38696 12481 38752
rect 10669 38628 12481 38696
rect 10669 38572 10679 38628
rect 10735 38572 10803 38628
rect 10859 38572 10927 38628
rect 10983 38572 11051 38628
rect 11107 38572 11175 38628
rect 11231 38572 11299 38628
rect 11355 38572 11423 38628
rect 11479 38572 11547 38628
rect 11603 38572 11671 38628
rect 11727 38572 11795 38628
rect 11851 38572 11919 38628
rect 11975 38572 12043 38628
rect 12099 38572 12167 38628
rect 12223 38572 12291 38628
rect 12347 38572 12415 38628
rect 12471 38572 12481 38628
rect 10669 38504 12481 38572
rect 10669 38448 10679 38504
rect 10735 38448 10803 38504
rect 10859 38448 10927 38504
rect 10983 38448 11051 38504
rect 11107 38448 11175 38504
rect 11231 38448 11299 38504
rect 11355 38448 11423 38504
rect 11479 38448 11547 38504
rect 11603 38448 11671 38504
rect 11727 38448 11795 38504
rect 11851 38448 11919 38504
rect 11975 38448 12043 38504
rect 12099 38448 12167 38504
rect 12223 38448 12291 38504
rect 12347 38448 12415 38504
rect 12471 38448 12481 38504
rect 10669 38438 12481 38448
rect 2517 37000 2593 37010
rect 2517 36944 2527 37000
rect 2583 36944 2593 37000
rect 2517 36876 2593 36944
rect 2517 36820 2527 36876
rect 2583 36820 2593 36876
rect 2517 36752 2593 36820
rect 2517 36696 2527 36752
rect 2583 36696 2593 36752
rect 2517 36628 2593 36696
rect 2517 36572 2527 36628
rect 2583 36572 2593 36628
rect 2517 36504 2593 36572
rect 2517 36448 2527 36504
rect 2583 36448 2593 36504
rect 2517 36380 2593 36448
rect 2517 36324 2527 36380
rect 2583 36324 2593 36380
rect 2517 36256 2593 36324
rect 2517 36200 2527 36256
rect 2583 36200 2593 36256
rect 2517 36132 2593 36200
rect 2517 36076 2527 36132
rect 2583 36076 2593 36132
rect 2517 36008 2593 36076
rect 2517 35952 2527 36008
rect 2583 35952 2593 36008
rect 2517 35884 2593 35952
rect 2517 35828 2527 35884
rect 2583 35828 2593 35884
rect 2517 35760 2593 35828
rect 2517 35704 2527 35760
rect 2583 35704 2593 35760
rect 2517 35636 2593 35704
rect 2517 35580 2527 35636
rect 2583 35580 2593 35636
rect 2517 35512 2593 35580
rect 2517 35456 2527 35512
rect 2583 35456 2593 35512
rect 2517 35388 2593 35456
rect 2517 35332 2527 35388
rect 2583 35332 2593 35388
rect 2517 35264 2593 35332
rect 2517 35208 2527 35264
rect 2583 35208 2593 35264
rect 2517 35140 2593 35208
rect 2517 35084 2527 35140
rect 2583 35084 2593 35140
rect 2517 35016 2593 35084
rect 2517 34960 2527 35016
rect 2583 34960 2593 35016
rect 2517 34892 2593 34960
rect 2517 34836 2527 34892
rect 2583 34836 2593 34892
rect 2517 34768 2593 34836
rect 2517 34712 2527 34768
rect 2583 34712 2593 34768
rect 2517 34644 2593 34712
rect 2517 34588 2527 34644
rect 2583 34588 2593 34644
rect 2517 34520 2593 34588
rect 2517 34464 2527 34520
rect 2583 34464 2593 34520
rect 2517 34396 2593 34464
rect 2517 34340 2527 34396
rect 2583 34340 2593 34396
rect 2517 34272 2593 34340
rect 2517 34216 2527 34272
rect 2583 34216 2593 34272
rect 2517 34148 2593 34216
rect 2517 34092 2527 34148
rect 2583 34092 2593 34148
rect 2517 34024 2593 34092
rect 2517 33968 2527 34024
rect 2583 33968 2593 34024
rect 2517 33900 2593 33968
rect 2517 33844 2527 33900
rect 2583 33844 2593 33900
rect 2517 33776 2593 33844
rect 1145 33766 1221 33776
rect 1145 33710 1155 33766
rect 1211 33710 1221 33766
rect 1145 33642 1221 33710
rect 2517 33720 2527 33776
rect 2583 33720 2593 33776
rect 2517 33652 2593 33720
rect 1145 33586 1155 33642
rect 1211 33586 1221 33642
rect 1145 33518 1221 33586
rect 1145 33462 1155 33518
rect 1211 33462 1221 33518
rect 1145 33394 1221 33462
rect 1145 33338 1155 33394
rect 1211 33338 1221 33394
rect 1145 33270 1221 33338
rect 1145 33214 1155 33270
rect 1211 33214 1221 33270
rect 1145 33146 1221 33214
rect 1145 33090 1155 33146
rect 1211 33090 1221 33146
rect 1145 33022 1221 33090
rect 1145 32966 1155 33022
rect 1211 32966 1221 33022
rect 1145 32898 1221 32966
rect 1145 32842 1155 32898
rect 1211 32842 1221 32898
rect 1145 32774 1221 32842
rect 1145 32718 1155 32774
rect 1211 32718 1221 32774
rect 1145 32650 1221 32718
rect 1145 32594 1155 32650
rect 1211 32594 1221 32650
rect 1145 32526 1221 32594
rect 1145 32470 1155 32526
rect 1211 32470 1221 32526
rect 1145 32402 1221 32470
rect 1145 32346 1155 32402
rect 1211 32346 1221 32402
rect 1145 32278 1221 32346
rect 1145 32222 1155 32278
rect 1211 32222 1221 32278
rect 1145 32154 1221 32222
rect 1145 32098 1155 32154
rect 1211 32098 1221 32154
rect 1145 32030 1221 32098
rect 1145 31974 1155 32030
rect 1211 31974 1221 32030
rect 1145 31906 1221 31974
rect 1145 31850 1155 31906
rect 1211 31850 1221 31906
rect 1145 31782 1221 31850
rect 1145 31726 1155 31782
rect 1211 31726 1221 31782
rect 1145 31658 1221 31726
rect 1145 31602 1155 31658
rect 1211 31602 1221 31658
rect 1145 31534 1221 31602
rect 1145 31478 1155 31534
rect 1211 31478 1221 31534
rect 1145 31410 1221 31478
rect 1145 31354 1155 31410
rect 1211 31354 1221 31410
rect 1145 31286 1221 31354
rect 1145 31230 1155 31286
rect 1211 31230 1221 31286
rect 1145 31162 1221 31230
rect 1145 31106 1155 31162
rect 1211 31106 1221 31162
rect 1145 31038 1221 31106
rect 1145 30982 1155 31038
rect 1211 30982 1221 31038
rect 1145 30914 1221 30982
rect 1145 30858 1155 30914
rect 1211 30858 1221 30914
rect 1145 30790 1221 30858
rect 1145 30734 1155 30790
rect 1211 30734 1221 30790
rect 1145 30666 1221 30734
rect 1145 30610 1155 30666
rect 1211 30610 1221 30666
rect 1145 30542 1221 30610
rect 1145 30486 1155 30542
rect 1211 30486 1221 30542
rect 1145 30418 1221 30486
rect 1145 30362 1155 30418
rect 1211 30362 1221 30418
rect 1145 30294 1221 30362
rect 1145 30238 1155 30294
rect 1211 30238 1221 30294
rect 1145 30170 1221 30238
rect 1145 30114 1155 30170
rect 1211 30114 1221 30170
rect 1145 30046 1221 30114
rect 1145 29990 1155 30046
rect 1211 29990 1221 30046
rect 1145 29922 1221 29990
rect 1145 29866 1155 29922
rect 1211 29866 1221 29922
rect 1145 29798 1221 29866
rect 1145 29742 1155 29798
rect 1211 29742 1221 29798
rect 1145 29732 1221 29742
rect 1269 33642 1345 33652
rect 1269 33586 1279 33642
rect 1335 33586 1345 33642
rect 1269 33518 1345 33586
rect 2517 33596 2527 33652
rect 2583 33596 2593 33652
rect 2517 33528 2593 33596
rect 1269 33462 1279 33518
rect 1335 33462 1345 33518
rect 1269 33394 1345 33462
rect 1269 33338 1279 33394
rect 1335 33338 1345 33394
rect 1269 33270 1345 33338
rect 1269 33214 1279 33270
rect 1335 33214 1345 33270
rect 1269 33146 1345 33214
rect 1269 33090 1279 33146
rect 1335 33090 1345 33146
rect 1269 33022 1345 33090
rect 1269 32966 1279 33022
rect 1335 32966 1345 33022
rect 1269 32898 1345 32966
rect 1269 32842 1279 32898
rect 1335 32842 1345 32898
rect 1269 32774 1345 32842
rect 1269 32718 1279 32774
rect 1335 32718 1345 32774
rect 1269 32650 1345 32718
rect 1269 32594 1279 32650
rect 1335 32594 1345 32650
rect 1269 32526 1345 32594
rect 1269 32470 1279 32526
rect 1335 32470 1345 32526
rect 1269 32402 1345 32470
rect 1269 32346 1279 32402
rect 1335 32346 1345 32402
rect 1269 32278 1345 32346
rect 1269 32222 1279 32278
rect 1335 32222 1345 32278
rect 1269 32154 1345 32222
rect 1269 32098 1279 32154
rect 1335 32098 1345 32154
rect 1269 32030 1345 32098
rect 1269 31974 1279 32030
rect 1335 31974 1345 32030
rect 1269 31906 1345 31974
rect 1269 31850 1279 31906
rect 1335 31850 1345 31906
rect 1269 31782 1345 31850
rect 1269 31726 1279 31782
rect 1335 31726 1345 31782
rect 1269 31658 1345 31726
rect 1269 31602 1279 31658
rect 1335 31602 1345 31658
rect 1269 31534 1345 31602
rect 1269 31478 1279 31534
rect 1335 31478 1345 31534
rect 1269 31410 1345 31478
rect 1269 31354 1279 31410
rect 1335 31354 1345 31410
rect 1269 31286 1345 31354
rect 1269 31230 1279 31286
rect 1335 31230 1345 31286
rect 1269 31162 1345 31230
rect 1269 31106 1279 31162
rect 1335 31106 1345 31162
rect 1269 31038 1345 31106
rect 1269 30982 1279 31038
rect 1335 30982 1345 31038
rect 1269 30914 1345 30982
rect 1269 30858 1279 30914
rect 1335 30858 1345 30914
rect 1269 30790 1345 30858
rect 1269 30734 1279 30790
rect 1335 30734 1345 30790
rect 1269 30666 1345 30734
rect 1269 30610 1279 30666
rect 1335 30610 1345 30666
rect 1269 30542 1345 30610
rect 1269 30486 1279 30542
rect 1335 30486 1345 30542
rect 1269 30418 1345 30486
rect 1269 30362 1279 30418
rect 1335 30362 1345 30418
rect 1269 30294 1345 30362
rect 1269 30238 1279 30294
rect 1335 30238 1345 30294
rect 1269 30170 1345 30238
rect 1269 30114 1279 30170
rect 1335 30114 1345 30170
rect 1269 30046 1345 30114
rect 1269 29990 1279 30046
rect 1335 29990 1345 30046
rect 1269 29922 1345 29990
rect 1269 29866 1279 29922
rect 1335 29866 1345 29922
rect 1269 29798 1345 29866
rect 1269 29742 1279 29798
rect 1335 29742 1345 29798
rect 1269 29674 1345 29742
rect 1269 29618 1279 29674
rect 1335 29618 1345 29674
rect 1269 29608 1345 29618
rect 1393 33518 1469 33528
rect 1393 33462 1403 33518
rect 1459 33462 1469 33518
rect 1393 33394 1469 33462
rect 2517 33472 2527 33528
rect 2583 33472 2593 33528
rect 2517 33404 2593 33472
rect 1393 33338 1403 33394
rect 1459 33338 1469 33394
rect 1393 33270 1469 33338
rect 1393 33214 1403 33270
rect 1459 33214 1469 33270
rect 1393 33146 1469 33214
rect 1393 33090 1403 33146
rect 1459 33090 1469 33146
rect 1393 33022 1469 33090
rect 1393 32966 1403 33022
rect 1459 32966 1469 33022
rect 1393 32898 1469 32966
rect 1393 32842 1403 32898
rect 1459 32842 1469 32898
rect 1393 32774 1469 32842
rect 1393 32718 1403 32774
rect 1459 32718 1469 32774
rect 1393 32650 1469 32718
rect 1393 32594 1403 32650
rect 1459 32594 1469 32650
rect 1393 32526 1469 32594
rect 1393 32470 1403 32526
rect 1459 32470 1469 32526
rect 1393 32402 1469 32470
rect 1393 32346 1403 32402
rect 1459 32346 1469 32402
rect 1393 32278 1469 32346
rect 1393 32222 1403 32278
rect 1459 32222 1469 32278
rect 1393 32154 1469 32222
rect 1393 32098 1403 32154
rect 1459 32098 1469 32154
rect 1393 32030 1469 32098
rect 1393 31974 1403 32030
rect 1459 31974 1469 32030
rect 1393 31906 1469 31974
rect 1393 31850 1403 31906
rect 1459 31850 1469 31906
rect 1393 31782 1469 31850
rect 1393 31726 1403 31782
rect 1459 31726 1469 31782
rect 1393 31658 1469 31726
rect 1393 31602 1403 31658
rect 1459 31602 1469 31658
rect 1393 31534 1469 31602
rect 1393 31478 1403 31534
rect 1459 31478 1469 31534
rect 1393 31410 1469 31478
rect 1393 31354 1403 31410
rect 1459 31354 1469 31410
rect 1393 31286 1469 31354
rect 1393 31230 1403 31286
rect 1459 31230 1469 31286
rect 1393 31162 1469 31230
rect 1393 31106 1403 31162
rect 1459 31106 1469 31162
rect 1393 31038 1469 31106
rect 1393 30982 1403 31038
rect 1459 30982 1469 31038
rect 1393 30914 1469 30982
rect 1393 30858 1403 30914
rect 1459 30858 1469 30914
rect 1393 30790 1469 30858
rect 1393 30734 1403 30790
rect 1459 30734 1469 30790
rect 1393 30666 1469 30734
rect 1393 30610 1403 30666
rect 1459 30610 1469 30666
rect 1393 30542 1469 30610
rect 1393 30486 1403 30542
rect 1459 30486 1469 30542
rect 1393 30418 1469 30486
rect 1393 30362 1403 30418
rect 1459 30362 1469 30418
rect 1393 30294 1469 30362
rect 1393 30238 1403 30294
rect 1459 30238 1469 30294
rect 1393 30170 1469 30238
rect 1393 30114 1403 30170
rect 1459 30114 1469 30170
rect 1393 30046 1469 30114
rect 1393 29990 1403 30046
rect 1459 29990 1469 30046
rect 1393 29922 1469 29990
rect 1393 29866 1403 29922
rect 1459 29866 1469 29922
rect 1393 29798 1469 29866
rect 1393 29742 1403 29798
rect 1459 29742 1469 29798
rect 1393 29674 1469 29742
rect 1393 29618 1403 29674
rect 1459 29618 1469 29674
rect 1393 29550 1469 29618
rect 1393 29494 1403 29550
rect 1459 29494 1469 29550
rect 1393 29484 1469 29494
rect 1517 33394 1593 33404
rect 1517 33338 1527 33394
rect 1583 33338 1593 33394
rect 1517 33270 1593 33338
rect 2517 33348 2527 33404
rect 2583 33348 2593 33404
rect 2517 33280 2593 33348
rect 1517 33214 1527 33270
rect 1583 33214 1593 33270
rect 1517 33146 1593 33214
rect 1517 33090 1527 33146
rect 1583 33090 1593 33146
rect 1517 33022 1593 33090
rect 1517 32966 1527 33022
rect 1583 32966 1593 33022
rect 1517 32898 1593 32966
rect 1517 32842 1527 32898
rect 1583 32842 1593 32898
rect 1517 32774 1593 32842
rect 1517 32718 1527 32774
rect 1583 32718 1593 32774
rect 1517 32650 1593 32718
rect 1517 32594 1527 32650
rect 1583 32594 1593 32650
rect 1517 32526 1593 32594
rect 1517 32470 1527 32526
rect 1583 32470 1593 32526
rect 1517 32402 1593 32470
rect 1517 32346 1527 32402
rect 1583 32346 1593 32402
rect 1517 32278 1593 32346
rect 1517 32222 1527 32278
rect 1583 32222 1593 32278
rect 1517 32154 1593 32222
rect 1517 32098 1527 32154
rect 1583 32098 1593 32154
rect 1517 32030 1593 32098
rect 1517 31974 1527 32030
rect 1583 31974 1593 32030
rect 1517 31906 1593 31974
rect 1517 31850 1527 31906
rect 1583 31850 1593 31906
rect 1517 31782 1593 31850
rect 1517 31726 1527 31782
rect 1583 31726 1593 31782
rect 1517 31658 1593 31726
rect 1517 31602 1527 31658
rect 1583 31602 1593 31658
rect 1517 31534 1593 31602
rect 1517 31478 1527 31534
rect 1583 31478 1593 31534
rect 1517 31410 1593 31478
rect 1517 31354 1527 31410
rect 1583 31354 1593 31410
rect 1517 31286 1593 31354
rect 1517 31230 1527 31286
rect 1583 31230 1593 31286
rect 1517 31162 1593 31230
rect 1517 31106 1527 31162
rect 1583 31106 1593 31162
rect 1517 31038 1593 31106
rect 1517 30982 1527 31038
rect 1583 30982 1593 31038
rect 1517 30914 1593 30982
rect 1517 30858 1527 30914
rect 1583 30858 1593 30914
rect 1517 30790 1593 30858
rect 1517 30734 1527 30790
rect 1583 30734 1593 30790
rect 1517 30666 1593 30734
rect 1517 30610 1527 30666
rect 1583 30610 1593 30666
rect 1517 30542 1593 30610
rect 1517 30486 1527 30542
rect 1583 30486 1593 30542
rect 1517 30418 1593 30486
rect 1517 30362 1527 30418
rect 1583 30362 1593 30418
rect 1517 30294 1593 30362
rect 1517 30238 1527 30294
rect 1583 30238 1593 30294
rect 1517 30170 1593 30238
rect 1517 30114 1527 30170
rect 1583 30114 1593 30170
rect 1517 30046 1593 30114
rect 1517 29990 1527 30046
rect 1583 29990 1593 30046
rect 1517 29922 1593 29990
rect 1517 29866 1527 29922
rect 1583 29866 1593 29922
rect 1517 29798 1593 29866
rect 1517 29742 1527 29798
rect 1583 29742 1593 29798
rect 1517 29674 1593 29742
rect 1517 29618 1527 29674
rect 1583 29618 1593 29674
rect 1517 29550 1593 29618
rect 1517 29494 1527 29550
rect 1583 29494 1593 29550
rect 1517 29426 1593 29494
rect 1517 29370 1527 29426
rect 1583 29370 1593 29426
rect 1517 29360 1593 29370
rect 1641 33270 1717 33280
rect 1641 33214 1651 33270
rect 1707 33214 1717 33270
rect 1641 33146 1717 33214
rect 2517 33224 2527 33280
rect 2583 33224 2593 33280
rect 2517 33156 2593 33224
rect 1641 33090 1651 33146
rect 1707 33090 1717 33146
rect 1641 33022 1717 33090
rect 1641 32966 1651 33022
rect 1707 32966 1717 33022
rect 1641 32898 1717 32966
rect 1641 32842 1651 32898
rect 1707 32842 1717 32898
rect 1641 32774 1717 32842
rect 1641 32718 1651 32774
rect 1707 32718 1717 32774
rect 1641 32650 1717 32718
rect 1641 32594 1651 32650
rect 1707 32594 1717 32650
rect 1641 32526 1717 32594
rect 1641 32470 1651 32526
rect 1707 32470 1717 32526
rect 1641 32402 1717 32470
rect 1641 32346 1651 32402
rect 1707 32346 1717 32402
rect 1641 32278 1717 32346
rect 1641 32222 1651 32278
rect 1707 32222 1717 32278
rect 1641 32154 1717 32222
rect 1641 32098 1651 32154
rect 1707 32098 1717 32154
rect 1641 32030 1717 32098
rect 1641 31974 1651 32030
rect 1707 31974 1717 32030
rect 1641 31906 1717 31974
rect 1641 31850 1651 31906
rect 1707 31850 1717 31906
rect 1641 31782 1717 31850
rect 1641 31726 1651 31782
rect 1707 31726 1717 31782
rect 1641 31658 1717 31726
rect 1641 31602 1651 31658
rect 1707 31602 1717 31658
rect 1641 31534 1717 31602
rect 1641 31478 1651 31534
rect 1707 31478 1717 31534
rect 1641 31410 1717 31478
rect 1641 31354 1651 31410
rect 1707 31354 1717 31410
rect 1641 31286 1717 31354
rect 1641 31230 1651 31286
rect 1707 31230 1717 31286
rect 1641 31162 1717 31230
rect 1641 31106 1651 31162
rect 1707 31106 1717 31162
rect 1641 31038 1717 31106
rect 1641 30982 1651 31038
rect 1707 30982 1717 31038
rect 1641 30914 1717 30982
rect 1641 30858 1651 30914
rect 1707 30858 1717 30914
rect 1641 30790 1717 30858
rect 1641 30734 1651 30790
rect 1707 30734 1717 30790
rect 1641 30666 1717 30734
rect 1641 30610 1651 30666
rect 1707 30610 1717 30666
rect 1641 30542 1717 30610
rect 1641 30486 1651 30542
rect 1707 30486 1717 30542
rect 1641 30418 1717 30486
rect 1641 30362 1651 30418
rect 1707 30362 1717 30418
rect 1641 30294 1717 30362
rect 1641 30238 1651 30294
rect 1707 30238 1717 30294
rect 1641 30170 1717 30238
rect 1641 30114 1651 30170
rect 1707 30114 1717 30170
rect 1641 30046 1717 30114
rect 1641 29990 1651 30046
rect 1707 29990 1717 30046
rect 1641 29922 1717 29990
rect 1641 29866 1651 29922
rect 1707 29866 1717 29922
rect 1641 29798 1717 29866
rect 1641 29742 1651 29798
rect 1707 29742 1717 29798
rect 1641 29674 1717 29742
rect 1641 29618 1651 29674
rect 1707 29618 1717 29674
rect 1641 29550 1717 29618
rect 1641 29494 1651 29550
rect 1707 29494 1717 29550
rect 1641 29426 1717 29494
rect 1641 29370 1651 29426
rect 1707 29370 1717 29426
rect 1117 29307 1193 29317
rect 1117 29251 1127 29307
rect 1183 29251 1193 29307
rect 1117 29183 1193 29251
rect 1641 29302 1717 29370
rect 1641 29246 1651 29302
rect 1707 29246 1717 29302
rect 1641 29236 1717 29246
rect 1765 33146 1841 33156
rect 1765 33090 1775 33146
rect 1831 33090 1841 33146
rect 1765 33022 1841 33090
rect 2517 33100 2527 33156
rect 2583 33100 2593 33156
rect 2517 33032 2593 33100
rect 1765 32966 1775 33022
rect 1831 32966 1841 33022
rect 1765 32898 1841 32966
rect 1765 32842 1775 32898
rect 1831 32842 1841 32898
rect 1765 32774 1841 32842
rect 1765 32718 1775 32774
rect 1831 32718 1841 32774
rect 1765 32650 1841 32718
rect 1765 32594 1775 32650
rect 1831 32594 1841 32650
rect 1765 32526 1841 32594
rect 1765 32470 1775 32526
rect 1831 32470 1841 32526
rect 1765 32402 1841 32470
rect 1765 32346 1775 32402
rect 1831 32346 1841 32402
rect 1765 32278 1841 32346
rect 1765 32222 1775 32278
rect 1831 32222 1841 32278
rect 1765 32154 1841 32222
rect 1765 32098 1775 32154
rect 1831 32098 1841 32154
rect 1765 32030 1841 32098
rect 1765 31974 1775 32030
rect 1831 31974 1841 32030
rect 1765 31906 1841 31974
rect 1765 31850 1775 31906
rect 1831 31850 1841 31906
rect 1765 31782 1841 31850
rect 1765 31726 1775 31782
rect 1831 31726 1841 31782
rect 1765 31658 1841 31726
rect 1765 31602 1775 31658
rect 1831 31602 1841 31658
rect 1765 31534 1841 31602
rect 1765 31478 1775 31534
rect 1831 31478 1841 31534
rect 1765 31410 1841 31478
rect 1765 31354 1775 31410
rect 1831 31354 1841 31410
rect 1765 31286 1841 31354
rect 1765 31230 1775 31286
rect 1831 31230 1841 31286
rect 1765 31162 1841 31230
rect 1765 31106 1775 31162
rect 1831 31106 1841 31162
rect 1765 31038 1841 31106
rect 1765 30982 1775 31038
rect 1831 30982 1841 31038
rect 1765 30914 1841 30982
rect 1765 30858 1775 30914
rect 1831 30858 1841 30914
rect 1765 30790 1841 30858
rect 1765 30734 1775 30790
rect 1831 30734 1841 30790
rect 1765 30666 1841 30734
rect 1765 30610 1775 30666
rect 1831 30610 1841 30666
rect 1765 30542 1841 30610
rect 1765 30486 1775 30542
rect 1831 30486 1841 30542
rect 1765 30418 1841 30486
rect 1765 30362 1775 30418
rect 1831 30362 1841 30418
rect 1765 30294 1841 30362
rect 1765 30238 1775 30294
rect 1831 30238 1841 30294
rect 1765 30170 1841 30238
rect 1765 30114 1775 30170
rect 1831 30114 1841 30170
rect 1765 30046 1841 30114
rect 1765 29990 1775 30046
rect 1831 29990 1841 30046
rect 1765 29922 1841 29990
rect 1765 29866 1775 29922
rect 1831 29866 1841 29922
rect 1765 29798 1841 29866
rect 1765 29742 1775 29798
rect 1831 29742 1841 29798
rect 1765 29674 1841 29742
rect 1765 29618 1775 29674
rect 1831 29618 1841 29674
rect 1765 29550 1841 29618
rect 1765 29494 1775 29550
rect 1831 29494 1841 29550
rect 1765 29426 1841 29494
rect 1765 29370 1775 29426
rect 1831 29370 1841 29426
rect 1765 29302 1841 29370
rect 1765 29246 1775 29302
rect 1831 29246 1841 29302
rect 1117 29127 1127 29183
rect 1183 29127 1193 29183
rect 1117 29059 1193 29127
rect 1117 29003 1127 29059
rect 1183 29003 1193 29059
rect 1117 28935 1193 29003
rect 1117 28879 1127 28935
rect 1183 28879 1193 28935
rect 1117 28811 1193 28879
rect 1117 28755 1127 28811
rect 1183 28755 1193 28811
rect 1117 28687 1193 28755
rect 1117 28631 1127 28687
rect 1183 28631 1193 28687
rect 1117 28563 1193 28631
rect 1117 28507 1127 28563
rect 1183 28507 1193 28563
rect 1117 28439 1193 28507
rect 1117 28383 1127 28439
rect 1183 28383 1193 28439
rect 1117 28315 1193 28383
rect 1117 28259 1127 28315
rect 1183 28259 1193 28315
rect 1117 28191 1193 28259
rect 1117 28135 1127 28191
rect 1183 28135 1193 28191
rect 1117 28067 1193 28135
rect 1117 28011 1127 28067
rect 1183 28011 1193 28067
rect 1117 27943 1193 28011
rect 1117 27887 1127 27943
rect 1183 27887 1193 27943
rect 1117 27819 1193 27887
rect 1117 27763 1127 27819
rect 1183 27763 1193 27819
rect 1117 27695 1193 27763
rect 1117 27639 1127 27695
rect 1183 27639 1193 27695
rect 1117 27571 1193 27639
rect 1117 27515 1127 27571
rect 1183 27515 1193 27571
rect 1117 27505 1193 27515
rect 1241 29183 1317 29193
rect 1241 29127 1251 29183
rect 1307 29127 1317 29183
rect 1241 29059 1317 29127
rect 1765 29178 1841 29246
rect 1765 29122 1775 29178
rect 1831 29122 1841 29178
rect 1765 29112 1841 29122
rect 1889 33022 1965 33032
rect 1889 32966 1899 33022
rect 1955 32966 1965 33022
rect 2517 32976 2527 33032
rect 2583 32976 2593 33032
rect 2517 32966 2593 32976
rect 2641 36876 2717 36886
rect 2641 36820 2651 36876
rect 2707 36820 2717 36876
rect 2641 36752 2717 36820
rect 2641 36696 2651 36752
rect 2707 36696 2717 36752
rect 2641 36628 2717 36696
rect 2641 36572 2651 36628
rect 2707 36572 2717 36628
rect 2641 36504 2717 36572
rect 2641 36448 2651 36504
rect 2707 36448 2717 36504
rect 2641 36380 2717 36448
rect 2641 36324 2651 36380
rect 2707 36324 2717 36380
rect 2641 36256 2717 36324
rect 2641 36200 2651 36256
rect 2707 36200 2717 36256
rect 2641 36132 2717 36200
rect 2641 36076 2651 36132
rect 2707 36076 2717 36132
rect 2641 36008 2717 36076
rect 2641 35952 2651 36008
rect 2707 35952 2717 36008
rect 2641 35884 2717 35952
rect 2641 35828 2651 35884
rect 2707 35828 2717 35884
rect 2641 35760 2717 35828
rect 2641 35704 2651 35760
rect 2707 35704 2717 35760
rect 2641 35636 2717 35704
rect 2641 35580 2651 35636
rect 2707 35580 2717 35636
rect 2641 35512 2717 35580
rect 2641 35456 2651 35512
rect 2707 35456 2717 35512
rect 2641 35388 2717 35456
rect 2641 35332 2651 35388
rect 2707 35332 2717 35388
rect 2641 35264 2717 35332
rect 2641 35208 2651 35264
rect 2707 35208 2717 35264
rect 2641 35140 2717 35208
rect 2641 35084 2651 35140
rect 2707 35084 2717 35140
rect 2641 35016 2717 35084
rect 2641 34960 2651 35016
rect 2707 34960 2717 35016
rect 2641 34892 2717 34960
rect 2641 34836 2651 34892
rect 2707 34836 2717 34892
rect 2641 34768 2717 34836
rect 2641 34712 2651 34768
rect 2707 34712 2717 34768
rect 2641 34644 2717 34712
rect 2641 34588 2651 34644
rect 2707 34588 2717 34644
rect 2641 34520 2717 34588
rect 2641 34464 2651 34520
rect 2707 34464 2717 34520
rect 2641 34396 2717 34464
rect 2641 34340 2651 34396
rect 2707 34340 2717 34396
rect 2641 34272 2717 34340
rect 2641 34216 2651 34272
rect 2707 34216 2717 34272
rect 2641 34148 2717 34216
rect 2641 34092 2651 34148
rect 2707 34092 2717 34148
rect 2641 34024 2717 34092
rect 2641 33968 2651 34024
rect 2707 33968 2717 34024
rect 2641 33900 2717 33968
rect 2641 33844 2651 33900
rect 2707 33844 2717 33900
rect 2641 33776 2717 33844
rect 2641 33720 2651 33776
rect 2707 33720 2717 33776
rect 2641 33652 2717 33720
rect 2641 33596 2651 33652
rect 2707 33596 2717 33652
rect 2641 33528 2717 33596
rect 2641 33472 2651 33528
rect 2707 33472 2717 33528
rect 2641 33404 2717 33472
rect 2641 33348 2651 33404
rect 2707 33348 2717 33404
rect 2641 33280 2717 33348
rect 2641 33224 2651 33280
rect 2707 33224 2717 33280
rect 2641 33156 2717 33224
rect 2641 33100 2651 33156
rect 2707 33100 2717 33156
rect 2641 33032 2717 33100
rect 2641 32976 2651 33032
rect 2707 32976 2717 33032
rect 1889 32898 1965 32966
rect 2641 32908 2717 32976
rect 1889 32842 1899 32898
rect 1955 32842 1965 32898
rect 1889 32774 1965 32842
rect 1889 32718 1899 32774
rect 1955 32718 1965 32774
rect 1889 32650 1965 32718
rect 1889 32594 1899 32650
rect 1955 32594 1965 32650
rect 1889 32526 1965 32594
rect 1889 32470 1899 32526
rect 1955 32470 1965 32526
rect 1889 32402 1965 32470
rect 1889 32346 1899 32402
rect 1955 32346 1965 32402
rect 1889 32278 1965 32346
rect 1889 32222 1899 32278
rect 1955 32222 1965 32278
rect 1889 32154 1965 32222
rect 1889 32098 1899 32154
rect 1955 32098 1965 32154
rect 1889 32030 1965 32098
rect 1889 31974 1899 32030
rect 1955 31974 1965 32030
rect 1889 31906 1965 31974
rect 1889 31850 1899 31906
rect 1955 31850 1965 31906
rect 1889 31782 1965 31850
rect 1889 31726 1899 31782
rect 1955 31726 1965 31782
rect 1889 31658 1965 31726
rect 1889 31602 1899 31658
rect 1955 31602 1965 31658
rect 1889 31534 1965 31602
rect 1889 31478 1899 31534
rect 1955 31478 1965 31534
rect 1889 31410 1965 31478
rect 1889 31354 1899 31410
rect 1955 31354 1965 31410
rect 1889 31286 1965 31354
rect 1889 31230 1899 31286
rect 1955 31230 1965 31286
rect 1889 31162 1965 31230
rect 1889 31106 1899 31162
rect 1955 31106 1965 31162
rect 1889 31038 1965 31106
rect 1889 30982 1899 31038
rect 1955 30982 1965 31038
rect 1889 30914 1965 30982
rect 1889 30858 1899 30914
rect 1955 30858 1965 30914
rect 1889 30790 1965 30858
rect 1889 30734 1899 30790
rect 1955 30734 1965 30790
rect 1889 30666 1965 30734
rect 1889 30610 1899 30666
rect 1955 30610 1965 30666
rect 1889 30542 1965 30610
rect 1889 30486 1899 30542
rect 1955 30486 1965 30542
rect 1889 30418 1965 30486
rect 1889 30362 1899 30418
rect 1955 30362 1965 30418
rect 1889 30294 1965 30362
rect 1889 30238 1899 30294
rect 1955 30238 1965 30294
rect 1889 30170 1965 30238
rect 1889 30114 1899 30170
rect 1955 30114 1965 30170
rect 1889 30046 1965 30114
rect 1889 29990 1899 30046
rect 1955 29990 1965 30046
rect 1889 29922 1965 29990
rect 1889 29866 1899 29922
rect 1955 29866 1965 29922
rect 1889 29798 1965 29866
rect 1889 29742 1899 29798
rect 1955 29742 1965 29798
rect 1889 29674 1965 29742
rect 1889 29618 1899 29674
rect 1955 29618 1965 29674
rect 1889 29550 1965 29618
rect 1889 29494 1899 29550
rect 1955 29494 1965 29550
rect 1889 29426 1965 29494
rect 1889 29370 1899 29426
rect 1955 29370 1965 29426
rect 1889 29302 1965 29370
rect 1889 29246 1899 29302
rect 1955 29246 1965 29302
rect 1889 29178 1965 29246
rect 1889 29122 1899 29178
rect 1955 29122 1965 29178
rect 1241 29003 1251 29059
rect 1307 29003 1317 29059
rect 1241 28935 1317 29003
rect 1241 28879 1251 28935
rect 1307 28879 1317 28935
rect 1241 28811 1317 28879
rect 1241 28755 1251 28811
rect 1307 28755 1317 28811
rect 1241 28687 1317 28755
rect 1241 28631 1251 28687
rect 1307 28631 1317 28687
rect 1241 28563 1317 28631
rect 1241 28507 1251 28563
rect 1307 28507 1317 28563
rect 1241 28439 1317 28507
rect 1241 28383 1251 28439
rect 1307 28383 1317 28439
rect 1241 28315 1317 28383
rect 1241 28259 1251 28315
rect 1307 28259 1317 28315
rect 1241 28191 1317 28259
rect 1241 28135 1251 28191
rect 1307 28135 1317 28191
rect 1241 28067 1317 28135
rect 1241 28011 1251 28067
rect 1307 28011 1317 28067
rect 1241 27943 1317 28011
rect 1241 27887 1251 27943
rect 1307 27887 1317 27943
rect 1241 27819 1317 27887
rect 1241 27763 1251 27819
rect 1307 27763 1317 27819
rect 1241 27695 1317 27763
rect 1241 27639 1251 27695
rect 1307 27639 1317 27695
rect 1241 27571 1317 27639
rect 1241 27515 1251 27571
rect 1307 27515 1317 27571
rect 1241 27447 1317 27515
rect 1241 27391 1251 27447
rect 1307 27391 1317 27447
rect 1241 27381 1317 27391
rect 1365 29059 1441 29069
rect 1365 29003 1375 29059
rect 1431 29003 1441 29059
rect 1365 28935 1441 29003
rect 1889 29054 1965 29122
rect 1889 28998 1899 29054
rect 1955 28998 1965 29054
rect 1889 28988 1965 28998
rect 2013 32898 2089 32908
rect 2013 32842 2023 32898
rect 2079 32842 2089 32898
rect 2641 32852 2651 32908
rect 2707 32852 2717 32908
rect 2641 32842 2717 32852
rect 2765 36752 2841 36762
rect 2765 36696 2775 36752
rect 2831 36696 2841 36752
rect 2765 36628 2841 36696
rect 2765 36572 2775 36628
rect 2831 36572 2841 36628
rect 2765 36504 2841 36572
rect 2765 36448 2775 36504
rect 2831 36448 2841 36504
rect 2765 36380 2841 36448
rect 2765 36324 2775 36380
rect 2831 36324 2841 36380
rect 2765 36256 2841 36324
rect 2765 36200 2775 36256
rect 2831 36200 2841 36256
rect 2765 36132 2841 36200
rect 2765 36076 2775 36132
rect 2831 36076 2841 36132
rect 2765 36008 2841 36076
rect 2765 35952 2775 36008
rect 2831 35952 2841 36008
rect 2765 35884 2841 35952
rect 2765 35828 2775 35884
rect 2831 35828 2841 35884
rect 2765 35760 2841 35828
rect 2765 35704 2775 35760
rect 2831 35704 2841 35760
rect 2765 35636 2841 35704
rect 2765 35580 2775 35636
rect 2831 35580 2841 35636
rect 2765 35512 2841 35580
rect 2765 35456 2775 35512
rect 2831 35456 2841 35512
rect 2765 35388 2841 35456
rect 2765 35332 2775 35388
rect 2831 35332 2841 35388
rect 2765 35264 2841 35332
rect 2765 35208 2775 35264
rect 2831 35208 2841 35264
rect 2765 35140 2841 35208
rect 2765 35084 2775 35140
rect 2831 35084 2841 35140
rect 2765 35016 2841 35084
rect 2765 34960 2775 35016
rect 2831 34960 2841 35016
rect 2765 34892 2841 34960
rect 2765 34836 2775 34892
rect 2831 34836 2841 34892
rect 2765 34768 2841 34836
rect 2765 34712 2775 34768
rect 2831 34712 2841 34768
rect 2765 34644 2841 34712
rect 2765 34588 2775 34644
rect 2831 34588 2841 34644
rect 2765 34520 2841 34588
rect 2765 34464 2775 34520
rect 2831 34464 2841 34520
rect 2765 34396 2841 34464
rect 2765 34340 2775 34396
rect 2831 34340 2841 34396
rect 2765 34272 2841 34340
rect 2765 34216 2775 34272
rect 2831 34216 2841 34272
rect 2765 34148 2841 34216
rect 2765 34092 2775 34148
rect 2831 34092 2841 34148
rect 2765 34024 2841 34092
rect 2765 33968 2775 34024
rect 2831 33968 2841 34024
rect 2765 33900 2841 33968
rect 2765 33844 2775 33900
rect 2831 33844 2841 33900
rect 2765 33776 2841 33844
rect 2765 33720 2775 33776
rect 2831 33720 2841 33776
rect 2765 33652 2841 33720
rect 2765 33596 2775 33652
rect 2831 33596 2841 33652
rect 2765 33528 2841 33596
rect 2765 33472 2775 33528
rect 2831 33472 2841 33528
rect 2765 33404 2841 33472
rect 2765 33348 2775 33404
rect 2831 33348 2841 33404
rect 2765 33280 2841 33348
rect 2765 33224 2775 33280
rect 2831 33224 2841 33280
rect 2765 33156 2841 33224
rect 2765 33100 2775 33156
rect 2831 33100 2841 33156
rect 2765 33032 2841 33100
rect 2765 32976 2775 33032
rect 2831 32976 2841 33032
rect 2765 32908 2841 32976
rect 2765 32852 2775 32908
rect 2831 32852 2841 32908
rect 2013 32774 2089 32842
rect 2013 32718 2023 32774
rect 2079 32718 2089 32774
rect 2765 32784 2841 32852
rect 2765 32728 2775 32784
rect 2831 32728 2841 32784
rect 2765 32718 2841 32728
rect 2889 36628 2965 36638
rect 2889 36572 2899 36628
rect 2955 36572 2965 36628
rect 2889 36504 2965 36572
rect 14757 36572 14833 36582
rect 2889 36448 2899 36504
rect 2955 36448 2965 36504
rect 2889 36380 2965 36448
rect 2889 36324 2899 36380
rect 2955 36324 2965 36380
rect 2889 36256 2965 36324
rect 2889 36200 2899 36256
rect 2955 36200 2965 36256
rect 2889 36132 2965 36200
rect 2889 36076 2899 36132
rect 2955 36076 2965 36132
rect 2889 36008 2965 36076
rect 2889 35952 2899 36008
rect 2955 35952 2965 36008
rect 2889 35884 2965 35952
rect 2889 35828 2899 35884
rect 2955 35828 2965 35884
rect 2889 35760 2965 35828
rect 2889 35704 2899 35760
rect 2955 35704 2965 35760
rect 2889 35636 2965 35704
rect 2889 35580 2899 35636
rect 2955 35580 2965 35636
rect 2889 35512 2965 35580
rect 2889 35456 2899 35512
rect 2955 35456 2965 35512
rect 2889 35388 2965 35456
rect 2889 35332 2899 35388
rect 2955 35332 2965 35388
rect 2889 35264 2965 35332
rect 2889 35208 2899 35264
rect 2955 35208 2965 35264
rect 2889 35140 2965 35208
rect 2889 35084 2899 35140
rect 2955 35084 2965 35140
rect 2889 35016 2965 35084
rect 2889 34960 2899 35016
rect 2955 34960 2965 35016
rect 2889 34892 2965 34960
rect 2889 34836 2899 34892
rect 2955 34836 2965 34892
rect 2889 34768 2965 34836
rect 2889 34712 2899 34768
rect 2955 34712 2965 34768
rect 2889 34644 2965 34712
rect 2889 34588 2899 34644
rect 2955 34588 2965 34644
rect 2889 34520 2965 34588
rect 2889 34464 2899 34520
rect 2955 34464 2965 34520
rect 2889 34396 2965 34464
rect 2889 34340 2899 34396
rect 2955 34340 2965 34396
rect 2889 34272 2965 34340
rect 2889 34216 2899 34272
rect 2955 34216 2965 34272
rect 2889 34148 2965 34216
rect 2889 34092 2899 34148
rect 2955 34092 2965 34148
rect 2889 34024 2965 34092
rect 2889 33968 2899 34024
rect 2955 33968 2965 34024
rect 2889 33900 2965 33968
rect 2889 33844 2899 33900
rect 2955 33844 2965 33900
rect 2889 33776 2965 33844
rect 2889 33720 2899 33776
rect 2955 33720 2965 33776
rect 2889 33652 2965 33720
rect 2889 33596 2899 33652
rect 2955 33596 2965 33652
rect 2889 33528 2965 33596
rect 2889 33472 2899 33528
rect 2955 33472 2965 33528
rect 2889 33404 2965 33472
rect 2889 33348 2899 33404
rect 2955 33348 2965 33404
rect 2889 33280 2965 33348
rect 2889 33224 2899 33280
rect 2955 33224 2965 33280
rect 2889 33156 2965 33224
rect 2889 33100 2899 33156
rect 2955 33100 2965 33156
rect 2889 33032 2965 33100
rect 2889 32976 2899 33032
rect 2955 32976 2965 33032
rect 2889 32908 2965 32976
rect 2889 32852 2899 32908
rect 2955 32852 2965 32908
rect 2889 32784 2965 32852
rect 2889 32728 2899 32784
rect 2955 32728 2965 32784
rect 2013 32650 2089 32718
rect 2013 32594 2023 32650
rect 2079 32594 2089 32650
rect 2889 32660 2965 32728
rect 2889 32604 2899 32660
rect 2955 32604 2965 32660
rect 2889 32594 2965 32604
rect 3013 36504 3089 36514
rect 3013 36448 3023 36504
rect 3079 36448 3089 36504
rect 3013 36380 3089 36448
rect 3013 36324 3023 36380
rect 3079 36324 3089 36380
rect 3013 36256 3089 36324
rect 3013 36200 3023 36256
rect 3079 36200 3089 36256
rect 3013 36132 3089 36200
rect 3013 36076 3023 36132
rect 3079 36076 3089 36132
rect 3013 36008 3089 36076
rect 3013 35952 3023 36008
rect 3079 35952 3089 36008
rect 3013 35884 3089 35952
rect 3013 35828 3023 35884
rect 3079 35828 3089 35884
rect 3013 35760 3089 35828
rect 3013 35704 3023 35760
rect 3079 35704 3089 35760
rect 3013 35636 3089 35704
rect 3013 35580 3023 35636
rect 3079 35580 3089 35636
rect 3013 35512 3089 35580
rect 3013 35456 3023 35512
rect 3079 35456 3089 35512
rect 3013 35388 3089 35456
rect 3013 35332 3023 35388
rect 3079 35332 3089 35388
rect 3013 35264 3089 35332
rect 3013 35208 3023 35264
rect 3079 35208 3089 35264
rect 3013 35140 3089 35208
rect 3013 35084 3023 35140
rect 3079 35084 3089 35140
rect 3013 35016 3089 35084
rect 3013 34960 3023 35016
rect 3079 34960 3089 35016
rect 3013 34892 3089 34960
rect 3013 34836 3023 34892
rect 3079 34836 3089 34892
rect 3013 34768 3089 34836
rect 3013 34712 3023 34768
rect 3079 34712 3089 34768
rect 3013 34644 3089 34712
rect 3013 34588 3023 34644
rect 3079 34588 3089 34644
rect 3013 34520 3089 34588
rect 3013 34464 3023 34520
rect 3079 34464 3089 34520
rect 3013 34396 3089 34464
rect 3013 34340 3023 34396
rect 3079 34340 3089 34396
rect 3013 34272 3089 34340
rect 3013 34216 3023 34272
rect 3079 34216 3089 34272
rect 3013 34148 3089 34216
rect 3013 34092 3023 34148
rect 3079 34092 3089 34148
rect 3013 34024 3089 34092
rect 3013 33968 3023 34024
rect 3079 33968 3089 34024
rect 3013 33900 3089 33968
rect 3013 33844 3023 33900
rect 3079 33844 3089 33900
rect 3013 33776 3089 33844
rect 3013 33720 3023 33776
rect 3079 33720 3089 33776
rect 3013 33652 3089 33720
rect 3013 33596 3023 33652
rect 3079 33596 3089 33652
rect 3013 33528 3089 33596
rect 3013 33472 3023 33528
rect 3079 33472 3089 33528
rect 3013 33404 3089 33472
rect 3013 33348 3023 33404
rect 3079 33348 3089 33404
rect 3013 33280 3089 33348
rect 3013 33224 3023 33280
rect 3079 33224 3089 33280
rect 3013 33156 3089 33224
rect 3013 33100 3023 33156
rect 3079 33100 3089 33156
rect 3013 33032 3089 33100
rect 3013 32976 3023 33032
rect 3079 32976 3089 33032
rect 3013 32908 3089 32976
rect 3013 32852 3023 32908
rect 3079 32852 3089 32908
rect 3013 32784 3089 32852
rect 3013 32728 3023 32784
rect 3079 32728 3089 32784
rect 3013 32660 3089 32728
rect 3013 32604 3023 32660
rect 3079 32604 3089 32660
rect 2013 32526 2089 32594
rect 2013 32470 2023 32526
rect 2079 32470 2089 32526
rect 3013 32536 3089 32604
rect 3013 32480 3023 32536
rect 3079 32480 3089 32536
rect 3013 32470 3089 32480
rect 3137 36380 3213 36390
rect 3137 36324 3147 36380
rect 3203 36324 3213 36380
rect 3137 36256 3213 36324
rect 3137 36200 3147 36256
rect 3203 36200 3213 36256
rect 3137 36132 3213 36200
rect 3137 36076 3147 36132
rect 3203 36076 3213 36132
rect 3137 36008 3213 36076
rect 3137 35952 3147 36008
rect 3203 35952 3213 36008
rect 3137 35884 3213 35952
rect 3137 35828 3147 35884
rect 3203 35828 3213 35884
rect 3137 35760 3213 35828
rect 3137 35704 3147 35760
rect 3203 35704 3213 35760
rect 3137 35636 3213 35704
rect 3137 35580 3147 35636
rect 3203 35580 3213 35636
rect 3137 35512 3213 35580
rect 3137 35456 3147 35512
rect 3203 35456 3213 35512
rect 3137 35388 3213 35456
rect 3137 35332 3147 35388
rect 3203 35332 3213 35388
rect 3137 35264 3213 35332
rect 3137 35208 3147 35264
rect 3203 35208 3213 35264
rect 3137 35140 3213 35208
rect 3137 35084 3147 35140
rect 3203 35084 3213 35140
rect 3137 35016 3213 35084
rect 3137 34960 3147 35016
rect 3203 34960 3213 35016
rect 3137 34892 3213 34960
rect 3137 34836 3147 34892
rect 3203 34836 3213 34892
rect 3137 34768 3213 34836
rect 3137 34712 3147 34768
rect 3203 34712 3213 34768
rect 3137 34644 3213 34712
rect 3137 34588 3147 34644
rect 3203 34588 3213 34644
rect 3137 34520 3213 34588
rect 3137 34464 3147 34520
rect 3203 34464 3213 34520
rect 3137 34396 3213 34464
rect 3137 34340 3147 34396
rect 3203 34340 3213 34396
rect 3137 34272 3213 34340
rect 3137 34216 3147 34272
rect 3203 34216 3213 34272
rect 3137 34148 3213 34216
rect 3137 34092 3147 34148
rect 3203 34092 3213 34148
rect 3137 34024 3213 34092
rect 3137 33968 3147 34024
rect 3203 33968 3213 34024
rect 3137 33900 3213 33968
rect 3137 33844 3147 33900
rect 3203 33844 3213 33900
rect 3137 33776 3213 33844
rect 3137 33720 3147 33776
rect 3203 33720 3213 33776
rect 3137 33652 3213 33720
rect 3137 33596 3147 33652
rect 3203 33596 3213 33652
rect 3137 33528 3213 33596
rect 3137 33472 3147 33528
rect 3203 33472 3213 33528
rect 3137 33404 3213 33472
rect 3137 33348 3147 33404
rect 3203 33348 3213 33404
rect 3137 33280 3213 33348
rect 3137 33224 3147 33280
rect 3203 33224 3213 33280
rect 3137 33156 3213 33224
rect 3137 33100 3147 33156
rect 3203 33100 3213 33156
rect 3137 33032 3213 33100
rect 3137 32976 3147 33032
rect 3203 32976 3213 33032
rect 3137 32908 3213 32976
rect 3137 32852 3147 32908
rect 3203 32852 3213 32908
rect 3137 32784 3213 32852
rect 3137 32728 3147 32784
rect 3203 32728 3213 32784
rect 3137 32660 3213 32728
rect 3137 32604 3147 32660
rect 3203 32604 3213 32660
rect 3137 32536 3213 32604
rect 3137 32480 3147 32536
rect 3203 32480 3213 32536
rect 2013 32402 2089 32470
rect 2013 32346 2023 32402
rect 2079 32346 2089 32402
rect 3137 32412 3213 32480
rect 3137 32356 3147 32412
rect 3203 32356 3213 32412
rect 3137 32346 3213 32356
rect 3261 36256 3337 36266
rect 3261 36200 3271 36256
rect 3327 36200 3337 36256
rect 3261 36132 3337 36200
rect 3261 36076 3271 36132
rect 3327 36076 3337 36132
rect 3261 36008 3337 36076
rect 3261 35952 3271 36008
rect 3327 35952 3337 36008
rect 3261 35884 3337 35952
rect 3261 35828 3271 35884
rect 3327 35828 3337 35884
rect 3261 35760 3337 35828
rect 3261 35704 3271 35760
rect 3327 35704 3337 35760
rect 3261 35636 3337 35704
rect 3261 35580 3271 35636
rect 3327 35580 3337 35636
rect 3261 35512 3337 35580
rect 3261 35456 3271 35512
rect 3327 35456 3337 35512
rect 3261 35388 3337 35456
rect 3261 35332 3271 35388
rect 3327 35332 3337 35388
rect 3261 35264 3337 35332
rect 3261 35208 3271 35264
rect 3327 35208 3337 35264
rect 3261 35140 3337 35208
rect 3261 35084 3271 35140
rect 3327 35084 3337 35140
rect 3261 35016 3337 35084
rect 3261 34960 3271 35016
rect 3327 34960 3337 35016
rect 3261 34892 3337 34960
rect 3261 34836 3271 34892
rect 3327 34836 3337 34892
rect 3261 34768 3337 34836
rect 3261 34712 3271 34768
rect 3327 34712 3337 34768
rect 3261 34644 3337 34712
rect 3261 34588 3271 34644
rect 3327 34588 3337 34644
rect 3261 34520 3337 34588
rect 3261 34464 3271 34520
rect 3327 34464 3337 34520
rect 3261 34396 3337 34464
rect 3261 34340 3271 34396
rect 3327 34340 3337 34396
rect 3261 34272 3337 34340
rect 3261 34216 3271 34272
rect 3327 34216 3337 34272
rect 3261 34148 3337 34216
rect 3261 34092 3271 34148
rect 3327 34092 3337 34148
rect 3261 34024 3337 34092
rect 3261 33968 3271 34024
rect 3327 33968 3337 34024
rect 3261 33900 3337 33968
rect 3261 33844 3271 33900
rect 3327 33844 3337 33900
rect 3261 33776 3337 33844
rect 3261 33720 3271 33776
rect 3327 33720 3337 33776
rect 3261 33652 3337 33720
rect 3261 33596 3271 33652
rect 3327 33596 3337 33652
rect 3261 33528 3337 33596
rect 3261 33472 3271 33528
rect 3327 33472 3337 33528
rect 3261 33404 3337 33472
rect 3261 33348 3271 33404
rect 3327 33348 3337 33404
rect 3261 33280 3337 33348
rect 3261 33224 3271 33280
rect 3327 33224 3337 33280
rect 3261 33156 3337 33224
rect 3261 33100 3271 33156
rect 3327 33100 3337 33156
rect 3261 33032 3337 33100
rect 3261 32976 3271 33032
rect 3327 32976 3337 33032
rect 3261 32908 3337 32976
rect 3261 32852 3271 32908
rect 3327 32852 3337 32908
rect 3261 32784 3337 32852
rect 3261 32728 3271 32784
rect 3327 32728 3337 32784
rect 3261 32660 3337 32728
rect 3261 32604 3271 32660
rect 3327 32604 3337 32660
rect 3261 32536 3337 32604
rect 3261 32480 3271 32536
rect 3327 32480 3337 32536
rect 3261 32412 3337 32480
rect 3261 32356 3271 32412
rect 3327 32356 3337 32412
rect 2013 32278 2089 32346
rect 2013 32222 2023 32278
rect 2079 32222 2089 32278
rect 3261 32288 3337 32356
rect 3261 32232 3271 32288
rect 3327 32232 3337 32288
rect 3261 32222 3337 32232
rect 3385 36132 3461 36142
rect 3385 36076 3395 36132
rect 3451 36076 3461 36132
rect 3385 36008 3461 36076
rect 3385 35952 3395 36008
rect 3451 35952 3461 36008
rect 3385 35884 3461 35952
rect 3385 35828 3395 35884
rect 3451 35828 3461 35884
rect 3385 35760 3461 35828
rect 3385 35704 3395 35760
rect 3451 35704 3461 35760
rect 3385 35636 3461 35704
rect 3385 35580 3395 35636
rect 3451 35580 3461 35636
rect 3385 35512 3461 35580
rect 3385 35456 3395 35512
rect 3451 35456 3461 35512
rect 3385 35388 3461 35456
rect 3385 35332 3395 35388
rect 3451 35332 3461 35388
rect 3385 35264 3461 35332
rect 3385 35208 3395 35264
rect 3451 35208 3461 35264
rect 3385 35140 3461 35208
rect 3385 35084 3395 35140
rect 3451 35084 3461 35140
rect 3385 35016 3461 35084
rect 3385 34960 3395 35016
rect 3451 34960 3461 35016
rect 3385 34892 3461 34960
rect 3385 34836 3395 34892
rect 3451 34836 3461 34892
rect 3385 34768 3461 34836
rect 3385 34712 3395 34768
rect 3451 34712 3461 34768
rect 3385 34644 3461 34712
rect 3385 34588 3395 34644
rect 3451 34588 3461 34644
rect 3385 34520 3461 34588
rect 3385 34464 3395 34520
rect 3451 34464 3461 34520
rect 3385 34396 3461 34464
rect 3385 34340 3395 34396
rect 3451 34340 3461 34396
rect 3385 34272 3461 34340
rect 3385 34216 3395 34272
rect 3451 34216 3461 34272
rect 3385 34148 3461 34216
rect 3385 34092 3395 34148
rect 3451 34092 3461 34148
rect 3385 34024 3461 34092
rect 3385 33968 3395 34024
rect 3451 33968 3461 34024
rect 3385 33900 3461 33968
rect 3385 33844 3395 33900
rect 3451 33844 3461 33900
rect 3385 33776 3461 33844
rect 3385 33720 3395 33776
rect 3451 33720 3461 33776
rect 3385 33652 3461 33720
rect 3385 33596 3395 33652
rect 3451 33596 3461 33652
rect 3385 33528 3461 33596
rect 3385 33472 3395 33528
rect 3451 33472 3461 33528
rect 3385 33404 3461 33472
rect 3385 33348 3395 33404
rect 3451 33348 3461 33404
rect 3385 33280 3461 33348
rect 3385 33224 3395 33280
rect 3451 33224 3461 33280
rect 3385 33156 3461 33224
rect 3385 33100 3395 33156
rect 3451 33100 3461 33156
rect 3385 33032 3461 33100
rect 3385 32976 3395 33032
rect 3451 32976 3461 33032
rect 3385 32908 3461 32976
rect 3385 32852 3395 32908
rect 3451 32852 3461 32908
rect 3385 32784 3461 32852
rect 3385 32728 3395 32784
rect 3451 32728 3461 32784
rect 3385 32660 3461 32728
rect 3385 32604 3395 32660
rect 3451 32604 3461 32660
rect 3385 32536 3461 32604
rect 3385 32480 3395 32536
rect 3451 32480 3461 32536
rect 3385 32412 3461 32480
rect 3385 32356 3395 32412
rect 3451 32356 3461 32412
rect 3385 32288 3461 32356
rect 3385 32232 3395 32288
rect 3451 32232 3461 32288
rect 2013 32154 2089 32222
rect 2013 32098 2023 32154
rect 2079 32098 2089 32154
rect 3385 32164 3461 32232
rect 3385 32108 3395 32164
rect 3451 32108 3461 32164
rect 3385 32098 3461 32108
rect 3509 35946 3585 35956
rect 3509 35890 3519 35946
rect 3575 35890 3585 35946
rect 3509 35822 3585 35890
rect 3509 35766 3519 35822
rect 3575 35766 3585 35822
rect 3509 35698 3585 35766
rect 3509 35642 3519 35698
rect 3575 35642 3585 35698
rect 3509 35574 3585 35642
rect 3509 35518 3519 35574
rect 3575 35518 3585 35574
rect 3509 35450 3585 35518
rect 3509 35394 3519 35450
rect 3575 35394 3585 35450
rect 3509 35326 3585 35394
rect 3509 35270 3519 35326
rect 3575 35270 3585 35326
rect 3509 35202 3585 35270
rect 3509 35146 3519 35202
rect 3575 35146 3585 35202
rect 3509 35078 3585 35146
rect 3509 35022 3519 35078
rect 3575 35022 3585 35078
rect 3509 34954 3585 35022
rect 3509 34898 3519 34954
rect 3575 34898 3585 34954
rect 3509 34830 3585 34898
rect 3509 34774 3519 34830
rect 3575 34774 3585 34830
rect 3509 34706 3585 34774
rect 3509 34650 3519 34706
rect 3575 34650 3585 34706
rect 3509 34582 3585 34650
rect 3509 34526 3519 34582
rect 3575 34526 3585 34582
rect 3509 34458 3585 34526
rect 3509 34402 3519 34458
rect 3575 34402 3585 34458
rect 3509 34334 3585 34402
rect 3509 34278 3519 34334
rect 3575 34278 3585 34334
rect 3509 34210 3585 34278
rect 3509 34154 3519 34210
rect 3575 34154 3585 34210
rect 3509 34086 3585 34154
rect 3509 34030 3519 34086
rect 3575 34030 3585 34086
rect 3509 33962 3585 34030
rect 3509 33906 3519 33962
rect 3575 33906 3585 33962
rect 3509 33838 3585 33906
rect 3509 33782 3519 33838
rect 3575 33782 3585 33838
rect 3509 33714 3585 33782
rect 3509 33658 3519 33714
rect 3575 33658 3585 33714
rect 3509 33590 3585 33658
rect 3509 33534 3519 33590
rect 3575 33534 3585 33590
rect 3509 33466 3585 33534
rect 3509 33410 3519 33466
rect 3575 33410 3585 33466
rect 3509 33342 3585 33410
rect 3509 33286 3519 33342
rect 3575 33286 3585 33342
rect 3509 33218 3585 33286
rect 3509 33162 3519 33218
rect 3575 33162 3585 33218
rect 3509 33094 3585 33162
rect 3509 33038 3519 33094
rect 3575 33038 3585 33094
rect 3509 32970 3585 33038
rect 3509 32914 3519 32970
rect 3575 32914 3585 32970
rect 3509 32846 3585 32914
rect 3509 32790 3519 32846
rect 3575 32790 3585 32846
rect 3509 32722 3585 32790
rect 3509 32666 3519 32722
rect 3575 32666 3585 32722
rect 3509 32598 3585 32666
rect 3509 32542 3519 32598
rect 3575 32542 3585 32598
rect 3509 32474 3585 32542
rect 3509 32418 3519 32474
rect 3575 32418 3585 32474
rect 3509 32350 3585 32418
rect 3509 32294 3519 32350
rect 3575 32294 3585 32350
rect 3509 32226 3585 32294
rect 3509 32170 3519 32226
rect 3575 32170 3585 32226
rect 3509 32102 3585 32170
rect 2013 32030 2089 32098
rect 3509 32046 3519 32102
rect 3575 32046 3585 32102
rect 3509 32036 3585 32046
rect 3633 35813 3709 35823
rect 3633 35757 3643 35813
rect 3699 35757 3709 35813
rect 3633 35689 3709 35757
rect 3633 35633 3643 35689
rect 3699 35633 3709 35689
rect 3633 35565 3709 35633
rect 3633 35509 3643 35565
rect 3699 35509 3709 35565
rect 3633 35441 3709 35509
rect 3633 35385 3643 35441
rect 3699 35385 3709 35441
rect 3633 35317 3709 35385
rect 3633 35261 3643 35317
rect 3699 35261 3709 35317
rect 3633 35193 3709 35261
rect 3633 35137 3643 35193
rect 3699 35137 3709 35193
rect 3633 35069 3709 35137
rect 3633 35013 3643 35069
rect 3699 35013 3709 35069
rect 3633 34945 3709 35013
rect 3633 34889 3643 34945
rect 3699 34889 3709 34945
rect 3633 34821 3709 34889
rect 3633 34765 3643 34821
rect 3699 34765 3709 34821
rect 3633 34697 3709 34765
rect 3633 34641 3643 34697
rect 3699 34641 3709 34697
rect 3633 34573 3709 34641
rect 3633 34517 3643 34573
rect 3699 34517 3709 34573
rect 3633 34449 3709 34517
rect 3633 34393 3643 34449
rect 3699 34393 3709 34449
rect 3633 34325 3709 34393
rect 3633 34269 3643 34325
rect 3699 34269 3709 34325
rect 3633 34201 3709 34269
rect 3633 34145 3643 34201
rect 3699 34145 3709 34201
rect 3633 34077 3709 34145
rect 3633 34021 3643 34077
rect 3699 34021 3709 34077
rect 3633 33953 3709 34021
rect 3633 33897 3643 33953
rect 3699 33897 3709 33953
rect 3633 33829 3709 33897
rect 3633 33773 3643 33829
rect 3699 33773 3709 33829
rect 3633 33705 3709 33773
rect 3633 33649 3643 33705
rect 3699 33649 3709 33705
rect 3633 33581 3709 33649
rect 3633 33525 3643 33581
rect 3699 33525 3709 33581
rect 3633 33457 3709 33525
rect 3633 33401 3643 33457
rect 3699 33401 3709 33457
rect 3633 33333 3709 33401
rect 3633 33277 3643 33333
rect 3699 33277 3709 33333
rect 3633 33209 3709 33277
rect 3633 33153 3643 33209
rect 3699 33153 3709 33209
rect 3633 33085 3709 33153
rect 3633 33029 3643 33085
rect 3699 33029 3709 33085
rect 3633 32961 3709 33029
rect 3633 32905 3643 32961
rect 3699 32905 3709 32961
rect 3633 32837 3709 32905
rect 3633 32781 3643 32837
rect 3699 32781 3709 32837
rect 3633 32713 3709 32781
rect 3633 32657 3643 32713
rect 3699 32657 3709 32713
rect 3633 32589 3709 32657
rect 3633 32533 3643 32589
rect 3699 32533 3709 32589
rect 3633 32465 3709 32533
rect 3633 32409 3643 32465
rect 3699 32409 3709 32465
rect 3633 32341 3709 32409
rect 3633 32285 3643 32341
rect 3699 32285 3709 32341
rect 3633 32217 3709 32285
rect 3633 32161 3643 32217
rect 3699 32161 3709 32217
rect 3633 32093 3709 32161
rect 3633 32037 3643 32093
rect 3699 32037 3709 32093
rect 3757 35710 3833 35720
rect 3757 35654 3767 35710
rect 3823 35654 3833 35710
rect 3757 35586 3833 35654
rect 3757 35530 3767 35586
rect 3823 35530 3833 35586
rect 3757 35462 3833 35530
rect 3757 35406 3767 35462
rect 3823 35406 3833 35462
rect 3757 35338 3833 35406
rect 3757 35282 3767 35338
rect 3823 35282 3833 35338
rect 3757 35214 3833 35282
rect 3757 35158 3767 35214
rect 3823 35158 3833 35214
rect 3757 35090 3833 35158
rect 3757 35034 3767 35090
rect 3823 35034 3833 35090
rect 3757 34966 3833 35034
rect 3757 34910 3767 34966
rect 3823 34910 3833 34966
rect 3757 34842 3833 34910
rect 3757 34786 3767 34842
rect 3823 34786 3833 34842
rect 3757 34718 3833 34786
rect 3757 34662 3767 34718
rect 3823 34662 3833 34718
rect 3757 34594 3833 34662
rect 3757 34538 3767 34594
rect 3823 34538 3833 34594
rect 3757 34470 3833 34538
rect 3757 34414 3767 34470
rect 3823 34414 3833 34470
rect 3757 34346 3833 34414
rect 3757 34290 3767 34346
rect 3823 34290 3833 34346
rect 3757 34222 3833 34290
rect 3757 34166 3767 34222
rect 3823 34166 3833 34222
rect 3757 34098 3833 34166
rect 3757 34042 3767 34098
rect 3823 34042 3833 34098
rect 3757 33974 3833 34042
rect 3757 33918 3767 33974
rect 3823 33918 3833 33974
rect 3757 33850 3833 33918
rect 3757 33794 3767 33850
rect 3823 33794 3833 33850
rect 3757 33726 3833 33794
rect 3757 33670 3767 33726
rect 3823 33670 3833 33726
rect 3757 33602 3833 33670
rect 3757 33546 3767 33602
rect 3823 33546 3833 33602
rect 3757 33478 3833 33546
rect 3757 33422 3767 33478
rect 3823 33422 3833 33478
rect 3757 33354 3833 33422
rect 3757 33298 3767 33354
rect 3823 33298 3833 33354
rect 3757 33230 3833 33298
rect 3757 33174 3767 33230
rect 3823 33174 3833 33230
rect 3757 33106 3833 33174
rect 3757 33050 3767 33106
rect 3823 33050 3833 33106
rect 3757 32982 3833 33050
rect 3757 32926 3767 32982
rect 3823 32926 3833 32982
rect 3757 32858 3833 32926
rect 3757 32802 3767 32858
rect 3823 32802 3833 32858
rect 3757 32734 3833 32802
rect 3757 32678 3767 32734
rect 3823 32678 3833 32734
rect 3757 32610 3833 32678
rect 3757 32554 3767 32610
rect 3823 32554 3833 32610
rect 3757 32486 3833 32554
rect 3757 32430 3767 32486
rect 3823 32430 3833 32486
rect 3757 32362 3833 32430
rect 3757 32306 3767 32362
rect 3823 32306 3833 32362
rect 3757 32238 3833 32306
rect 3757 32182 3767 32238
rect 3823 32182 3833 32238
rect 3757 32114 3833 32182
rect 3757 32058 3767 32114
rect 3823 32058 3833 32114
rect 3881 35606 3957 35616
rect 3881 35550 3891 35606
rect 3947 35550 3957 35606
rect 3881 35482 3957 35550
rect 3881 35426 3891 35482
rect 3947 35426 3957 35482
rect 3881 35358 3957 35426
rect 3881 35302 3891 35358
rect 3947 35302 3957 35358
rect 3881 35234 3957 35302
rect 3881 35178 3891 35234
rect 3947 35178 3957 35234
rect 3881 35110 3957 35178
rect 3881 35054 3891 35110
rect 3947 35054 3957 35110
rect 3881 34986 3957 35054
rect 3881 34930 3891 34986
rect 3947 34930 3957 34986
rect 3881 34862 3957 34930
rect 3881 34806 3891 34862
rect 3947 34806 3957 34862
rect 3881 34738 3957 34806
rect 3881 34682 3891 34738
rect 3947 34682 3957 34738
rect 3881 34614 3957 34682
rect 3881 34558 3891 34614
rect 3947 34558 3957 34614
rect 3881 34490 3957 34558
rect 3881 34434 3891 34490
rect 3947 34434 3957 34490
rect 3881 34366 3957 34434
rect 3881 34310 3891 34366
rect 3947 34310 3957 34366
rect 3881 34242 3957 34310
rect 3881 34186 3891 34242
rect 3947 34186 3957 34242
rect 3881 34118 3957 34186
rect 3881 34062 3891 34118
rect 3947 34062 3957 34118
rect 3881 33994 3957 34062
rect 3881 33938 3891 33994
rect 3947 33938 3957 33994
rect 3881 33870 3957 33938
rect 3881 33814 3891 33870
rect 3947 33814 3957 33870
rect 3881 33746 3957 33814
rect 3881 33690 3891 33746
rect 3947 33690 3957 33746
rect 3881 33622 3957 33690
rect 3881 33566 3891 33622
rect 3947 33566 3957 33622
rect 3881 33498 3957 33566
rect 3881 33442 3891 33498
rect 3947 33442 3957 33498
rect 3881 33374 3957 33442
rect 3881 33318 3891 33374
rect 3947 33318 3957 33374
rect 3881 33250 3957 33318
rect 3881 33194 3891 33250
rect 3947 33194 3957 33250
rect 3881 33126 3957 33194
rect 3881 33070 3891 33126
rect 3947 33070 3957 33126
rect 3881 33002 3957 33070
rect 3881 32946 3891 33002
rect 3947 32946 3957 33002
rect 3881 32878 3957 32946
rect 3881 32822 3891 32878
rect 3947 32822 3957 32878
rect 3881 32754 3957 32822
rect 3881 32698 3891 32754
rect 3947 32698 3957 32754
rect 3881 32630 3957 32698
rect 3881 32574 3891 32630
rect 3947 32574 3957 32630
rect 3881 32506 3957 32574
rect 3881 32450 3891 32506
rect 3947 32450 3957 32506
rect 3881 32382 3957 32450
rect 3881 32326 3891 32382
rect 3947 32326 3957 32382
rect 3881 32258 3957 32326
rect 3881 32202 3891 32258
rect 3947 32202 3957 32258
rect 3881 32134 3957 32202
rect 3881 32078 3891 32134
rect 3947 32078 3957 32134
rect 3881 32068 3957 32078
rect 4005 35535 4081 35545
rect 4005 35479 4015 35535
rect 4071 35479 4081 35535
rect 4005 35411 4081 35479
rect 4005 35355 4015 35411
rect 4071 35355 4081 35411
rect 4005 35287 4081 35355
rect 4005 35231 4015 35287
rect 4071 35231 4081 35287
rect 4005 35163 4081 35231
rect 4005 35107 4015 35163
rect 4071 35107 4081 35163
rect 4005 35039 4081 35107
rect 4005 34983 4015 35039
rect 4071 34983 4081 35039
rect 4005 34915 4081 34983
rect 4005 34859 4015 34915
rect 4071 34859 4081 34915
rect 4005 34791 4081 34859
rect 4005 34735 4015 34791
rect 4071 34735 4081 34791
rect 4005 34667 4081 34735
rect 4005 34611 4015 34667
rect 4071 34611 4081 34667
rect 4005 34543 4081 34611
rect 4005 34487 4015 34543
rect 4071 34487 4081 34543
rect 4005 34419 4081 34487
rect 4005 34363 4015 34419
rect 4071 34363 4081 34419
rect 4005 34295 4081 34363
rect 4005 34239 4015 34295
rect 4071 34239 4081 34295
rect 4005 34171 4081 34239
rect 4005 34115 4015 34171
rect 4071 34115 4081 34171
rect 4005 34047 4081 34115
rect 4005 33991 4015 34047
rect 4071 33991 4081 34047
rect 4005 33923 4081 33991
rect 4005 33867 4015 33923
rect 4071 33867 4081 33923
rect 4005 33799 4081 33867
rect 4005 33743 4015 33799
rect 4071 33743 4081 33799
rect 4005 33675 4081 33743
rect 4005 33619 4015 33675
rect 4071 33619 4081 33675
rect 4005 33551 4081 33619
rect 4005 33495 4015 33551
rect 4071 33495 4081 33551
rect 4005 33427 4081 33495
rect 4005 33371 4015 33427
rect 4071 33371 4081 33427
rect 4005 33303 4081 33371
rect 4005 33247 4015 33303
rect 4071 33247 4081 33303
rect 4005 33179 4081 33247
rect 4005 33123 4015 33179
rect 4071 33123 4081 33179
rect 4005 33055 4081 33123
rect 4005 32999 4015 33055
rect 4071 32999 4081 33055
rect 4005 32931 4081 32999
rect 4005 32875 4015 32931
rect 4071 32875 4081 32931
rect 4005 32807 4081 32875
rect 4005 32751 4015 32807
rect 4071 32751 4081 32807
rect 4005 32683 4081 32751
rect 4005 32627 4015 32683
rect 4071 32627 4081 32683
rect 4005 32559 4081 32627
rect 4005 32503 4015 32559
rect 4071 32503 4081 32559
rect 4005 32435 4081 32503
rect 4005 32379 4015 32435
rect 4071 32379 4081 32435
rect 4005 32311 4081 32379
rect 4005 32255 4015 32311
rect 4071 32255 4081 32311
rect 4005 32187 4081 32255
rect 4005 32131 4015 32187
rect 4071 32131 4081 32187
rect 3757 32048 3833 32058
rect 4005 32063 4081 32131
rect 2013 31974 2023 32030
rect 2079 31974 2089 32030
rect 3633 32027 3709 32037
rect 4005 32007 4015 32063
rect 4071 32007 4081 32063
rect 4005 31997 4081 32007
rect 4129 35417 4205 35427
rect 4129 35361 4139 35417
rect 4195 35361 4205 35417
rect 4129 35293 4205 35361
rect 4129 35237 4139 35293
rect 4195 35237 4205 35293
rect 4129 35169 4205 35237
rect 14757 35220 14767 36572
rect 14823 35220 14833 36572
rect 14757 35210 14833 35220
rect 4129 35113 4139 35169
rect 4195 35113 4205 35169
rect 4129 35045 4205 35113
rect 4129 34989 4139 35045
rect 4195 34989 4205 35045
rect 4129 34921 4205 34989
rect 4129 34865 4139 34921
rect 4195 34865 4205 34921
rect 4129 34797 4205 34865
rect 4129 34741 4139 34797
rect 4195 34741 4205 34797
rect 4129 34673 4205 34741
rect 4129 34617 4139 34673
rect 4195 34617 4205 34673
rect 4129 34549 4205 34617
rect 4129 34493 4139 34549
rect 4195 34493 4205 34549
rect 4129 34425 4205 34493
rect 4129 34369 4139 34425
rect 4195 34369 4205 34425
rect 4129 34301 4205 34369
rect 4129 34245 4139 34301
rect 4195 34245 4205 34301
rect 4129 34177 4205 34245
rect 4129 34121 4139 34177
rect 4195 34121 4205 34177
rect 4129 34053 4205 34121
rect 4129 33997 4139 34053
rect 4195 33997 4205 34053
rect 4129 33929 4205 33997
rect 4129 33873 4139 33929
rect 4195 33873 4205 33929
rect 4129 33805 4205 33873
rect 4129 33749 4139 33805
rect 4195 33749 4205 33805
rect 4129 33681 4205 33749
rect 4129 33625 4139 33681
rect 4195 33625 4205 33681
rect 4129 33557 4205 33625
rect 4129 33501 4139 33557
rect 4195 33501 4205 33557
rect 4129 33433 4205 33501
rect 4129 33377 4139 33433
rect 4195 33377 4205 33433
rect 4129 33309 4205 33377
rect 4129 33253 4139 33309
rect 4195 33253 4205 33309
rect 4129 33185 4205 33253
rect 4129 33129 4139 33185
rect 4195 33129 4205 33185
rect 4129 33061 4205 33129
rect 4129 33005 4139 33061
rect 4195 33005 4205 33061
rect 4129 32937 4205 33005
rect 4129 32881 4139 32937
rect 4195 32881 4205 32937
rect 4129 32813 4205 32881
rect 4129 32757 4139 32813
rect 4195 32757 4205 32813
rect 4129 32689 4205 32757
rect 4129 32633 4139 32689
rect 4195 32633 4205 32689
rect 4129 32565 4205 32633
rect 4129 32509 4139 32565
rect 4195 32509 4205 32565
rect 4129 32441 4205 32509
rect 4129 32385 4139 32441
rect 4195 32385 4205 32441
rect 4129 32317 4205 32385
rect 4129 32261 4139 32317
rect 4195 32261 4205 32317
rect 4129 32193 4205 32261
rect 4129 32137 4139 32193
rect 4195 32137 4205 32193
rect 4129 32069 4205 32137
rect 4129 32013 4139 32069
rect 4195 32013 4205 32069
rect 6358 34950 7426 34960
rect 6358 34894 6368 34950
rect 6424 34894 6492 34950
rect 6548 34894 6616 34950
rect 6672 34894 6740 34950
rect 6796 34894 6864 34950
rect 6920 34894 6988 34950
rect 7044 34894 7112 34950
rect 7168 34894 7236 34950
rect 7292 34894 7360 34950
rect 7416 34894 7426 34950
rect 6358 34826 7426 34894
rect 6358 34770 6368 34826
rect 6424 34770 6492 34826
rect 6548 34770 6616 34826
rect 6672 34770 6740 34826
rect 6796 34770 6864 34826
rect 6920 34770 6988 34826
rect 7044 34770 7112 34826
rect 7168 34770 7236 34826
rect 7292 34770 7360 34826
rect 7416 34770 7426 34826
rect 6358 34702 7426 34770
rect 6358 34646 6368 34702
rect 6424 34646 6492 34702
rect 6548 34646 6616 34702
rect 6672 34646 6740 34702
rect 6796 34646 6864 34702
rect 6920 34646 6988 34702
rect 7044 34646 7112 34702
rect 7168 34646 7236 34702
rect 7292 34646 7360 34702
rect 7416 34646 7426 34702
rect 6358 34578 7426 34646
rect 6358 34522 6368 34578
rect 6424 34522 6492 34578
rect 6548 34522 6616 34578
rect 6672 34522 6740 34578
rect 6796 34522 6864 34578
rect 6920 34522 6988 34578
rect 7044 34522 7112 34578
rect 7168 34522 7236 34578
rect 7292 34522 7360 34578
rect 7416 34522 7426 34578
rect 6358 34454 7426 34522
rect 6358 34398 6368 34454
rect 6424 34398 6492 34454
rect 6548 34398 6616 34454
rect 6672 34398 6740 34454
rect 6796 34398 6864 34454
rect 6920 34398 6988 34454
rect 7044 34398 7112 34454
rect 7168 34398 7236 34454
rect 7292 34398 7360 34454
rect 7416 34398 7426 34454
rect 6358 34330 7426 34398
rect 6358 34274 6368 34330
rect 6424 34274 6492 34330
rect 6548 34274 6616 34330
rect 6672 34274 6740 34330
rect 6796 34274 6864 34330
rect 6920 34274 6988 34330
rect 7044 34274 7112 34330
rect 7168 34274 7236 34330
rect 7292 34274 7360 34330
rect 7416 34274 7426 34330
rect 6358 34206 7426 34274
rect 6358 34150 6368 34206
rect 6424 34150 6492 34206
rect 6548 34150 6616 34206
rect 6672 34150 6740 34206
rect 6796 34150 6864 34206
rect 6920 34150 6988 34206
rect 7044 34150 7112 34206
rect 7168 34150 7236 34206
rect 7292 34150 7360 34206
rect 7416 34150 7426 34206
rect 6358 34082 7426 34150
rect 6358 34026 6368 34082
rect 6424 34026 6492 34082
rect 6548 34026 6616 34082
rect 6672 34026 6740 34082
rect 6796 34026 6864 34082
rect 6920 34026 6988 34082
rect 7044 34026 7112 34082
rect 7168 34026 7236 34082
rect 7292 34026 7360 34082
rect 7416 34026 7426 34082
rect 6358 33958 7426 34026
rect 6358 33902 6368 33958
rect 6424 33902 6492 33958
rect 6548 33902 6616 33958
rect 6672 33902 6740 33958
rect 6796 33902 6864 33958
rect 6920 33902 6988 33958
rect 7044 33902 7112 33958
rect 7168 33902 7236 33958
rect 7292 33902 7360 33958
rect 7416 33902 7426 33958
rect 6358 33834 7426 33902
rect 6358 33778 6368 33834
rect 6424 33778 6492 33834
rect 6548 33778 6616 33834
rect 6672 33778 6740 33834
rect 6796 33778 6864 33834
rect 6920 33778 6988 33834
rect 7044 33778 7112 33834
rect 7168 33778 7236 33834
rect 7292 33778 7360 33834
rect 7416 33778 7426 33834
rect 6358 33710 7426 33778
rect 6358 33654 6368 33710
rect 6424 33654 6492 33710
rect 6548 33654 6616 33710
rect 6672 33654 6740 33710
rect 6796 33654 6864 33710
rect 6920 33654 6988 33710
rect 7044 33654 7112 33710
rect 7168 33654 7236 33710
rect 7292 33654 7360 33710
rect 7416 33654 7426 33710
rect 6358 33586 7426 33654
rect 6358 33530 6368 33586
rect 6424 33530 6492 33586
rect 6548 33530 6616 33586
rect 6672 33530 6740 33586
rect 6796 33530 6864 33586
rect 6920 33530 6988 33586
rect 7044 33530 7112 33586
rect 7168 33530 7236 33586
rect 7292 33530 7360 33586
rect 7416 33530 7426 33586
rect 6358 33462 7426 33530
rect 6358 33406 6368 33462
rect 6424 33406 6492 33462
rect 6548 33406 6616 33462
rect 6672 33406 6740 33462
rect 6796 33406 6864 33462
rect 6920 33406 6988 33462
rect 7044 33406 7112 33462
rect 7168 33406 7236 33462
rect 7292 33406 7360 33462
rect 7416 33406 7426 33462
rect 6358 33338 7426 33406
rect 6358 33282 6368 33338
rect 6424 33282 6492 33338
rect 6548 33282 6616 33338
rect 6672 33282 6740 33338
rect 6796 33282 6864 33338
rect 6920 33282 6988 33338
rect 7044 33282 7112 33338
rect 7168 33282 7236 33338
rect 7292 33282 7360 33338
rect 7416 33282 7426 33338
rect 6358 33214 7426 33282
rect 6358 33158 6368 33214
rect 6424 33158 6492 33214
rect 6548 33158 6616 33214
rect 6672 33158 6740 33214
rect 6796 33158 6864 33214
rect 6920 33158 6988 33214
rect 7044 33158 7112 33214
rect 7168 33158 7236 33214
rect 7292 33158 7360 33214
rect 7416 33158 7426 33214
rect 6358 33090 7426 33158
rect 6358 33034 6368 33090
rect 6424 33034 6492 33090
rect 6548 33034 6616 33090
rect 6672 33034 6740 33090
rect 6796 33034 6864 33090
rect 6920 33034 6988 33090
rect 7044 33034 7112 33090
rect 7168 33034 7236 33090
rect 7292 33034 7360 33090
rect 7416 33034 7426 33090
rect 6358 32966 7426 33034
rect 6358 32910 6368 32966
rect 6424 32910 6492 32966
rect 6548 32910 6616 32966
rect 6672 32910 6740 32966
rect 6796 32910 6864 32966
rect 6920 32910 6988 32966
rect 7044 32910 7112 32966
rect 7168 32910 7236 32966
rect 7292 32910 7360 32966
rect 7416 32910 7426 32966
rect 6358 32842 7426 32910
rect 6358 32786 6368 32842
rect 6424 32786 6492 32842
rect 6548 32786 6616 32842
rect 6672 32786 6740 32842
rect 6796 32786 6864 32842
rect 6920 32786 6988 32842
rect 7044 32786 7112 32842
rect 7168 32786 7236 32842
rect 7292 32786 7360 32842
rect 7416 32786 7426 32842
rect 6358 32718 7426 32786
rect 6358 32662 6368 32718
rect 6424 32662 6492 32718
rect 6548 32662 6616 32718
rect 6672 32662 6740 32718
rect 6796 32662 6864 32718
rect 6920 32662 6988 32718
rect 7044 32662 7112 32718
rect 7168 32662 7236 32718
rect 7292 32662 7360 32718
rect 7416 32662 7426 32718
rect 6358 32594 7426 32662
rect 6358 32538 6368 32594
rect 6424 32538 6492 32594
rect 6548 32538 6616 32594
rect 6672 32538 6740 32594
rect 6796 32538 6864 32594
rect 6920 32538 6988 32594
rect 7044 32538 7112 32594
rect 7168 32538 7236 32594
rect 7292 32538 7360 32594
rect 7416 32538 7426 32594
rect 6358 32470 7426 32538
rect 6358 32414 6368 32470
rect 6424 32414 6492 32470
rect 6548 32414 6616 32470
rect 6672 32414 6740 32470
rect 6796 32414 6864 32470
rect 6920 32414 6988 32470
rect 7044 32414 7112 32470
rect 7168 32414 7236 32470
rect 7292 32414 7360 32470
rect 7416 32414 7426 32470
rect 6358 32346 7426 32414
rect 6358 32290 6368 32346
rect 6424 32290 6492 32346
rect 6548 32290 6616 32346
rect 6672 32290 6740 32346
rect 6796 32290 6864 32346
rect 6920 32290 6988 32346
rect 7044 32290 7112 32346
rect 7168 32290 7236 32346
rect 7292 32290 7360 32346
rect 7416 32290 7426 32346
rect 6358 32222 7426 32290
rect 6358 32166 6368 32222
rect 6424 32166 6492 32222
rect 6548 32166 6616 32222
rect 6672 32166 6740 32222
rect 6796 32166 6864 32222
rect 6920 32166 6988 32222
rect 7044 32166 7112 32222
rect 7168 32166 7236 32222
rect 7292 32166 7360 32222
rect 7416 32166 7426 32222
rect 6358 32098 7426 32166
rect 6358 32042 6368 32098
rect 6424 32042 6492 32098
rect 6548 32042 6616 32098
rect 6672 32042 6740 32098
rect 6796 32042 6864 32098
rect 6920 32042 6988 32098
rect 7044 32042 7112 32098
rect 7168 32042 7236 32098
rect 7292 32042 7360 32098
rect 7416 32042 7426 32098
rect 6358 32032 7426 32042
rect 8741 34950 10553 34960
rect 8741 34894 8751 34950
rect 8807 34894 8875 34950
rect 8931 34894 8999 34950
rect 9055 34894 9123 34950
rect 9179 34894 9247 34950
rect 9303 34894 9371 34950
rect 9427 34894 9495 34950
rect 9551 34894 9619 34950
rect 9675 34894 9743 34950
rect 9799 34894 9867 34950
rect 9923 34894 9991 34950
rect 10047 34894 10115 34950
rect 10171 34894 10239 34950
rect 10295 34894 10363 34950
rect 10419 34894 10487 34950
rect 10543 34894 10553 34950
rect 8741 34826 10553 34894
rect 8741 34770 8751 34826
rect 8807 34770 8875 34826
rect 8931 34770 8999 34826
rect 9055 34770 9123 34826
rect 9179 34770 9247 34826
rect 9303 34770 9371 34826
rect 9427 34770 9495 34826
rect 9551 34770 9619 34826
rect 9675 34770 9743 34826
rect 9799 34770 9867 34826
rect 9923 34770 9991 34826
rect 10047 34770 10115 34826
rect 10171 34770 10239 34826
rect 10295 34770 10363 34826
rect 10419 34770 10487 34826
rect 10543 34770 10553 34826
rect 8741 34702 10553 34770
rect 8741 34646 8751 34702
rect 8807 34646 8875 34702
rect 8931 34646 8999 34702
rect 9055 34646 9123 34702
rect 9179 34646 9247 34702
rect 9303 34646 9371 34702
rect 9427 34646 9495 34702
rect 9551 34646 9619 34702
rect 9675 34646 9743 34702
rect 9799 34646 9867 34702
rect 9923 34646 9991 34702
rect 10047 34646 10115 34702
rect 10171 34646 10239 34702
rect 10295 34646 10363 34702
rect 10419 34646 10487 34702
rect 10543 34646 10553 34702
rect 8741 34578 10553 34646
rect 8741 34522 8751 34578
rect 8807 34522 8875 34578
rect 8931 34522 8999 34578
rect 9055 34522 9123 34578
rect 9179 34522 9247 34578
rect 9303 34522 9371 34578
rect 9427 34522 9495 34578
rect 9551 34522 9619 34578
rect 9675 34522 9743 34578
rect 9799 34522 9867 34578
rect 9923 34522 9991 34578
rect 10047 34522 10115 34578
rect 10171 34522 10239 34578
rect 10295 34522 10363 34578
rect 10419 34522 10487 34578
rect 10543 34522 10553 34578
rect 8741 34454 10553 34522
rect 8741 34398 8751 34454
rect 8807 34398 8875 34454
rect 8931 34398 8999 34454
rect 9055 34398 9123 34454
rect 9179 34398 9247 34454
rect 9303 34398 9371 34454
rect 9427 34398 9495 34454
rect 9551 34398 9619 34454
rect 9675 34398 9743 34454
rect 9799 34398 9867 34454
rect 9923 34398 9991 34454
rect 10047 34398 10115 34454
rect 10171 34398 10239 34454
rect 10295 34398 10363 34454
rect 10419 34398 10487 34454
rect 10543 34398 10553 34454
rect 8741 34330 10553 34398
rect 8741 34274 8751 34330
rect 8807 34274 8875 34330
rect 8931 34274 8999 34330
rect 9055 34274 9123 34330
rect 9179 34274 9247 34330
rect 9303 34274 9371 34330
rect 9427 34274 9495 34330
rect 9551 34274 9619 34330
rect 9675 34274 9743 34330
rect 9799 34274 9867 34330
rect 9923 34274 9991 34330
rect 10047 34274 10115 34330
rect 10171 34274 10239 34330
rect 10295 34274 10363 34330
rect 10419 34274 10487 34330
rect 10543 34274 10553 34330
rect 8741 34206 10553 34274
rect 8741 34150 8751 34206
rect 8807 34150 8875 34206
rect 8931 34150 8999 34206
rect 9055 34150 9123 34206
rect 9179 34150 9247 34206
rect 9303 34150 9371 34206
rect 9427 34150 9495 34206
rect 9551 34150 9619 34206
rect 9675 34150 9743 34206
rect 9799 34150 9867 34206
rect 9923 34150 9991 34206
rect 10047 34150 10115 34206
rect 10171 34150 10239 34206
rect 10295 34150 10363 34206
rect 10419 34150 10487 34206
rect 10543 34150 10553 34206
rect 8741 34082 10553 34150
rect 8741 34026 8751 34082
rect 8807 34026 8875 34082
rect 8931 34026 8999 34082
rect 9055 34026 9123 34082
rect 9179 34026 9247 34082
rect 9303 34026 9371 34082
rect 9427 34026 9495 34082
rect 9551 34026 9619 34082
rect 9675 34026 9743 34082
rect 9799 34026 9867 34082
rect 9923 34026 9991 34082
rect 10047 34026 10115 34082
rect 10171 34026 10239 34082
rect 10295 34026 10363 34082
rect 10419 34026 10487 34082
rect 10543 34026 10553 34082
rect 8741 33958 10553 34026
rect 8741 33902 8751 33958
rect 8807 33902 8875 33958
rect 8931 33902 8999 33958
rect 9055 33902 9123 33958
rect 9179 33902 9247 33958
rect 9303 33902 9371 33958
rect 9427 33902 9495 33958
rect 9551 33902 9619 33958
rect 9675 33902 9743 33958
rect 9799 33902 9867 33958
rect 9923 33902 9991 33958
rect 10047 33902 10115 33958
rect 10171 33902 10239 33958
rect 10295 33902 10363 33958
rect 10419 33902 10487 33958
rect 10543 33902 10553 33958
rect 8741 33834 10553 33902
rect 8741 33778 8751 33834
rect 8807 33778 8875 33834
rect 8931 33778 8999 33834
rect 9055 33778 9123 33834
rect 9179 33778 9247 33834
rect 9303 33778 9371 33834
rect 9427 33778 9495 33834
rect 9551 33778 9619 33834
rect 9675 33778 9743 33834
rect 9799 33778 9867 33834
rect 9923 33778 9991 33834
rect 10047 33778 10115 33834
rect 10171 33778 10239 33834
rect 10295 33778 10363 33834
rect 10419 33778 10487 33834
rect 10543 33778 10553 33834
rect 8741 33710 10553 33778
rect 8741 33654 8751 33710
rect 8807 33654 8875 33710
rect 8931 33654 8999 33710
rect 9055 33654 9123 33710
rect 9179 33654 9247 33710
rect 9303 33654 9371 33710
rect 9427 33654 9495 33710
rect 9551 33654 9619 33710
rect 9675 33654 9743 33710
rect 9799 33654 9867 33710
rect 9923 33654 9991 33710
rect 10047 33654 10115 33710
rect 10171 33654 10239 33710
rect 10295 33654 10363 33710
rect 10419 33654 10487 33710
rect 10543 33654 10553 33710
rect 8741 33586 10553 33654
rect 8741 33530 8751 33586
rect 8807 33530 8875 33586
rect 8931 33530 8999 33586
rect 9055 33530 9123 33586
rect 9179 33530 9247 33586
rect 9303 33530 9371 33586
rect 9427 33530 9495 33586
rect 9551 33530 9619 33586
rect 9675 33530 9743 33586
rect 9799 33530 9867 33586
rect 9923 33530 9991 33586
rect 10047 33530 10115 33586
rect 10171 33530 10239 33586
rect 10295 33530 10363 33586
rect 10419 33530 10487 33586
rect 10543 33530 10553 33586
rect 8741 33462 10553 33530
rect 8741 33406 8751 33462
rect 8807 33406 8875 33462
rect 8931 33406 8999 33462
rect 9055 33406 9123 33462
rect 9179 33406 9247 33462
rect 9303 33406 9371 33462
rect 9427 33406 9495 33462
rect 9551 33406 9619 33462
rect 9675 33406 9743 33462
rect 9799 33406 9867 33462
rect 9923 33406 9991 33462
rect 10047 33406 10115 33462
rect 10171 33406 10239 33462
rect 10295 33406 10363 33462
rect 10419 33406 10487 33462
rect 10543 33406 10553 33462
rect 8741 33338 10553 33406
rect 8741 33282 8751 33338
rect 8807 33282 8875 33338
rect 8931 33282 8999 33338
rect 9055 33282 9123 33338
rect 9179 33282 9247 33338
rect 9303 33282 9371 33338
rect 9427 33282 9495 33338
rect 9551 33282 9619 33338
rect 9675 33282 9743 33338
rect 9799 33282 9867 33338
rect 9923 33282 9991 33338
rect 10047 33282 10115 33338
rect 10171 33282 10239 33338
rect 10295 33282 10363 33338
rect 10419 33282 10487 33338
rect 10543 33282 10553 33338
rect 8741 33214 10553 33282
rect 8741 33158 8751 33214
rect 8807 33158 8875 33214
rect 8931 33158 8999 33214
rect 9055 33158 9123 33214
rect 9179 33158 9247 33214
rect 9303 33158 9371 33214
rect 9427 33158 9495 33214
rect 9551 33158 9619 33214
rect 9675 33158 9743 33214
rect 9799 33158 9867 33214
rect 9923 33158 9991 33214
rect 10047 33158 10115 33214
rect 10171 33158 10239 33214
rect 10295 33158 10363 33214
rect 10419 33158 10487 33214
rect 10543 33158 10553 33214
rect 8741 33090 10553 33158
rect 8741 33034 8751 33090
rect 8807 33034 8875 33090
rect 8931 33034 8999 33090
rect 9055 33034 9123 33090
rect 9179 33034 9247 33090
rect 9303 33034 9371 33090
rect 9427 33034 9495 33090
rect 9551 33034 9619 33090
rect 9675 33034 9743 33090
rect 9799 33034 9867 33090
rect 9923 33034 9991 33090
rect 10047 33034 10115 33090
rect 10171 33034 10239 33090
rect 10295 33034 10363 33090
rect 10419 33034 10487 33090
rect 10543 33034 10553 33090
rect 8741 32966 10553 33034
rect 8741 32910 8751 32966
rect 8807 32910 8875 32966
rect 8931 32910 8999 32966
rect 9055 32910 9123 32966
rect 9179 32910 9247 32966
rect 9303 32910 9371 32966
rect 9427 32910 9495 32966
rect 9551 32910 9619 32966
rect 9675 32910 9743 32966
rect 9799 32910 9867 32966
rect 9923 32910 9991 32966
rect 10047 32910 10115 32966
rect 10171 32910 10239 32966
rect 10295 32910 10363 32966
rect 10419 32910 10487 32966
rect 10543 32910 10553 32966
rect 8741 32842 10553 32910
rect 8741 32786 8751 32842
rect 8807 32786 8875 32842
rect 8931 32786 8999 32842
rect 9055 32786 9123 32842
rect 9179 32786 9247 32842
rect 9303 32786 9371 32842
rect 9427 32786 9495 32842
rect 9551 32786 9619 32842
rect 9675 32786 9743 32842
rect 9799 32786 9867 32842
rect 9923 32786 9991 32842
rect 10047 32786 10115 32842
rect 10171 32786 10239 32842
rect 10295 32786 10363 32842
rect 10419 32786 10487 32842
rect 10543 32786 10553 32842
rect 8741 32718 10553 32786
rect 8741 32662 8751 32718
rect 8807 32662 8875 32718
rect 8931 32662 8999 32718
rect 9055 32662 9123 32718
rect 9179 32662 9247 32718
rect 9303 32662 9371 32718
rect 9427 32662 9495 32718
rect 9551 32662 9619 32718
rect 9675 32662 9743 32718
rect 9799 32662 9867 32718
rect 9923 32662 9991 32718
rect 10047 32662 10115 32718
rect 10171 32662 10239 32718
rect 10295 32662 10363 32718
rect 10419 32662 10487 32718
rect 10543 32662 10553 32718
rect 8741 32594 10553 32662
rect 8741 32538 8751 32594
rect 8807 32538 8875 32594
rect 8931 32538 8999 32594
rect 9055 32538 9123 32594
rect 9179 32538 9247 32594
rect 9303 32538 9371 32594
rect 9427 32538 9495 32594
rect 9551 32538 9619 32594
rect 9675 32538 9743 32594
rect 9799 32538 9867 32594
rect 9923 32538 9991 32594
rect 10047 32538 10115 32594
rect 10171 32538 10239 32594
rect 10295 32538 10363 32594
rect 10419 32538 10487 32594
rect 10543 32538 10553 32594
rect 8741 32470 10553 32538
rect 8741 32414 8751 32470
rect 8807 32414 8875 32470
rect 8931 32414 8999 32470
rect 9055 32414 9123 32470
rect 9179 32414 9247 32470
rect 9303 32414 9371 32470
rect 9427 32414 9495 32470
rect 9551 32414 9619 32470
rect 9675 32414 9743 32470
rect 9799 32414 9867 32470
rect 9923 32414 9991 32470
rect 10047 32414 10115 32470
rect 10171 32414 10239 32470
rect 10295 32414 10363 32470
rect 10419 32414 10487 32470
rect 10543 32414 10553 32470
rect 8741 32346 10553 32414
rect 8741 32290 8751 32346
rect 8807 32290 8875 32346
rect 8931 32290 8999 32346
rect 9055 32290 9123 32346
rect 9179 32290 9247 32346
rect 9303 32290 9371 32346
rect 9427 32290 9495 32346
rect 9551 32290 9619 32346
rect 9675 32290 9743 32346
rect 9799 32290 9867 32346
rect 9923 32290 9991 32346
rect 10047 32290 10115 32346
rect 10171 32290 10239 32346
rect 10295 32290 10363 32346
rect 10419 32290 10487 32346
rect 10543 32290 10553 32346
rect 8741 32222 10553 32290
rect 8741 32166 8751 32222
rect 8807 32166 8875 32222
rect 8931 32166 8999 32222
rect 9055 32166 9123 32222
rect 9179 32166 9247 32222
rect 9303 32166 9371 32222
rect 9427 32166 9495 32222
rect 9551 32166 9619 32222
rect 9675 32166 9743 32222
rect 9799 32166 9867 32222
rect 9923 32166 9991 32222
rect 10047 32166 10115 32222
rect 10171 32166 10239 32222
rect 10295 32166 10363 32222
rect 10419 32166 10487 32222
rect 10543 32166 10553 32222
rect 8741 32098 10553 32166
rect 8741 32042 8751 32098
rect 8807 32042 8875 32098
rect 8931 32042 8999 32098
rect 9055 32042 9123 32098
rect 9179 32042 9247 32098
rect 9303 32042 9371 32098
rect 9427 32042 9495 32098
rect 9551 32042 9619 32098
rect 9675 32042 9743 32098
rect 9799 32042 9867 32098
rect 9923 32042 9991 32098
rect 10047 32042 10115 32098
rect 10171 32042 10239 32098
rect 10295 32042 10363 32098
rect 10419 32042 10487 32098
rect 10543 32042 10553 32098
rect 8741 32032 10553 32042
rect 12842 34950 13910 34960
rect 12842 34894 12852 34950
rect 12908 34894 12976 34950
rect 13032 34894 13100 34950
rect 13156 34894 13224 34950
rect 13280 34894 13348 34950
rect 13404 34894 13472 34950
rect 13528 34894 13596 34950
rect 13652 34894 13720 34950
rect 13776 34894 13844 34950
rect 13900 34894 13910 34950
rect 12842 34826 13910 34894
rect 12842 34770 12852 34826
rect 12908 34770 12976 34826
rect 13032 34770 13100 34826
rect 13156 34770 13224 34826
rect 13280 34770 13348 34826
rect 13404 34770 13472 34826
rect 13528 34770 13596 34826
rect 13652 34770 13720 34826
rect 13776 34770 13844 34826
rect 13900 34770 13910 34826
rect 12842 34702 13910 34770
rect 12842 34646 12852 34702
rect 12908 34646 12976 34702
rect 13032 34646 13100 34702
rect 13156 34646 13224 34702
rect 13280 34646 13348 34702
rect 13404 34646 13472 34702
rect 13528 34646 13596 34702
rect 13652 34646 13720 34702
rect 13776 34646 13844 34702
rect 13900 34646 13910 34702
rect 12842 34578 13910 34646
rect 12842 34522 12852 34578
rect 12908 34522 12976 34578
rect 13032 34522 13100 34578
rect 13156 34522 13224 34578
rect 13280 34522 13348 34578
rect 13404 34522 13472 34578
rect 13528 34522 13596 34578
rect 13652 34522 13720 34578
rect 13776 34522 13844 34578
rect 13900 34522 13910 34578
rect 12842 34454 13910 34522
rect 12842 34398 12852 34454
rect 12908 34398 12976 34454
rect 13032 34398 13100 34454
rect 13156 34398 13224 34454
rect 13280 34398 13348 34454
rect 13404 34398 13472 34454
rect 13528 34398 13596 34454
rect 13652 34398 13720 34454
rect 13776 34398 13844 34454
rect 13900 34398 13910 34454
rect 12842 34330 13910 34398
rect 12842 34274 12852 34330
rect 12908 34274 12976 34330
rect 13032 34274 13100 34330
rect 13156 34274 13224 34330
rect 13280 34274 13348 34330
rect 13404 34274 13472 34330
rect 13528 34274 13596 34330
rect 13652 34274 13720 34330
rect 13776 34274 13844 34330
rect 13900 34274 13910 34330
rect 12842 34206 13910 34274
rect 12842 34150 12852 34206
rect 12908 34150 12976 34206
rect 13032 34150 13100 34206
rect 13156 34150 13224 34206
rect 13280 34150 13348 34206
rect 13404 34150 13472 34206
rect 13528 34150 13596 34206
rect 13652 34150 13720 34206
rect 13776 34150 13844 34206
rect 13900 34150 13910 34206
rect 12842 34082 13910 34150
rect 12842 34026 12852 34082
rect 12908 34026 12976 34082
rect 13032 34026 13100 34082
rect 13156 34026 13224 34082
rect 13280 34026 13348 34082
rect 13404 34026 13472 34082
rect 13528 34026 13596 34082
rect 13652 34026 13720 34082
rect 13776 34026 13844 34082
rect 13900 34026 13910 34082
rect 12842 33958 13910 34026
rect 12842 33902 12852 33958
rect 12908 33902 12976 33958
rect 13032 33902 13100 33958
rect 13156 33902 13224 33958
rect 13280 33902 13348 33958
rect 13404 33902 13472 33958
rect 13528 33902 13596 33958
rect 13652 33902 13720 33958
rect 13776 33902 13844 33958
rect 13900 33902 13910 33958
rect 12842 33834 13910 33902
rect 12842 33778 12852 33834
rect 12908 33778 12976 33834
rect 13032 33778 13100 33834
rect 13156 33778 13224 33834
rect 13280 33778 13348 33834
rect 13404 33778 13472 33834
rect 13528 33778 13596 33834
rect 13652 33778 13720 33834
rect 13776 33778 13844 33834
rect 13900 33778 13910 33834
rect 12842 33710 13910 33778
rect 12842 33654 12852 33710
rect 12908 33654 12976 33710
rect 13032 33654 13100 33710
rect 13156 33654 13224 33710
rect 13280 33654 13348 33710
rect 13404 33654 13472 33710
rect 13528 33654 13596 33710
rect 13652 33654 13720 33710
rect 13776 33654 13844 33710
rect 13900 33654 13910 33710
rect 12842 33586 13910 33654
rect 12842 33530 12852 33586
rect 12908 33530 12976 33586
rect 13032 33530 13100 33586
rect 13156 33530 13224 33586
rect 13280 33530 13348 33586
rect 13404 33530 13472 33586
rect 13528 33530 13596 33586
rect 13652 33530 13720 33586
rect 13776 33530 13844 33586
rect 13900 33530 13910 33586
rect 12842 33462 13910 33530
rect 12842 33406 12852 33462
rect 12908 33406 12976 33462
rect 13032 33406 13100 33462
rect 13156 33406 13224 33462
rect 13280 33406 13348 33462
rect 13404 33406 13472 33462
rect 13528 33406 13596 33462
rect 13652 33406 13720 33462
rect 13776 33406 13844 33462
rect 13900 33406 13910 33462
rect 12842 33338 13910 33406
rect 12842 33282 12852 33338
rect 12908 33282 12976 33338
rect 13032 33282 13100 33338
rect 13156 33282 13224 33338
rect 13280 33282 13348 33338
rect 13404 33282 13472 33338
rect 13528 33282 13596 33338
rect 13652 33282 13720 33338
rect 13776 33282 13844 33338
rect 13900 33282 13910 33338
rect 12842 33214 13910 33282
rect 12842 33158 12852 33214
rect 12908 33158 12976 33214
rect 13032 33158 13100 33214
rect 13156 33158 13224 33214
rect 13280 33158 13348 33214
rect 13404 33158 13472 33214
rect 13528 33158 13596 33214
rect 13652 33158 13720 33214
rect 13776 33158 13844 33214
rect 13900 33158 13910 33214
rect 12842 33090 13910 33158
rect 12842 33034 12852 33090
rect 12908 33034 12976 33090
rect 13032 33034 13100 33090
rect 13156 33034 13224 33090
rect 13280 33034 13348 33090
rect 13404 33034 13472 33090
rect 13528 33034 13596 33090
rect 13652 33034 13720 33090
rect 13776 33034 13844 33090
rect 13900 33034 13910 33090
rect 12842 32966 13910 33034
rect 12842 32910 12852 32966
rect 12908 32910 12976 32966
rect 13032 32910 13100 32966
rect 13156 32910 13224 32966
rect 13280 32910 13348 32966
rect 13404 32910 13472 32966
rect 13528 32910 13596 32966
rect 13652 32910 13720 32966
rect 13776 32910 13844 32966
rect 13900 32910 13910 32966
rect 12842 32842 13910 32910
rect 12842 32786 12852 32842
rect 12908 32786 12976 32842
rect 13032 32786 13100 32842
rect 13156 32786 13224 32842
rect 13280 32786 13348 32842
rect 13404 32786 13472 32842
rect 13528 32786 13596 32842
rect 13652 32786 13720 32842
rect 13776 32786 13844 32842
rect 13900 32786 13910 32842
rect 12842 32718 13910 32786
rect 12842 32662 12852 32718
rect 12908 32662 12976 32718
rect 13032 32662 13100 32718
rect 13156 32662 13224 32718
rect 13280 32662 13348 32718
rect 13404 32662 13472 32718
rect 13528 32662 13596 32718
rect 13652 32662 13720 32718
rect 13776 32662 13844 32718
rect 13900 32662 13910 32718
rect 12842 32594 13910 32662
rect 12842 32538 12852 32594
rect 12908 32538 12976 32594
rect 13032 32538 13100 32594
rect 13156 32538 13224 32594
rect 13280 32538 13348 32594
rect 13404 32538 13472 32594
rect 13528 32538 13596 32594
rect 13652 32538 13720 32594
rect 13776 32538 13844 32594
rect 13900 32538 13910 32594
rect 12842 32470 13910 32538
rect 12842 32414 12852 32470
rect 12908 32414 12976 32470
rect 13032 32414 13100 32470
rect 13156 32414 13224 32470
rect 13280 32414 13348 32470
rect 13404 32414 13472 32470
rect 13528 32414 13596 32470
rect 13652 32414 13720 32470
rect 13776 32414 13844 32470
rect 13900 32414 13910 32470
rect 12842 32346 13910 32414
rect 12842 32290 12852 32346
rect 12908 32290 12976 32346
rect 13032 32290 13100 32346
rect 13156 32290 13224 32346
rect 13280 32290 13348 32346
rect 13404 32290 13472 32346
rect 13528 32290 13596 32346
rect 13652 32290 13720 32346
rect 13776 32290 13844 32346
rect 13900 32290 13910 32346
rect 12842 32222 13910 32290
rect 12842 32166 12852 32222
rect 12908 32166 12976 32222
rect 13032 32166 13100 32222
rect 13156 32166 13224 32222
rect 13280 32166 13348 32222
rect 13404 32166 13472 32222
rect 13528 32166 13596 32222
rect 13652 32166 13720 32222
rect 13776 32166 13844 32222
rect 13900 32166 13910 32222
rect 12842 32098 13910 32166
rect 12842 32042 12852 32098
rect 12908 32042 12976 32098
rect 13032 32042 13100 32098
rect 13156 32042 13224 32098
rect 13280 32042 13348 32098
rect 13404 32042 13472 32098
rect 13528 32042 13596 32098
rect 13652 32042 13720 32098
rect 13776 32042 13844 32098
rect 13900 32042 13910 32098
rect 12842 32032 13910 32042
rect 4129 32003 4205 32013
rect 2013 31906 2089 31974
rect 2013 31850 2023 31906
rect 2079 31850 2089 31906
rect 2013 31782 2089 31850
rect 2013 31726 2023 31782
rect 2079 31726 2089 31782
rect 2013 31658 2089 31726
rect 2013 31602 2023 31658
rect 2079 31602 2089 31658
rect 2013 31534 2089 31602
rect 2013 31478 2023 31534
rect 2079 31478 2089 31534
rect 2013 31410 2089 31478
rect 2013 31354 2023 31410
rect 2079 31354 2089 31410
rect 2013 31286 2089 31354
rect 2013 31230 2023 31286
rect 2079 31230 2089 31286
rect 2013 31162 2089 31230
rect 2013 31106 2023 31162
rect 2079 31106 2089 31162
rect 2013 31038 2089 31106
rect 2013 30982 2023 31038
rect 2079 30982 2089 31038
rect 2013 30914 2089 30982
rect 2013 30858 2023 30914
rect 2079 30858 2089 30914
rect 2013 30790 2089 30858
rect 2013 30734 2023 30790
rect 2079 30734 2089 30790
rect 2013 30666 2089 30734
rect 2013 30610 2023 30666
rect 2079 30610 2089 30666
rect 2013 30542 2089 30610
rect 2013 30486 2023 30542
rect 2079 30486 2089 30542
rect 2013 30418 2089 30486
rect 2013 30362 2023 30418
rect 2079 30362 2089 30418
rect 2013 30294 2089 30362
rect 2013 30238 2023 30294
rect 2079 30238 2089 30294
rect 2013 30170 2089 30238
rect 2013 30114 2023 30170
rect 2079 30114 2089 30170
rect 2013 30046 2089 30114
rect 2013 29990 2023 30046
rect 2079 29990 2089 30046
rect 2013 29922 2089 29990
rect 2013 29866 2023 29922
rect 2079 29866 2089 29922
rect 2013 29798 2089 29866
rect 2013 29742 2023 29798
rect 2079 29742 2089 29798
rect 2013 29674 2089 29742
rect 2013 29618 2023 29674
rect 2079 29618 2089 29674
rect 2013 29550 2089 29618
rect 2013 29494 2023 29550
rect 2079 29494 2089 29550
rect 2013 29426 2089 29494
rect 2013 29370 2023 29426
rect 2079 29370 2089 29426
rect 2013 29302 2089 29370
rect 2013 29246 2023 29302
rect 2079 29246 2089 29302
rect 2013 29178 2089 29246
rect 2013 29122 2023 29178
rect 2079 29122 2089 29178
rect 2013 29054 2089 29122
rect 2013 28998 2023 29054
rect 2079 28998 2089 29054
rect 1365 28879 1375 28935
rect 1431 28879 1441 28935
rect 1365 28811 1441 28879
rect 1365 28755 1375 28811
rect 1431 28755 1441 28811
rect 1365 28687 1441 28755
rect 1365 28631 1375 28687
rect 1431 28631 1441 28687
rect 1365 28563 1441 28631
rect 1365 28507 1375 28563
rect 1431 28507 1441 28563
rect 1365 28439 1441 28507
rect 1365 28383 1375 28439
rect 1431 28383 1441 28439
rect 1365 28315 1441 28383
rect 1365 28259 1375 28315
rect 1431 28259 1441 28315
rect 1365 28191 1441 28259
rect 1365 28135 1375 28191
rect 1431 28135 1441 28191
rect 1365 28067 1441 28135
rect 1365 28011 1375 28067
rect 1431 28011 1441 28067
rect 1365 27943 1441 28011
rect 1365 27887 1375 27943
rect 1431 27887 1441 27943
rect 1365 27819 1441 27887
rect 1365 27763 1375 27819
rect 1431 27763 1441 27819
rect 1365 27695 1441 27763
rect 1365 27639 1375 27695
rect 1431 27639 1441 27695
rect 1365 27571 1441 27639
rect 1365 27515 1375 27571
rect 1431 27515 1441 27571
rect 1365 27447 1441 27515
rect 1365 27391 1375 27447
rect 1431 27391 1441 27447
rect 1365 27323 1441 27391
rect 1365 27267 1375 27323
rect 1431 27267 1441 27323
rect 1365 27257 1441 27267
rect 1489 28922 1565 28932
rect 1489 28866 1499 28922
rect 1555 28866 1565 28922
rect 1489 28798 1565 28866
rect 2013 28930 2089 28998
rect 2013 28874 2023 28930
rect 2079 28874 2089 28930
rect 2013 28864 2089 28874
rect 4425 31750 6237 31760
rect 4425 31694 4435 31750
rect 4491 31694 4559 31750
rect 4615 31694 4683 31750
rect 4739 31694 4807 31750
rect 4863 31694 4931 31750
rect 4987 31694 5055 31750
rect 5111 31694 5179 31750
rect 5235 31694 5303 31750
rect 5359 31694 5427 31750
rect 5483 31694 5551 31750
rect 5607 31694 5675 31750
rect 5731 31694 5799 31750
rect 5855 31694 5923 31750
rect 5979 31694 6047 31750
rect 6103 31694 6171 31750
rect 6227 31694 6237 31750
rect 4425 31626 6237 31694
rect 4425 31570 4435 31626
rect 4491 31570 4559 31626
rect 4615 31570 4683 31626
rect 4739 31570 4807 31626
rect 4863 31570 4931 31626
rect 4987 31570 5055 31626
rect 5111 31570 5179 31626
rect 5235 31570 5303 31626
rect 5359 31570 5427 31626
rect 5483 31570 5551 31626
rect 5607 31570 5675 31626
rect 5731 31570 5799 31626
rect 5855 31570 5923 31626
rect 5979 31570 6047 31626
rect 6103 31570 6171 31626
rect 6227 31570 6237 31626
rect 4425 31502 6237 31570
rect 4425 31446 4435 31502
rect 4491 31446 4559 31502
rect 4615 31446 4683 31502
rect 4739 31446 4807 31502
rect 4863 31446 4931 31502
rect 4987 31446 5055 31502
rect 5111 31446 5179 31502
rect 5235 31446 5303 31502
rect 5359 31446 5427 31502
rect 5483 31446 5551 31502
rect 5607 31446 5675 31502
rect 5731 31446 5799 31502
rect 5855 31446 5923 31502
rect 5979 31446 6047 31502
rect 6103 31446 6171 31502
rect 6227 31446 6237 31502
rect 4425 31378 6237 31446
rect 4425 31322 4435 31378
rect 4491 31322 4559 31378
rect 4615 31322 4683 31378
rect 4739 31322 4807 31378
rect 4863 31322 4931 31378
rect 4987 31322 5055 31378
rect 5111 31322 5179 31378
rect 5235 31322 5303 31378
rect 5359 31322 5427 31378
rect 5483 31322 5551 31378
rect 5607 31322 5675 31378
rect 5731 31322 5799 31378
rect 5855 31322 5923 31378
rect 5979 31322 6047 31378
rect 6103 31322 6171 31378
rect 6227 31322 6237 31378
rect 4425 31254 6237 31322
rect 4425 31198 4435 31254
rect 4491 31198 4559 31254
rect 4615 31198 4683 31254
rect 4739 31198 4807 31254
rect 4863 31198 4931 31254
rect 4987 31198 5055 31254
rect 5111 31198 5179 31254
rect 5235 31198 5303 31254
rect 5359 31198 5427 31254
rect 5483 31198 5551 31254
rect 5607 31198 5675 31254
rect 5731 31198 5799 31254
rect 5855 31198 5923 31254
rect 5979 31198 6047 31254
rect 6103 31198 6171 31254
rect 6227 31198 6237 31254
rect 4425 31130 6237 31198
rect 4425 31074 4435 31130
rect 4491 31074 4559 31130
rect 4615 31074 4683 31130
rect 4739 31074 4807 31130
rect 4863 31074 4931 31130
rect 4987 31074 5055 31130
rect 5111 31074 5179 31130
rect 5235 31074 5303 31130
rect 5359 31074 5427 31130
rect 5483 31074 5551 31130
rect 5607 31074 5675 31130
rect 5731 31074 5799 31130
rect 5855 31074 5923 31130
rect 5979 31074 6047 31130
rect 6103 31074 6171 31130
rect 6227 31074 6237 31130
rect 4425 31006 6237 31074
rect 4425 30950 4435 31006
rect 4491 30950 4559 31006
rect 4615 30950 4683 31006
rect 4739 30950 4807 31006
rect 4863 30950 4931 31006
rect 4987 30950 5055 31006
rect 5111 30950 5179 31006
rect 5235 30950 5303 31006
rect 5359 30950 5427 31006
rect 5483 30950 5551 31006
rect 5607 30950 5675 31006
rect 5731 30950 5799 31006
rect 5855 30950 5923 31006
rect 5979 30950 6047 31006
rect 6103 30950 6171 31006
rect 6227 30950 6237 31006
rect 4425 30882 6237 30950
rect 4425 30826 4435 30882
rect 4491 30826 4559 30882
rect 4615 30826 4683 30882
rect 4739 30826 4807 30882
rect 4863 30826 4931 30882
rect 4987 30826 5055 30882
rect 5111 30826 5179 30882
rect 5235 30826 5303 30882
rect 5359 30826 5427 30882
rect 5483 30826 5551 30882
rect 5607 30826 5675 30882
rect 5731 30826 5799 30882
rect 5855 30826 5923 30882
rect 5979 30826 6047 30882
rect 6103 30826 6171 30882
rect 6227 30826 6237 30882
rect 4425 30758 6237 30826
rect 4425 30702 4435 30758
rect 4491 30702 4559 30758
rect 4615 30702 4683 30758
rect 4739 30702 4807 30758
rect 4863 30702 4931 30758
rect 4987 30702 5055 30758
rect 5111 30702 5179 30758
rect 5235 30702 5303 30758
rect 5359 30702 5427 30758
rect 5483 30702 5551 30758
rect 5607 30702 5675 30758
rect 5731 30702 5799 30758
rect 5855 30702 5923 30758
rect 5979 30702 6047 30758
rect 6103 30702 6171 30758
rect 6227 30702 6237 30758
rect 4425 30634 6237 30702
rect 4425 30578 4435 30634
rect 4491 30578 4559 30634
rect 4615 30578 4683 30634
rect 4739 30578 4807 30634
rect 4863 30578 4931 30634
rect 4987 30578 5055 30634
rect 5111 30578 5179 30634
rect 5235 30578 5303 30634
rect 5359 30578 5427 30634
rect 5483 30578 5551 30634
rect 5607 30578 5675 30634
rect 5731 30578 5799 30634
rect 5855 30578 5923 30634
rect 5979 30578 6047 30634
rect 6103 30578 6171 30634
rect 6227 30578 6237 30634
rect 4425 30510 6237 30578
rect 4425 30454 4435 30510
rect 4491 30454 4559 30510
rect 4615 30454 4683 30510
rect 4739 30454 4807 30510
rect 4863 30454 4931 30510
rect 4987 30454 5055 30510
rect 5111 30454 5179 30510
rect 5235 30454 5303 30510
rect 5359 30454 5427 30510
rect 5483 30454 5551 30510
rect 5607 30454 5675 30510
rect 5731 30454 5799 30510
rect 5855 30454 5923 30510
rect 5979 30454 6047 30510
rect 6103 30454 6171 30510
rect 6227 30454 6237 30510
rect 4425 30386 6237 30454
rect 4425 30330 4435 30386
rect 4491 30330 4559 30386
rect 4615 30330 4683 30386
rect 4739 30330 4807 30386
rect 4863 30330 4931 30386
rect 4987 30330 5055 30386
rect 5111 30330 5179 30386
rect 5235 30330 5303 30386
rect 5359 30330 5427 30386
rect 5483 30330 5551 30386
rect 5607 30330 5675 30386
rect 5731 30330 5799 30386
rect 5855 30330 5923 30386
rect 5979 30330 6047 30386
rect 6103 30330 6171 30386
rect 6227 30330 6237 30386
rect 4425 30262 6237 30330
rect 4425 30206 4435 30262
rect 4491 30206 4559 30262
rect 4615 30206 4683 30262
rect 4739 30206 4807 30262
rect 4863 30206 4931 30262
rect 4987 30206 5055 30262
rect 5111 30206 5179 30262
rect 5235 30206 5303 30262
rect 5359 30206 5427 30262
rect 5483 30206 5551 30262
rect 5607 30206 5675 30262
rect 5731 30206 5799 30262
rect 5855 30206 5923 30262
rect 5979 30206 6047 30262
rect 6103 30206 6171 30262
rect 6227 30206 6237 30262
rect 4425 30138 6237 30206
rect 4425 30082 4435 30138
rect 4491 30082 4559 30138
rect 4615 30082 4683 30138
rect 4739 30082 4807 30138
rect 4863 30082 4931 30138
rect 4987 30082 5055 30138
rect 5111 30082 5179 30138
rect 5235 30082 5303 30138
rect 5359 30082 5427 30138
rect 5483 30082 5551 30138
rect 5607 30082 5675 30138
rect 5731 30082 5799 30138
rect 5855 30082 5923 30138
rect 5979 30082 6047 30138
rect 6103 30082 6171 30138
rect 6227 30082 6237 30138
rect 4425 30014 6237 30082
rect 4425 29958 4435 30014
rect 4491 29958 4559 30014
rect 4615 29958 4683 30014
rect 4739 29958 4807 30014
rect 4863 29958 4931 30014
rect 4987 29958 5055 30014
rect 5111 29958 5179 30014
rect 5235 29958 5303 30014
rect 5359 29958 5427 30014
rect 5483 29958 5551 30014
rect 5607 29958 5675 30014
rect 5731 29958 5799 30014
rect 5855 29958 5923 30014
rect 5979 29958 6047 30014
rect 6103 29958 6171 30014
rect 6227 29958 6237 30014
rect 4425 29890 6237 29958
rect 4425 29834 4435 29890
rect 4491 29834 4559 29890
rect 4615 29834 4683 29890
rect 4739 29834 4807 29890
rect 4863 29834 4931 29890
rect 4987 29834 5055 29890
rect 5111 29834 5179 29890
rect 5235 29834 5303 29890
rect 5359 29834 5427 29890
rect 5483 29834 5551 29890
rect 5607 29834 5675 29890
rect 5731 29834 5799 29890
rect 5855 29834 5923 29890
rect 5979 29834 6047 29890
rect 6103 29834 6171 29890
rect 6227 29834 6237 29890
rect 4425 29766 6237 29834
rect 4425 29710 4435 29766
rect 4491 29710 4559 29766
rect 4615 29710 4683 29766
rect 4739 29710 4807 29766
rect 4863 29710 4931 29766
rect 4987 29710 5055 29766
rect 5111 29710 5179 29766
rect 5235 29710 5303 29766
rect 5359 29710 5427 29766
rect 5483 29710 5551 29766
rect 5607 29710 5675 29766
rect 5731 29710 5799 29766
rect 5855 29710 5923 29766
rect 5979 29710 6047 29766
rect 6103 29710 6171 29766
rect 6227 29710 6237 29766
rect 4425 29642 6237 29710
rect 4425 29586 4435 29642
rect 4491 29586 4559 29642
rect 4615 29586 4683 29642
rect 4739 29586 4807 29642
rect 4863 29586 4931 29642
rect 4987 29586 5055 29642
rect 5111 29586 5179 29642
rect 5235 29586 5303 29642
rect 5359 29586 5427 29642
rect 5483 29586 5551 29642
rect 5607 29586 5675 29642
rect 5731 29586 5799 29642
rect 5855 29586 5923 29642
rect 5979 29586 6047 29642
rect 6103 29586 6171 29642
rect 6227 29586 6237 29642
rect 4425 29518 6237 29586
rect 4425 29462 4435 29518
rect 4491 29462 4559 29518
rect 4615 29462 4683 29518
rect 4739 29462 4807 29518
rect 4863 29462 4931 29518
rect 4987 29462 5055 29518
rect 5111 29462 5179 29518
rect 5235 29462 5303 29518
rect 5359 29462 5427 29518
rect 5483 29462 5551 29518
rect 5607 29462 5675 29518
rect 5731 29462 5799 29518
rect 5855 29462 5923 29518
rect 5979 29462 6047 29518
rect 6103 29462 6171 29518
rect 6227 29462 6237 29518
rect 4425 29394 6237 29462
rect 4425 29338 4435 29394
rect 4491 29338 4559 29394
rect 4615 29338 4683 29394
rect 4739 29338 4807 29394
rect 4863 29338 4931 29394
rect 4987 29338 5055 29394
rect 5111 29338 5179 29394
rect 5235 29338 5303 29394
rect 5359 29338 5427 29394
rect 5483 29338 5551 29394
rect 5607 29338 5675 29394
rect 5731 29338 5799 29394
rect 5855 29338 5923 29394
rect 5979 29338 6047 29394
rect 6103 29338 6171 29394
rect 6227 29338 6237 29394
rect 4425 29270 6237 29338
rect 4425 29214 4435 29270
rect 4491 29214 4559 29270
rect 4615 29214 4683 29270
rect 4739 29214 4807 29270
rect 4863 29214 4931 29270
rect 4987 29214 5055 29270
rect 5111 29214 5179 29270
rect 5235 29214 5303 29270
rect 5359 29214 5427 29270
rect 5483 29214 5551 29270
rect 5607 29214 5675 29270
rect 5731 29214 5799 29270
rect 5855 29214 5923 29270
rect 5979 29214 6047 29270
rect 6103 29214 6171 29270
rect 6227 29214 6237 29270
rect 4425 29146 6237 29214
rect 4425 29090 4435 29146
rect 4491 29090 4559 29146
rect 4615 29090 4683 29146
rect 4739 29090 4807 29146
rect 4863 29090 4931 29146
rect 4987 29090 5055 29146
rect 5111 29090 5179 29146
rect 5235 29090 5303 29146
rect 5359 29090 5427 29146
rect 5483 29090 5551 29146
rect 5607 29090 5675 29146
rect 5731 29090 5799 29146
rect 5855 29090 5923 29146
rect 5979 29090 6047 29146
rect 6103 29090 6171 29146
rect 6227 29090 6237 29146
rect 4425 29022 6237 29090
rect 4425 28966 4435 29022
rect 4491 28966 4559 29022
rect 4615 28966 4683 29022
rect 4739 28966 4807 29022
rect 4863 28966 4931 29022
rect 4987 28966 5055 29022
rect 5111 28966 5179 29022
rect 5235 28966 5303 29022
rect 5359 28966 5427 29022
rect 5483 28966 5551 29022
rect 5607 28966 5675 29022
rect 5731 28966 5799 29022
rect 5855 28966 5923 29022
rect 5979 28966 6047 29022
rect 6103 28966 6171 29022
rect 6227 28966 6237 29022
rect 4425 28898 6237 28966
rect 4425 28842 4435 28898
rect 4491 28842 4559 28898
rect 4615 28842 4683 28898
rect 4739 28842 4807 28898
rect 4863 28842 4931 28898
rect 4987 28842 5055 28898
rect 5111 28842 5179 28898
rect 5235 28842 5303 28898
rect 5359 28842 5427 28898
rect 5483 28842 5551 28898
rect 5607 28842 5675 28898
rect 5731 28842 5799 28898
rect 5855 28842 5923 28898
rect 5979 28842 6047 28898
rect 6103 28842 6171 28898
rect 6227 28842 6237 28898
rect 4425 28832 6237 28842
rect 7552 31750 8620 31760
rect 7552 31694 7562 31750
rect 7618 31694 7686 31750
rect 7742 31694 7810 31750
rect 7866 31694 7934 31750
rect 7990 31694 8058 31750
rect 8114 31694 8182 31750
rect 8238 31694 8306 31750
rect 8362 31694 8430 31750
rect 8486 31694 8554 31750
rect 8610 31694 8620 31750
rect 7552 31626 8620 31694
rect 7552 31570 7562 31626
rect 7618 31570 7686 31626
rect 7742 31570 7810 31626
rect 7866 31570 7934 31626
rect 7990 31570 8058 31626
rect 8114 31570 8182 31626
rect 8238 31570 8306 31626
rect 8362 31570 8430 31626
rect 8486 31570 8554 31626
rect 8610 31570 8620 31626
rect 7552 31502 8620 31570
rect 7552 31446 7562 31502
rect 7618 31446 7686 31502
rect 7742 31446 7810 31502
rect 7866 31446 7934 31502
rect 7990 31446 8058 31502
rect 8114 31446 8182 31502
rect 8238 31446 8306 31502
rect 8362 31446 8430 31502
rect 8486 31446 8554 31502
rect 8610 31446 8620 31502
rect 7552 31378 8620 31446
rect 7552 31322 7562 31378
rect 7618 31322 7686 31378
rect 7742 31322 7810 31378
rect 7866 31322 7934 31378
rect 7990 31322 8058 31378
rect 8114 31322 8182 31378
rect 8238 31322 8306 31378
rect 8362 31322 8430 31378
rect 8486 31322 8554 31378
rect 8610 31322 8620 31378
rect 7552 31254 8620 31322
rect 7552 31198 7562 31254
rect 7618 31198 7686 31254
rect 7742 31198 7810 31254
rect 7866 31198 7934 31254
rect 7990 31198 8058 31254
rect 8114 31198 8182 31254
rect 8238 31198 8306 31254
rect 8362 31198 8430 31254
rect 8486 31198 8554 31254
rect 8610 31198 8620 31254
rect 7552 31130 8620 31198
rect 7552 31074 7562 31130
rect 7618 31074 7686 31130
rect 7742 31074 7810 31130
rect 7866 31074 7934 31130
rect 7990 31074 8058 31130
rect 8114 31074 8182 31130
rect 8238 31074 8306 31130
rect 8362 31074 8430 31130
rect 8486 31074 8554 31130
rect 8610 31074 8620 31130
rect 7552 31006 8620 31074
rect 7552 30950 7562 31006
rect 7618 30950 7686 31006
rect 7742 30950 7810 31006
rect 7866 30950 7934 31006
rect 7990 30950 8058 31006
rect 8114 30950 8182 31006
rect 8238 30950 8306 31006
rect 8362 30950 8430 31006
rect 8486 30950 8554 31006
rect 8610 30950 8620 31006
rect 7552 30882 8620 30950
rect 7552 30826 7562 30882
rect 7618 30826 7686 30882
rect 7742 30826 7810 30882
rect 7866 30826 7934 30882
rect 7990 30826 8058 30882
rect 8114 30826 8182 30882
rect 8238 30826 8306 30882
rect 8362 30826 8430 30882
rect 8486 30826 8554 30882
rect 8610 30826 8620 30882
rect 7552 30758 8620 30826
rect 7552 30702 7562 30758
rect 7618 30702 7686 30758
rect 7742 30702 7810 30758
rect 7866 30702 7934 30758
rect 7990 30702 8058 30758
rect 8114 30702 8182 30758
rect 8238 30702 8306 30758
rect 8362 30702 8430 30758
rect 8486 30702 8554 30758
rect 8610 30702 8620 30758
rect 7552 30634 8620 30702
rect 7552 30578 7562 30634
rect 7618 30578 7686 30634
rect 7742 30578 7810 30634
rect 7866 30578 7934 30634
rect 7990 30578 8058 30634
rect 8114 30578 8182 30634
rect 8238 30578 8306 30634
rect 8362 30578 8430 30634
rect 8486 30578 8554 30634
rect 8610 30578 8620 30634
rect 7552 30510 8620 30578
rect 7552 30454 7562 30510
rect 7618 30454 7686 30510
rect 7742 30454 7810 30510
rect 7866 30454 7934 30510
rect 7990 30454 8058 30510
rect 8114 30454 8182 30510
rect 8238 30454 8306 30510
rect 8362 30454 8430 30510
rect 8486 30454 8554 30510
rect 8610 30454 8620 30510
rect 7552 30386 8620 30454
rect 7552 30330 7562 30386
rect 7618 30330 7686 30386
rect 7742 30330 7810 30386
rect 7866 30330 7934 30386
rect 7990 30330 8058 30386
rect 8114 30330 8182 30386
rect 8238 30330 8306 30386
rect 8362 30330 8430 30386
rect 8486 30330 8554 30386
rect 8610 30330 8620 30386
rect 7552 30262 8620 30330
rect 7552 30206 7562 30262
rect 7618 30206 7686 30262
rect 7742 30206 7810 30262
rect 7866 30206 7934 30262
rect 7990 30206 8058 30262
rect 8114 30206 8182 30262
rect 8238 30206 8306 30262
rect 8362 30206 8430 30262
rect 8486 30206 8554 30262
rect 8610 30206 8620 30262
rect 7552 30138 8620 30206
rect 7552 30082 7562 30138
rect 7618 30082 7686 30138
rect 7742 30082 7810 30138
rect 7866 30082 7934 30138
rect 7990 30082 8058 30138
rect 8114 30082 8182 30138
rect 8238 30082 8306 30138
rect 8362 30082 8430 30138
rect 8486 30082 8554 30138
rect 8610 30082 8620 30138
rect 7552 30014 8620 30082
rect 7552 29958 7562 30014
rect 7618 29958 7686 30014
rect 7742 29958 7810 30014
rect 7866 29958 7934 30014
rect 7990 29958 8058 30014
rect 8114 29958 8182 30014
rect 8238 29958 8306 30014
rect 8362 29958 8430 30014
rect 8486 29958 8554 30014
rect 8610 29958 8620 30014
rect 7552 29890 8620 29958
rect 7552 29834 7562 29890
rect 7618 29834 7686 29890
rect 7742 29834 7810 29890
rect 7866 29834 7934 29890
rect 7990 29834 8058 29890
rect 8114 29834 8182 29890
rect 8238 29834 8306 29890
rect 8362 29834 8430 29890
rect 8486 29834 8554 29890
rect 8610 29834 8620 29890
rect 7552 29766 8620 29834
rect 7552 29710 7562 29766
rect 7618 29710 7686 29766
rect 7742 29710 7810 29766
rect 7866 29710 7934 29766
rect 7990 29710 8058 29766
rect 8114 29710 8182 29766
rect 8238 29710 8306 29766
rect 8362 29710 8430 29766
rect 8486 29710 8554 29766
rect 8610 29710 8620 29766
rect 7552 29642 8620 29710
rect 7552 29586 7562 29642
rect 7618 29586 7686 29642
rect 7742 29586 7810 29642
rect 7866 29586 7934 29642
rect 7990 29586 8058 29642
rect 8114 29586 8182 29642
rect 8238 29586 8306 29642
rect 8362 29586 8430 29642
rect 8486 29586 8554 29642
rect 8610 29586 8620 29642
rect 7552 29518 8620 29586
rect 7552 29462 7562 29518
rect 7618 29462 7686 29518
rect 7742 29462 7810 29518
rect 7866 29462 7934 29518
rect 7990 29462 8058 29518
rect 8114 29462 8182 29518
rect 8238 29462 8306 29518
rect 8362 29462 8430 29518
rect 8486 29462 8554 29518
rect 8610 29462 8620 29518
rect 7552 29394 8620 29462
rect 7552 29338 7562 29394
rect 7618 29338 7686 29394
rect 7742 29338 7810 29394
rect 7866 29338 7934 29394
rect 7990 29338 8058 29394
rect 8114 29338 8182 29394
rect 8238 29338 8306 29394
rect 8362 29338 8430 29394
rect 8486 29338 8554 29394
rect 8610 29338 8620 29394
rect 7552 29270 8620 29338
rect 7552 29214 7562 29270
rect 7618 29214 7686 29270
rect 7742 29214 7810 29270
rect 7866 29214 7934 29270
rect 7990 29214 8058 29270
rect 8114 29214 8182 29270
rect 8238 29214 8306 29270
rect 8362 29214 8430 29270
rect 8486 29214 8554 29270
rect 8610 29214 8620 29270
rect 7552 29146 8620 29214
rect 7552 29090 7562 29146
rect 7618 29090 7686 29146
rect 7742 29090 7810 29146
rect 7866 29090 7934 29146
rect 7990 29090 8058 29146
rect 8114 29090 8182 29146
rect 8238 29090 8306 29146
rect 8362 29090 8430 29146
rect 8486 29090 8554 29146
rect 8610 29090 8620 29146
rect 7552 29022 8620 29090
rect 7552 28966 7562 29022
rect 7618 28966 7686 29022
rect 7742 28966 7810 29022
rect 7866 28966 7934 29022
rect 7990 28966 8058 29022
rect 8114 28966 8182 29022
rect 8238 28966 8306 29022
rect 8362 28966 8430 29022
rect 8486 28966 8554 29022
rect 8610 28966 8620 29022
rect 7552 28898 8620 28966
rect 7552 28842 7562 28898
rect 7618 28842 7686 28898
rect 7742 28842 7810 28898
rect 7866 28842 7934 28898
rect 7990 28842 8058 28898
rect 8114 28842 8182 28898
rect 8238 28842 8306 28898
rect 8362 28842 8430 28898
rect 8486 28842 8554 28898
rect 8610 28842 8620 28898
rect 7552 28832 8620 28842
rect 10669 31750 12481 31760
rect 10669 31694 10679 31750
rect 10735 31694 10803 31750
rect 10859 31694 10927 31750
rect 10983 31694 11051 31750
rect 11107 31694 11175 31750
rect 11231 31694 11299 31750
rect 11355 31694 11423 31750
rect 11479 31694 11547 31750
rect 11603 31694 11671 31750
rect 11727 31694 11795 31750
rect 11851 31694 11919 31750
rect 11975 31694 12043 31750
rect 12099 31694 12167 31750
rect 12223 31694 12291 31750
rect 12347 31694 12415 31750
rect 12471 31694 12481 31750
rect 10669 31626 12481 31694
rect 10669 31570 10679 31626
rect 10735 31570 10803 31626
rect 10859 31570 10927 31626
rect 10983 31570 11051 31626
rect 11107 31570 11175 31626
rect 11231 31570 11299 31626
rect 11355 31570 11423 31626
rect 11479 31570 11547 31626
rect 11603 31570 11671 31626
rect 11727 31570 11795 31626
rect 11851 31570 11919 31626
rect 11975 31570 12043 31626
rect 12099 31570 12167 31626
rect 12223 31570 12291 31626
rect 12347 31570 12415 31626
rect 12471 31570 12481 31626
rect 10669 31502 12481 31570
rect 10669 31446 10679 31502
rect 10735 31446 10803 31502
rect 10859 31446 10927 31502
rect 10983 31446 11051 31502
rect 11107 31446 11175 31502
rect 11231 31446 11299 31502
rect 11355 31446 11423 31502
rect 11479 31446 11547 31502
rect 11603 31446 11671 31502
rect 11727 31446 11795 31502
rect 11851 31446 11919 31502
rect 11975 31446 12043 31502
rect 12099 31446 12167 31502
rect 12223 31446 12291 31502
rect 12347 31446 12415 31502
rect 12471 31446 12481 31502
rect 10669 31378 12481 31446
rect 10669 31322 10679 31378
rect 10735 31322 10803 31378
rect 10859 31322 10927 31378
rect 10983 31322 11051 31378
rect 11107 31322 11175 31378
rect 11231 31322 11299 31378
rect 11355 31322 11423 31378
rect 11479 31322 11547 31378
rect 11603 31322 11671 31378
rect 11727 31322 11795 31378
rect 11851 31322 11919 31378
rect 11975 31322 12043 31378
rect 12099 31322 12167 31378
rect 12223 31322 12291 31378
rect 12347 31322 12415 31378
rect 12471 31322 12481 31378
rect 10669 31254 12481 31322
rect 10669 31198 10679 31254
rect 10735 31198 10803 31254
rect 10859 31198 10927 31254
rect 10983 31198 11051 31254
rect 11107 31198 11175 31254
rect 11231 31198 11299 31254
rect 11355 31198 11423 31254
rect 11479 31198 11547 31254
rect 11603 31198 11671 31254
rect 11727 31198 11795 31254
rect 11851 31198 11919 31254
rect 11975 31198 12043 31254
rect 12099 31198 12167 31254
rect 12223 31198 12291 31254
rect 12347 31198 12415 31254
rect 12471 31198 12481 31254
rect 10669 31130 12481 31198
rect 10669 31074 10679 31130
rect 10735 31074 10803 31130
rect 10859 31074 10927 31130
rect 10983 31074 11051 31130
rect 11107 31074 11175 31130
rect 11231 31074 11299 31130
rect 11355 31074 11423 31130
rect 11479 31074 11547 31130
rect 11603 31074 11671 31130
rect 11727 31074 11795 31130
rect 11851 31074 11919 31130
rect 11975 31074 12043 31130
rect 12099 31074 12167 31130
rect 12223 31074 12291 31130
rect 12347 31074 12415 31130
rect 12471 31074 12481 31130
rect 10669 31006 12481 31074
rect 10669 30950 10679 31006
rect 10735 30950 10803 31006
rect 10859 30950 10927 31006
rect 10983 30950 11051 31006
rect 11107 30950 11175 31006
rect 11231 30950 11299 31006
rect 11355 30950 11423 31006
rect 11479 30950 11547 31006
rect 11603 30950 11671 31006
rect 11727 30950 11795 31006
rect 11851 30950 11919 31006
rect 11975 30950 12043 31006
rect 12099 30950 12167 31006
rect 12223 30950 12291 31006
rect 12347 30950 12415 31006
rect 12471 30950 12481 31006
rect 10669 30882 12481 30950
rect 10669 30826 10679 30882
rect 10735 30826 10803 30882
rect 10859 30826 10927 30882
rect 10983 30826 11051 30882
rect 11107 30826 11175 30882
rect 11231 30826 11299 30882
rect 11355 30826 11423 30882
rect 11479 30826 11547 30882
rect 11603 30826 11671 30882
rect 11727 30826 11795 30882
rect 11851 30826 11919 30882
rect 11975 30826 12043 30882
rect 12099 30826 12167 30882
rect 12223 30826 12291 30882
rect 12347 30826 12415 30882
rect 12471 30826 12481 30882
rect 10669 30758 12481 30826
rect 10669 30702 10679 30758
rect 10735 30702 10803 30758
rect 10859 30702 10927 30758
rect 10983 30702 11051 30758
rect 11107 30702 11175 30758
rect 11231 30702 11299 30758
rect 11355 30702 11423 30758
rect 11479 30702 11547 30758
rect 11603 30702 11671 30758
rect 11727 30702 11795 30758
rect 11851 30702 11919 30758
rect 11975 30702 12043 30758
rect 12099 30702 12167 30758
rect 12223 30702 12291 30758
rect 12347 30702 12415 30758
rect 12471 30702 12481 30758
rect 10669 30634 12481 30702
rect 10669 30578 10679 30634
rect 10735 30578 10803 30634
rect 10859 30578 10927 30634
rect 10983 30578 11051 30634
rect 11107 30578 11175 30634
rect 11231 30578 11299 30634
rect 11355 30578 11423 30634
rect 11479 30578 11547 30634
rect 11603 30578 11671 30634
rect 11727 30578 11795 30634
rect 11851 30578 11919 30634
rect 11975 30578 12043 30634
rect 12099 30578 12167 30634
rect 12223 30578 12291 30634
rect 12347 30578 12415 30634
rect 12471 30578 12481 30634
rect 10669 30510 12481 30578
rect 10669 30454 10679 30510
rect 10735 30454 10803 30510
rect 10859 30454 10927 30510
rect 10983 30454 11051 30510
rect 11107 30454 11175 30510
rect 11231 30454 11299 30510
rect 11355 30454 11423 30510
rect 11479 30454 11547 30510
rect 11603 30454 11671 30510
rect 11727 30454 11795 30510
rect 11851 30454 11919 30510
rect 11975 30454 12043 30510
rect 12099 30454 12167 30510
rect 12223 30454 12291 30510
rect 12347 30454 12415 30510
rect 12471 30454 12481 30510
rect 10669 30386 12481 30454
rect 10669 30330 10679 30386
rect 10735 30330 10803 30386
rect 10859 30330 10927 30386
rect 10983 30330 11051 30386
rect 11107 30330 11175 30386
rect 11231 30330 11299 30386
rect 11355 30330 11423 30386
rect 11479 30330 11547 30386
rect 11603 30330 11671 30386
rect 11727 30330 11795 30386
rect 11851 30330 11919 30386
rect 11975 30330 12043 30386
rect 12099 30330 12167 30386
rect 12223 30330 12291 30386
rect 12347 30330 12415 30386
rect 12471 30330 12481 30386
rect 10669 30262 12481 30330
rect 10669 30206 10679 30262
rect 10735 30206 10803 30262
rect 10859 30206 10927 30262
rect 10983 30206 11051 30262
rect 11107 30206 11175 30262
rect 11231 30206 11299 30262
rect 11355 30206 11423 30262
rect 11479 30206 11547 30262
rect 11603 30206 11671 30262
rect 11727 30206 11795 30262
rect 11851 30206 11919 30262
rect 11975 30206 12043 30262
rect 12099 30206 12167 30262
rect 12223 30206 12291 30262
rect 12347 30206 12415 30262
rect 12471 30206 12481 30262
rect 10669 30138 12481 30206
rect 10669 30082 10679 30138
rect 10735 30082 10803 30138
rect 10859 30082 10927 30138
rect 10983 30082 11051 30138
rect 11107 30082 11175 30138
rect 11231 30082 11299 30138
rect 11355 30082 11423 30138
rect 11479 30082 11547 30138
rect 11603 30082 11671 30138
rect 11727 30082 11795 30138
rect 11851 30082 11919 30138
rect 11975 30082 12043 30138
rect 12099 30082 12167 30138
rect 12223 30082 12291 30138
rect 12347 30082 12415 30138
rect 12471 30082 12481 30138
rect 10669 30014 12481 30082
rect 10669 29958 10679 30014
rect 10735 29958 10803 30014
rect 10859 29958 10927 30014
rect 10983 29958 11051 30014
rect 11107 29958 11175 30014
rect 11231 29958 11299 30014
rect 11355 29958 11423 30014
rect 11479 29958 11547 30014
rect 11603 29958 11671 30014
rect 11727 29958 11795 30014
rect 11851 29958 11919 30014
rect 11975 29958 12043 30014
rect 12099 29958 12167 30014
rect 12223 29958 12291 30014
rect 12347 29958 12415 30014
rect 12471 29958 12481 30014
rect 10669 29890 12481 29958
rect 10669 29834 10679 29890
rect 10735 29834 10803 29890
rect 10859 29834 10927 29890
rect 10983 29834 11051 29890
rect 11107 29834 11175 29890
rect 11231 29834 11299 29890
rect 11355 29834 11423 29890
rect 11479 29834 11547 29890
rect 11603 29834 11671 29890
rect 11727 29834 11795 29890
rect 11851 29834 11919 29890
rect 11975 29834 12043 29890
rect 12099 29834 12167 29890
rect 12223 29834 12291 29890
rect 12347 29834 12415 29890
rect 12471 29834 12481 29890
rect 10669 29766 12481 29834
rect 10669 29710 10679 29766
rect 10735 29710 10803 29766
rect 10859 29710 10927 29766
rect 10983 29710 11051 29766
rect 11107 29710 11175 29766
rect 11231 29710 11299 29766
rect 11355 29710 11423 29766
rect 11479 29710 11547 29766
rect 11603 29710 11671 29766
rect 11727 29710 11795 29766
rect 11851 29710 11919 29766
rect 11975 29710 12043 29766
rect 12099 29710 12167 29766
rect 12223 29710 12291 29766
rect 12347 29710 12415 29766
rect 12471 29710 12481 29766
rect 10669 29642 12481 29710
rect 10669 29586 10679 29642
rect 10735 29586 10803 29642
rect 10859 29586 10927 29642
rect 10983 29586 11051 29642
rect 11107 29586 11175 29642
rect 11231 29586 11299 29642
rect 11355 29586 11423 29642
rect 11479 29586 11547 29642
rect 11603 29586 11671 29642
rect 11727 29586 11795 29642
rect 11851 29586 11919 29642
rect 11975 29586 12043 29642
rect 12099 29586 12167 29642
rect 12223 29586 12291 29642
rect 12347 29586 12415 29642
rect 12471 29586 12481 29642
rect 10669 29518 12481 29586
rect 10669 29462 10679 29518
rect 10735 29462 10803 29518
rect 10859 29462 10927 29518
rect 10983 29462 11051 29518
rect 11107 29462 11175 29518
rect 11231 29462 11299 29518
rect 11355 29462 11423 29518
rect 11479 29462 11547 29518
rect 11603 29462 11671 29518
rect 11727 29462 11795 29518
rect 11851 29462 11919 29518
rect 11975 29462 12043 29518
rect 12099 29462 12167 29518
rect 12223 29462 12291 29518
rect 12347 29462 12415 29518
rect 12471 29462 12481 29518
rect 10669 29394 12481 29462
rect 10669 29338 10679 29394
rect 10735 29338 10803 29394
rect 10859 29338 10927 29394
rect 10983 29338 11051 29394
rect 11107 29338 11175 29394
rect 11231 29338 11299 29394
rect 11355 29338 11423 29394
rect 11479 29338 11547 29394
rect 11603 29338 11671 29394
rect 11727 29338 11795 29394
rect 11851 29338 11919 29394
rect 11975 29338 12043 29394
rect 12099 29338 12167 29394
rect 12223 29338 12291 29394
rect 12347 29338 12415 29394
rect 12471 29338 12481 29394
rect 10669 29270 12481 29338
rect 10669 29214 10679 29270
rect 10735 29214 10803 29270
rect 10859 29214 10927 29270
rect 10983 29214 11051 29270
rect 11107 29214 11175 29270
rect 11231 29214 11299 29270
rect 11355 29214 11423 29270
rect 11479 29214 11547 29270
rect 11603 29214 11671 29270
rect 11727 29214 11795 29270
rect 11851 29214 11919 29270
rect 11975 29214 12043 29270
rect 12099 29214 12167 29270
rect 12223 29214 12291 29270
rect 12347 29214 12415 29270
rect 12471 29214 12481 29270
rect 10669 29146 12481 29214
rect 10669 29090 10679 29146
rect 10735 29090 10803 29146
rect 10859 29090 10927 29146
rect 10983 29090 11051 29146
rect 11107 29090 11175 29146
rect 11231 29090 11299 29146
rect 11355 29090 11423 29146
rect 11479 29090 11547 29146
rect 11603 29090 11671 29146
rect 11727 29090 11795 29146
rect 11851 29090 11919 29146
rect 11975 29090 12043 29146
rect 12099 29090 12167 29146
rect 12223 29090 12291 29146
rect 12347 29090 12415 29146
rect 12471 29090 12481 29146
rect 10669 29022 12481 29090
rect 10669 28966 10679 29022
rect 10735 28966 10803 29022
rect 10859 28966 10927 29022
rect 10983 28966 11051 29022
rect 11107 28966 11175 29022
rect 11231 28966 11299 29022
rect 11355 28966 11423 29022
rect 11479 28966 11547 29022
rect 11603 28966 11671 29022
rect 11727 28966 11795 29022
rect 11851 28966 11919 29022
rect 11975 28966 12043 29022
rect 12099 28966 12167 29022
rect 12223 28966 12291 29022
rect 12347 28966 12415 29022
rect 12471 28966 12481 29022
rect 10669 28898 12481 28966
rect 10669 28842 10679 28898
rect 10735 28842 10803 28898
rect 10859 28842 10927 28898
rect 10983 28842 11051 28898
rect 11107 28842 11175 28898
rect 11231 28842 11299 28898
rect 11355 28842 11423 28898
rect 11479 28842 11547 28898
rect 11603 28842 11671 28898
rect 11727 28842 11795 28898
rect 11851 28842 11919 28898
rect 11975 28842 12043 28898
rect 12099 28842 12167 28898
rect 12223 28842 12291 28898
rect 12347 28842 12415 28898
rect 12471 28842 12481 28898
rect 10669 28832 12481 28842
rect 1489 28742 1499 28798
rect 1555 28742 1565 28798
rect 1489 28674 1565 28742
rect 1489 28618 1499 28674
rect 1555 28618 1565 28674
rect 1489 28550 1565 28618
rect 1489 28494 1499 28550
rect 1555 28494 1565 28550
rect 1489 28426 1565 28494
rect 1489 28370 1499 28426
rect 1555 28370 1565 28426
rect 1489 28302 1565 28370
rect 1489 28246 1499 28302
rect 1555 28246 1565 28302
rect 1489 28178 1565 28246
rect 1489 28122 1499 28178
rect 1555 28122 1565 28178
rect 1489 28054 1565 28122
rect 1489 27998 1499 28054
rect 1555 27998 1565 28054
rect 1489 27930 1565 27998
rect 1489 27874 1499 27930
rect 1555 27874 1565 27930
rect 1489 27806 1565 27874
rect 1489 27750 1499 27806
rect 1555 27750 1565 27806
rect 1489 27682 1565 27750
rect 1489 27626 1499 27682
rect 1555 27626 1565 27682
rect 1489 27558 1565 27626
rect 1489 27502 1499 27558
rect 1555 27502 1565 27558
rect 1489 27434 1565 27502
rect 1489 27378 1499 27434
rect 1555 27378 1565 27434
rect 1489 27310 1565 27378
rect 1489 27254 1499 27310
rect 1555 27254 1565 27310
rect 1613 28808 1689 28818
rect 1613 28752 1623 28808
rect 1679 28752 1689 28808
rect 1613 28684 1689 28752
rect 1613 28628 1623 28684
rect 1679 28628 1689 28684
rect 1613 28560 1689 28628
rect 1613 28504 1623 28560
rect 1679 28504 1689 28560
rect 1613 28436 1689 28504
rect 1613 28380 1623 28436
rect 1679 28380 1689 28436
rect 1613 28312 1689 28380
rect 1613 28256 1623 28312
rect 1679 28256 1689 28312
rect 1613 28188 1689 28256
rect 1613 28132 1623 28188
rect 1679 28132 1689 28188
rect 1613 28064 1689 28132
rect 1613 28008 1623 28064
rect 1679 28008 1689 28064
rect 1613 27940 1689 28008
rect 1613 27884 1623 27940
rect 1679 27884 1689 27940
rect 1613 27816 1689 27884
rect 1613 27760 1623 27816
rect 1679 27760 1689 27816
rect 1613 27692 1689 27760
rect 1613 27636 1623 27692
rect 1679 27636 1689 27692
rect 1613 27568 1689 27636
rect 1613 27512 1623 27568
rect 1679 27512 1689 27568
rect 1613 27444 1689 27512
rect 1613 27388 1623 27444
rect 1679 27388 1689 27444
rect 1613 27320 1689 27388
rect 1613 27264 1623 27320
rect 1679 27264 1689 27320
rect 1613 27254 1689 27264
rect 1737 28653 1813 28663
rect 1737 28597 1747 28653
rect 1803 28597 1813 28653
rect 1737 28529 1813 28597
rect 1737 28473 1747 28529
rect 1803 28473 1813 28529
rect 1737 28405 1813 28473
rect 1737 28349 1747 28405
rect 1803 28349 1813 28405
rect 1737 28281 1813 28349
rect 1737 28225 1747 28281
rect 1803 28225 1813 28281
rect 1737 28157 1813 28225
rect 1737 28101 1747 28157
rect 1803 28101 1813 28157
rect 1737 28033 1813 28101
rect 1737 27977 1747 28033
rect 1803 27977 1813 28033
rect 1737 27909 1813 27977
rect 1737 27853 1747 27909
rect 1803 27853 1813 27909
rect 1737 27785 1813 27853
rect 1737 27729 1747 27785
rect 1803 27729 1813 27785
rect 1737 27661 1813 27729
rect 1737 27605 1747 27661
rect 1803 27605 1813 27661
rect 1737 27537 1813 27605
rect 1737 27481 1747 27537
rect 1803 27481 1813 27537
rect 1737 27413 1813 27481
rect 1737 27357 1747 27413
rect 1803 27357 1813 27413
rect 1737 27289 1813 27357
rect 1489 27244 1565 27254
rect 1737 27233 1747 27289
rect 1803 27233 1813 27289
rect 1861 28539 1937 28549
rect 1861 28483 1871 28539
rect 1927 28483 1937 28539
rect 1861 28415 1937 28483
rect 1861 28359 1871 28415
rect 1927 28359 1937 28415
rect 1861 28291 1937 28359
rect 1861 28235 1871 28291
rect 1927 28235 1937 28291
rect 1861 28167 1937 28235
rect 1861 28111 1871 28167
rect 1927 28111 1937 28167
rect 1861 28043 1937 28111
rect 1861 27987 1871 28043
rect 1927 27987 1937 28043
rect 1861 27919 1937 27987
rect 1861 27863 1871 27919
rect 1927 27863 1937 27919
rect 1861 27795 1937 27863
rect 1861 27739 1871 27795
rect 1927 27739 1937 27795
rect 1861 27671 1937 27739
rect 1861 27615 1871 27671
rect 1927 27615 1937 27671
rect 1861 27547 1937 27615
rect 1861 27491 1871 27547
rect 1927 27491 1937 27547
rect 1861 27423 1937 27491
rect 1861 27367 1871 27423
rect 1927 27367 1937 27423
rect 1861 27299 1937 27367
rect 1861 27243 1871 27299
rect 1927 27243 1937 27299
rect 1861 27233 1937 27243
rect 1985 28537 2061 28547
rect 1985 28481 1995 28537
rect 2051 28481 2061 28537
rect 1985 28413 2061 28481
rect 1985 28357 1995 28413
rect 2051 28357 2061 28413
rect 1985 28289 2061 28357
rect 1985 28233 1995 28289
rect 2051 28233 2061 28289
rect 1985 28165 2061 28233
rect 1985 28109 1995 28165
rect 2051 28109 2061 28165
rect 1985 28041 2061 28109
rect 1985 27985 1995 28041
rect 2051 27985 2061 28041
rect 1985 27917 2061 27985
rect 1985 27861 1995 27917
rect 2051 27861 2061 27917
rect 1985 27793 2061 27861
rect 1985 27737 1995 27793
rect 2051 27737 2061 27793
rect 1985 27669 2061 27737
rect 1985 27613 1995 27669
rect 2051 27613 2061 27669
rect 1985 27545 2061 27613
rect 1985 27489 1995 27545
rect 2051 27489 2061 27545
rect 1985 27421 2061 27489
rect 1985 27365 1995 27421
rect 2051 27365 2061 27421
rect 1985 27297 2061 27365
rect 1985 27241 1995 27297
rect 2051 27241 2061 27297
rect 1737 27223 1813 27233
rect 1985 27231 2061 27241
rect 4425 28544 6237 28554
rect 4425 28488 4435 28544
rect 4491 28488 4559 28544
rect 4615 28488 4683 28544
rect 4739 28488 4807 28544
rect 4863 28488 4931 28544
rect 4987 28488 5055 28544
rect 5111 28488 5179 28544
rect 5235 28488 5303 28544
rect 5359 28488 5427 28544
rect 5483 28488 5551 28544
rect 5607 28488 5675 28544
rect 5731 28488 5799 28544
rect 5855 28488 5923 28544
rect 5979 28488 6047 28544
rect 6103 28488 6171 28544
rect 6227 28488 6237 28544
rect 4425 28420 6237 28488
rect 4425 28364 4435 28420
rect 4491 28364 4559 28420
rect 4615 28364 4683 28420
rect 4739 28364 4807 28420
rect 4863 28364 4931 28420
rect 4987 28364 5055 28420
rect 5111 28364 5179 28420
rect 5235 28364 5303 28420
rect 5359 28364 5427 28420
rect 5483 28364 5551 28420
rect 5607 28364 5675 28420
rect 5731 28364 5799 28420
rect 5855 28364 5923 28420
rect 5979 28364 6047 28420
rect 6103 28364 6171 28420
rect 6227 28364 6237 28420
rect 4425 28296 6237 28364
rect 4425 28240 4435 28296
rect 4491 28240 4559 28296
rect 4615 28240 4683 28296
rect 4739 28240 4807 28296
rect 4863 28240 4931 28296
rect 4987 28240 5055 28296
rect 5111 28240 5179 28296
rect 5235 28240 5303 28296
rect 5359 28240 5427 28296
rect 5483 28240 5551 28296
rect 5607 28240 5675 28296
rect 5731 28240 5799 28296
rect 5855 28240 5923 28296
rect 5979 28240 6047 28296
rect 6103 28240 6171 28296
rect 6227 28240 6237 28296
rect 4425 28172 6237 28240
rect 4425 28116 4435 28172
rect 4491 28116 4559 28172
rect 4615 28116 4683 28172
rect 4739 28116 4807 28172
rect 4863 28116 4931 28172
rect 4987 28116 5055 28172
rect 5111 28116 5179 28172
rect 5235 28116 5303 28172
rect 5359 28116 5427 28172
rect 5483 28116 5551 28172
rect 5607 28116 5675 28172
rect 5731 28116 5799 28172
rect 5855 28116 5923 28172
rect 5979 28116 6047 28172
rect 6103 28116 6171 28172
rect 6227 28116 6237 28172
rect 4425 28048 6237 28116
rect 4425 27992 4435 28048
rect 4491 27992 4559 28048
rect 4615 27992 4683 28048
rect 4739 27992 4807 28048
rect 4863 27992 4931 28048
rect 4987 27992 5055 28048
rect 5111 27992 5179 28048
rect 5235 27992 5303 28048
rect 5359 27992 5427 28048
rect 5483 27992 5551 28048
rect 5607 27992 5675 28048
rect 5731 27992 5799 28048
rect 5855 27992 5923 28048
rect 5979 27992 6047 28048
rect 6103 27992 6171 28048
rect 6227 27992 6237 28048
rect 4425 27924 6237 27992
rect 4425 27868 4435 27924
rect 4491 27868 4559 27924
rect 4615 27868 4683 27924
rect 4739 27868 4807 27924
rect 4863 27868 4931 27924
rect 4987 27868 5055 27924
rect 5111 27868 5179 27924
rect 5235 27868 5303 27924
rect 5359 27868 5427 27924
rect 5483 27868 5551 27924
rect 5607 27868 5675 27924
rect 5731 27868 5799 27924
rect 5855 27868 5923 27924
rect 5979 27868 6047 27924
rect 6103 27868 6171 27924
rect 6227 27868 6237 27924
rect 4425 27800 6237 27868
rect 4425 27744 4435 27800
rect 4491 27744 4559 27800
rect 4615 27744 4683 27800
rect 4739 27744 4807 27800
rect 4863 27744 4931 27800
rect 4987 27744 5055 27800
rect 5111 27744 5179 27800
rect 5235 27744 5303 27800
rect 5359 27744 5427 27800
rect 5483 27744 5551 27800
rect 5607 27744 5675 27800
rect 5731 27744 5799 27800
rect 5855 27744 5923 27800
rect 5979 27744 6047 27800
rect 6103 27744 6171 27800
rect 6227 27744 6237 27800
rect 4425 27676 6237 27744
rect 4425 27620 4435 27676
rect 4491 27620 4559 27676
rect 4615 27620 4683 27676
rect 4739 27620 4807 27676
rect 4863 27620 4931 27676
rect 4987 27620 5055 27676
rect 5111 27620 5179 27676
rect 5235 27620 5303 27676
rect 5359 27620 5427 27676
rect 5483 27620 5551 27676
rect 5607 27620 5675 27676
rect 5731 27620 5799 27676
rect 5855 27620 5923 27676
rect 5979 27620 6047 27676
rect 6103 27620 6171 27676
rect 6227 27620 6237 27676
rect 4425 27552 6237 27620
rect 4425 27496 4435 27552
rect 4491 27496 4559 27552
rect 4615 27496 4683 27552
rect 4739 27496 4807 27552
rect 4863 27496 4931 27552
rect 4987 27496 5055 27552
rect 5111 27496 5179 27552
rect 5235 27496 5303 27552
rect 5359 27496 5427 27552
rect 5483 27496 5551 27552
rect 5607 27496 5675 27552
rect 5731 27496 5799 27552
rect 5855 27496 5923 27552
rect 5979 27496 6047 27552
rect 6103 27496 6171 27552
rect 6227 27496 6237 27552
rect 4425 27428 6237 27496
rect 4425 27372 4435 27428
rect 4491 27372 4559 27428
rect 4615 27372 4683 27428
rect 4739 27372 4807 27428
rect 4863 27372 4931 27428
rect 4987 27372 5055 27428
rect 5111 27372 5179 27428
rect 5235 27372 5303 27428
rect 5359 27372 5427 27428
rect 5483 27372 5551 27428
rect 5607 27372 5675 27428
rect 5731 27372 5799 27428
rect 5855 27372 5923 27428
rect 5979 27372 6047 27428
rect 6103 27372 6171 27428
rect 6227 27372 6237 27428
rect 4425 27304 6237 27372
rect 4425 27248 4435 27304
rect 4491 27248 4559 27304
rect 4615 27248 4683 27304
rect 4739 27248 4807 27304
rect 4863 27248 4931 27304
rect 4987 27248 5055 27304
rect 5111 27248 5179 27304
rect 5235 27248 5303 27304
rect 5359 27248 5427 27304
rect 5483 27248 5551 27304
rect 5607 27248 5675 27304
rect 5731 27248 5799 27304
rect 5855 27248 5923 27304
rect 5979 27248 6047 27304
rect 6103 27248 6171 27304
rect 6227 27248 6237 27304
rect 4425 27238 6237 27248
rect 7552 28544 8620 28554
rect 7552 28488 7562 28544
rect 7618 28488 7686 28544
rect 7742 28488 7810 28544
rect 7866 28488 7934 28544
rect 7990 28488 8058 28544
rect 8114 28488 8182 28544
rect 8238 28488 8306 28544
rect 8362 28488 8430 28544
rect 8486 28488 8554 28544
rect 8610 28488 8620 28544
rect 7552 28420 8620 28488
rect 7552 28364 7562 28420
rect 7618 28364 7686 28420
rect 7742 28364 7810 28420
rect 7866 28364 7934 28420
rect 7990 28364 8058 28420
rect 8114 28364 8182 28420
rect 8238 28364 8306 28420
rect 8362 28364 8430 28420
rect 8486 28364 8554 28420
rect 8610 28364 8620 28420
rect 7552 28296 8620 28364
rect 7552 28240 7562 28296
rect 7618 28240 7686 28296
rect 7742 28240 7810 28296
rect 7866 28240 7934 28296
rect 7990 28240 8058 28296
rect 8114 28240 8182 28296
rect 8238 28240 8306 28296
rect 8362 28240 8430 28296
rect 8486 28240 8554 28296
rect 8610 28240 8620 28296
rect 7552 28172 8620 28240
rect 7552 28116 7562 28172
rect 7618 28116 7686 28172
rect 7742 28116 7810 28172
rect 7866 28116 7934 28172
rect 7990 28116 8058 28172
rect 8114 28116 8182 28172
rect 8238 28116 8306 28172
rect 8362 28116 8430 28172
rect 8486 28116 8554 28172
rect 8610 28116 8620 28172
rect 7552 28048 8620 28116
rect 7552 27992 7562 28048
rect 7618 27992 7686 28048
rect 7742 27992 7810 28048
rect 7866 27992 7934 28048
rect 7990 27992 8058 28048
rect 8114 27992 8182 28048
rect 8238 27992 8306 28048
rect 8362 27992 8430 28048
rect 8486 27992 8554 28048
rect 8610 27992 8620 28048
rect 7552 27924 8620 27992
rect 7552 27868 7562 27924
rect 7618 27868 7686 27924
rect 7742 27868 7810 27924
rect 7866 27868 7934 27924
rect 7990 27868 8058 27924
rect 8114 27868 8182 27924
rect 8238 27868 8306 27924
rect 8362 27868 8430 27924
rect 8486 27868 8554 27924
rect 8610 27868 8620 27924
rect 7552 27800 8620 27868
rect 7552 27744 7562 27800
rect 7618 27744 7686 27800
rect 7742 27744 7810 27800
rect 7866 27744 7934 27800
rect 7990 27744 8058 27800
rect 8114 27744 8182 27800
rect 8238 27744 8306 27800
rect 8362 27744 8430 27800
rect 8486 27744 8554 27800
rect 8610 27744 8620 27800
rect 7552 27676 8620 27744
rect 7552 27620 7562 27676
rect 7618 27620 7686 27676
rect 7742 27620 7810 27676
rect 7866 27620 7934 27676
rect 7990 27620 8058 27676
rect 8114 27620 8182 27676
rect 8238 27620 8306 27676
rect 8362 27620 8430 27676
rect 8486 27620 8554 27676
rect 8610 27620 8620 27676
rect 7552 27552 8620 27620
rect 7552 27496 7562 27552
rect 7618 27496 7686 27552
rect 7742 27496 7810 27552
rect 7866 27496 7934 27552
rect 7990 27496 8058 27552
rect 8114 27496 8182 27552
rect 8238 27496 8306 27552
rect 8362 27496 8430 27552
rect 8486 27496 8554 27552
rect 8610 27496 8620 27552
rect 7552 27428 8620 27496
rect 7552 27372 7562 27428
rect 7618 27372 7686 27428
rect 7742 27372 7810 27428
rect 7866 27372 7934 27428
rect 7990 27372 8058 27428
rect 8114 27372 8182 27428
rect 8238 27372 8306 27428
rect 8362 27372 8430 27428
rect 8486 27372 8554 27428
rect 8610 27372 8620 27428
rect 7552 27304 8620 27372
rect 7552 27248 7562 27304
rect 7618 27248 7686 27304
rect 7742 27248 7810 27304
rect 7866 27248 7934 27304
rect 7990 27248 8058 27304
rect 8114 27248 8182 27304
rect 8238 27248 8306 27304
rect 8362 27248 8430 27304
rect 8486 27248 8554 27304
rect 8610 27248 8620 27304
rect 7552 27238 8620 27248
rect 10669 28544 12481 28554
rect 10669 28488 10679 28544
rect 10735 28488 10803 28544
rect 10859 28488 10927 28544
rect 10983 28488 11051 28544
rect 11107 28488 11175 28544
rect 11231 28488 11299 28544
rect 11355 28488 11423 28544
rect 11479 28488 11547 28544
rect 11603 28488 11671 28544
rect 11727 28488 11795 28544
rect 11851 28488 11919 28544
rect 11975 28488 12043 28544
rect 12099 28488 12167 28544
rect 12223 28488 12291 28544
rect 12347 28488 12415 28544
rect 12471 28488 12481 28544
rect 10669 28420 12481 28488
rect 10669 28364 10679 28420
rect 10735 28364 10803 28420
rect 10859 28364 10927 28420
rect 10983 28364 11051 28420
rect 11107 28364 11175 28420
rect 11231 28364 11299 28420
rect 11355 28364 11423 28420
rect 11479 28364 11547 28420
rect 11603 28364 11671 28420
rect 11727 28364 11795 28420
rect 11851 28364 11919 28420
rect 11975 28364 12043 28420
rect 12099 28364 12167 28420
rect 12223 28364 12291 28420
rect 12347 28364 12415 28420
rect 12471 28364 12481 28420
rect 10669 28296 12481 28364
rect 10669 28240 10679 28296
rect 10735 28240 10803 28296
rect 10859 28240 10927 28296
rect 10983 28240 11051 28296
rect 11107 28240 11175 28296
rect 11231 28240 11299 28296
rect 11355 28240 11423 28296
rect 11479 28240 11547 28296
rect 11603 28240 11671 28296
rect 11727 28240 11795 28296
rect 11851 28240 11919 28296
rect 11975 28240 12043 28296
rect 12099 28240 12167 28296
rect 12223 28240 12291 28296
rect 12347 28240 12415 28296
rect 12471 28240 12481 28296
rect 10669 28172 12481 28240
rect 10669 28116 10679 28172
rect 10735 28116 10803 28172
rect 10859 28116 10927 28172
rect 10983 28116 11051 28172
rect 11107 28116 11175 28172
rect 11231 28116 11299 28172
rect 11355 28116 11423 28172
rect 11479 28116 11547 28172
rect 11603 28116 11671 28172
rect 11727 28116 11795 28172
rect 11851 28116 11919 28172
rect 11975 28116 12043 28172
rect 12099 28116 12167 28172
rect 12223 28116 12291 28172
rect 12347 28116 12415 28172
rect 12471 28116 12481 28172
rect 10669 28048 12481 28116
rect 10669 27992 10679 28048
rect 10735 27992 10803 28048
rect 10859 27992 10927 28048
rect 10983 27992 11051 28048
rect 11107 27992 11175 28048
rect 11231 27992 11299 28048
rect 11355 27992 11423 28048
rect 11479 27992 11547 28048
rect 11603 27992 11671 28048
rect 11727 27992 11795 28048
rect 11851 27992 11919 28048
rect 11975 27992 12043 28048
rect 12099 27992 12167 28048
rect 12223 27992 12291 28048
rect 12347 27992 12415 28048
rect 12471 27992 12481 28048
rect 10669 27924 12481 27992
rect 10669 27868 10679 27924
rect 10735 27868 10803 27924
rect 10859 27868 10927 27924
rect 10983 27868 11051 27924
rect 11107 27868 11175 27924
rect 11231 27868 11299 27924
rect 11355 27868 11423 27924
rect 11479 27868 11547 27924
rect 11603 27868 11671 27924
rect 11727 27868 11795 27924
rect 11851 27868 11919 27924
rect 11975 27868 12043 27924
rect 12099 27868 12167 27924
rect 12223 27868 12291 27924
rect 12347 27868 12415 27924
rect 12471 27868 12481 27924
rect 10669 27800 12481 27868
rect 10669 27744 10679 27800
rect 10735 27744 10803 27800
rect 10859 27744 10927 27800
rect 10983 27744 11051 27800
rect 11107 27744 11175 27800
rect 11231 27744 11299 27800
rect 11355 27744 11423 27800
rect 11479 27744 11547 27800
rect 11603 27744 11671 27800
rect 11727 27744 11795 27800
rect 11851 27744 11919 27800
rect 11975 27744 12043 27800
rect 12099 27744 12167 27800
rect 12223 27744 12291 27800
rect 12347 27744 12415 27800
rect 12471 27744 12481 27800
rect 10669 27676 12481 27744
rect 10669 27620 10679 27676
rect 10735 27620 10803 27676
rect 10859 27620 10927 27676
rect 10983 27620 11051 27676
rect 11107 27620 11175 27676
rect 11231 27620 11299 27676
rect 11355 27620 11423 27676
rect 11479 27620 11547 27676
rect 11603 27620 11671 27676
rect 11727 27620 11795 27676
rect 11851 27620 11919 27676
rect 11975 27620 12043 27676
rect 12099 27620 12167 27676
rect 12223 27620 12291 27676
rect 12347 27620 12415 27676
rect 12471 27620 12481 27676
rect 10669 27552 12481 27620
rect 10669 27496 10679 27552
rect 10735 27496 10803 27552
rect 10859 27496 10927 27552
rect 10983 27496 11051 27552
rect 11107 27496 11175 27552
rect 11231 27496 11299 27552
rect 11355 27496 11423 27552
rect 11479 27496 11547 27552
rect 11603 27496 11671 27552
rect 11727 27496 11795 27552
rect 11851 27496 11919 27552
rect 11975 27496 12043 27552
rect 12099 27496 12167 27552
rect 12223 27496 12291 27552
rect 12347 27496 12415 27552
rect 12471 27496 12481 27552
rect 10669 27428 12481 27496
rect 10669 27372 10679 27428
rect 10735 27372 10803 27428
rect 10859 27372 10927 27428
rect 10983 27372 11051 27428
rect 11107 27372 11175 27428
rect 11231 27372 11299 27428
rect 11355 27372 11423 27428
rect 11479 27372 11547 27428
rect 11603 27372 11671 27428
rect 11727 27372 11795 27428
rect 11851 27372 11919 27428
rect 11975 27372 12043 27428
rect 12099 27372 12167 27428
rect 12223 27372 12291 27428
rect 12347 27372 12415 27428
rect 12471 27372 12481 27428
rect 10669 27304 12481 27372
rect 10669 27248 10679 27304
rect 10735 27248 10803 27304
rect 10859 27248 10927 27304
rect 10983 27248 11051 27304
rect 11107 27248 11175 27304
rect 11231 27248 11299 27304
rect 11355 27248 11423 27304
rect 11479 27248 11547 27304
rect 11603 27248 11671 27304
rect 11727 27248 11795 27304
rect 11851 27248 11919 27304
rect 11975 27248 12043 27304
rect 12099 27248 12167 27304
rect 12223 27248 12291 27304
rect 12347 27248 12415 27304
rect 12471 27248 12481 27304
rect 10669 27238 12481 27248
rect 2497 26944 4309 26954
rect 2497 26888 2507 26944
rect 2563 26888 2631 26944
rect 2687 26888 2755 26944
rect 2811 26888 2879 26944
rect 2935 26888 3003 26944
rect 3059 26888 3127 26944
rect 3183 26888 3251 26944
rect 3307 26888 3375 26944
rect 3431 26888 3499 26944
rect 3555 26888 3623 26944
rect 3679 26888 3747 26944
rect 3803 26888 3871 26944
rect 3927 26888 3995 26944
rect 4051 26888 4119 26944
rect 4175 26888 4243 26944
rect 4299 26888 4309 26944
rect 2497 26820 4309 26888
rect 2497 26764 2507 26820
rect 2563 26764 2631 26820
rect 2687 26764 2755 26820
rect 2811 26764 2879 26820
rect 2935 26764 3003 26820
rect 3059 26764 3127 26820
rect 3183 26764 3251 26820
rect 3307 26764 3375 26820
rect 3431 26764 3499 26820
rect 3555 26764 3623 26820
rect 3679 26764 3747 26820
rect 3803 26764 3871 26820
rect 3927 26764 3995 26820
rect 4051 26764 4119 26820
rect 4175 26764 4243 26820
rect 4299 26764 4309 26820
rect 2497 26696 4309 26764
rect 2497 26640 2507 26696
rect 2563 26640 2631 26696
rect 2687 26640 2755 26696
rect 2811 26640 2879 26696
rect 2935 26640 3003 26696
rect 3059 26640 3127 26696
rect 3183 26640 3251 26696
rect 3307 26640 3375 26696
rect 3431 26640 3499 26696
rect 3555 26640 3623 26696
rect 3679 26640 3747 26696
rect 3803 26640 3871 26696
rect 3927 26640 3995 26696
rect 4051 26640 4119 26696
rect 4175 26640 4243 26696
rect 4299 26640 4309 26696
rect 2497 26572 4309 26640
rect 2497 26516 2507 26572
rect 2563 26516 2631 26572
rect 2687 26516 2755 26572
rect 2811 26516 2879 26572
rect 2935 26516 3003 26572
rect 3059 26516 3127 26572
rect 3183 26516 3251 26572
rect 3307 26516 3375 26572
rect 3431 26516 3499 26572
rect 3555 26516 3623 26572
rect 3679 26516 3747 26572
rect 3803 26516 3871 26572
rect 3927 26516 3995 26572
rect 4051 26516 4119 26572
rect 4175 26516 4243 26572
rect 4299 26516 4309 26572
rect 2497 26448 4309 26516
rect 2497 26392 2507 26448
rect 2563 26392 2631 26448
rect 2687 26392 2755 26448
rect 2811 26392 2879 26448
rect 2935 26392 3003 26448
rect 3059 26392 3127 26448
rect 3183 26392 3251 26448
rect 3307 26392 3375 26448
rect 3431 26392 3499 26448
rect 3555 26392 3623 26448
rect 3679 26392 3747 26448
rect 3803 26392 3871 26448
rect 3927 26392 3995 26448
rect 4051 26392 4119 26448
rect 4175 26392 4243 26448
rect 4299 26392 4309 26448
rect 2497 26324 4309 26392
rect 2497 26268 2507 26324
rect 2563 26268 2631 26324
rect 2687 26268 2755 26324
rect 2811 26268 2879 26324
rect 2935 26268 3003 26324
rect 3059 26268 3127 26324
rect 3183 26268 3251 26324
rect 3307 26268 3375 26324
rect 3431 26268 3499 26324
rect 3555 26268 3623 26324
rect 3679 26268 3747 26324
rect 3803 26268 3871 26324
rect 3927 26268 3995 26324
rect 4051 26268 4119 26324
rect 4175 26268 4243 26324
rect 4299 26268 4309 26324
rect 2497 26200 4309 26268
rect 2497 26144 2507 26200
rect 2563 26144 2631 26200
rect 2687 26144 2755 26200
rect 2811 26144 2879 26200
rect 2935 26144 3003 26200
rect 3059 26144 3127 26200
rect 3183 26144 3251 26200
rect 3307 26144 3375 26200
rect 3431 26144 3499 26200
rect 3555 26144 3623 26200
rect 3679 26144 3747 26200
rect 3803 26144 3871 26200
rect 3927 26144 3995 26200
rect 4051 26144 4119 26200
rect 4175 26144 4243 26200
rect 4299 26144 4309 26200
rect 2497 26076 4309 26144
rect 2497 26020 2507 26076
rect 2563 26020 2631 26076
rect 2687 26020 2755 26076
rect 2811 26020 2879 26076
rect 2935 26020 3003 26076
rect 3059 26020 3127 26076
rect 3183 26020 3251 26076
rect 3307 26020 3375 26076
rect 3431 26020 3499 26076
rect 3555 26020 3623 26076
rect 3679 26020 3747 26076
rect 3803 26020 3871 26076
rect 3927 26020 3995 26076
rect 4051 26020 4119 26076
rect 4175 26020 4243 26076
rect 4299 26020 4309 26076
rect 2497 25952 4309 26020
rect 2497 25896 2507 25952
rect 2563 25896 2631 25952
rect 2687 25896 2755 25952
rect 2811 25896 2879 25952
rect 2935 25896 3003 25952
rect 3059 25896 3127 25952
rect 3183 25896 3251 25952
rect 3307 25896 3375 25952
rect 3431 25896 3499 25952
rect 3555 25896 3623 25952
rect 3679 25896 3747 25952
rect 3803 25896 3871 25952
rect 3927 25896 3995 25952
rect 4051 25896 4119 25952
rect 4175 25896 4243 25952
rect 4299 25896 4309 25952
rect 2497 25828 4309 25896
rect 2497 25772 2507 25828
rect 2563 25772 2631 25828
rect 2687 25772 2755 25828
rect 2811 25772 2879 25828
rect 2935 25772 3003 25828
rect 3059 25772 3127 25828
rect 3183 25772 3251 25828
rect 3307 25772 3375 25828
rect 3431 25772 3499 25828
rect 3555 25772 3623 25828
rect 3679 25772 3747 25828
rect 3803 25772 3871 25828
rect 3927 25772 3995 25828
rect 4051 25772 4119 25828
rect 4175 25772 4243 25828
rect 4299 25772 4309 25828
rect 2497 25704 4309 25772
rect 2497 25648 2507 25704
rect 2563 25648 2631 25704
rect 2687 25648 2755 25704
rect 2811 25648 2879 25704
rect 2935 25648 3003 25704
rect 3059 25648 3127 25704
rect 3183 25648 3251 25704
rect 3307 25648 3375 25704
rect 3431 25648 3499 25704
rect 3555 25648 3623 25704
rect 3679 25648 3747 25704
rect 3803 25648 3871 25704
rect 3927 25648 3995 25704
rect 4051 25648 4119 25704
rect 4175 25648 4243 25704
rect 4299 25648 4309 25704
rect 2497 25638 4309 25648
rect 6358 26944 7426 26954
rect 6358 26888 6368 26944
rect 6424 26888 6492 26944
rect 6548 26888 6616 26944
rect 6672 26888 6740 26944
rect 6796 26888 6864 26944
rect 6920 26888 6988 26944
rect 7044 26888 7112 26944
rect 7168 26888 7236 26944
rect 7292 26888 7360 26944
rect 7416 26888 7426 26944
rect 6358 26820 7426 26888
rect 6358 26764 6368 26820
rect 6424 26764 6492 26820
rect 6548 26764 6616 26820
rect 6672 26764 6740 26820
rect 6796 26764 6864 26820
rect 6920 26764 6988 26820
rect 7044 26764 7112 26820
rect 7168 26764 7236 26820
rect 7292 26764 7360 26820
rect 7416 26764 7426 26820
rect 6358 26696 7426 26764
rect 6358 26640 6368 26696
rect 6424 26640 6492 26696
rect 6548 26640 6616 26696
rect 6672 26640 6740 26696
rect 6796 26640 6864 26696
rect 6920 26640 6988 26696
rect 7044 26640 7112 26696
rect 7168 26640 7236 26696
rect 7292 26640 7360 26696
rect 7416 26640 7426 26696
rect 6358 26572 7426 26640
rect 6358 26516 6368 26572
rect 6424 26516 6492 26572
rect 6548 26516 6616 26572
rect 6672 26516 6740 26572
rect 6796 26516 6864 26572
rect 6920 26516 6988 26572
rect 7044 26516 7112 26572
rect 7168 26516 7236 26572
rect 7292 26516 7360 26572
rect 7416 26516 7426 26572
rect 6358 26448 7426 26516
rect 6358 26392 6368 26448
rect 6424 26392 6492 26448
rect 6548 26392 6616 26448
rect 6672 26392 6740 26448
rect 6796 26392 6864 26448
rect 6920 26392 6988 26448
rect 7044 26392 7112 26448
rect 7168 26392 7236 26448
rect 7292 26392 7360 26448
rect 7416 26392 7426 26448
rect 6358 26324 7426 26392
rect 6358 26268 6368 26324
rect 6424 26268 6492 26324
rect 6548 26268 6616 26324
rect 6672 26268 6740 26324
rect 6796 26268 6864 26324
rect 6920 26268 6988 26324
rect 7044 26268 7112 26324
rect 7168 26268 7236 26324
rect 7292 26268 7360 26324
rect 7416 26268 7426 26324
rect 6358 26200 7426 26268
rect 6358 26144 6368 26200
rect 6424 26144 6492 26200
rect 6548 26144 6616 26200
rect 6672 26144 6740 26200
rect 6796 26144 6864 26200
rect 6920 26144 6988 26200
rect 7044 26144 7112 26200
rect 7168 26144 7236 26200
rect 7292 26144 7360 26200
rect 7416 26144 7426 26200
rect 6358 26076 7426 26144
rect 6358 26020 6368 26076
rect 6424 26020 6492 26076
rect 6548 26020 6616 26076
rect 6672 26020 6740 26076
rect 6796 26020 6864 26076
rect 6920 26020 6988 26076
rect 7044 26020 7112 26076
rect 7168 26020 7236 26076
rect 7292 26020 7360 26076
rect 7416 26020 7426 26076
rect 6358 25952 7426 26020
rect 6358 25896 6368 25952
rect 6424 25896 6492 25952
rect 6548 25896 6616 25952
rect 6672 25896 6740 25952
rect 6796 25896 6864 25952
rect 6920 25896 6988 25952
rect 7044 25896 7112 25952
rect 7168 25896 7236 25952
rect 7292 25896 7360 25952
rect 7416 25896 7426 25952
rect 6358 25828 7426 25896
rect 6358 25772 6368 25828
rect 6424 25772 6492 25828
rect 6548 25772 6616 25828
rect 6672 25772 6740 25828
rect 6796 25772 6864 25828
rect 6920 25772 6988 25828
rect 7044 25772 7112 25828
rect 7168 25772 7236 25828
rect 7292 25772 7360 25828
rect 7416 25772 7426 25828
rect 6358 25704 7426 25772
rect 6358 25648 6368 25704
rect 6424 25648 6492 25704
rect 6548 25648 6616 25704
rect 6672 25648 6740 25704
rect 6796 25648 6864 25704
rect 6920 25648 6988 25704
rect 7044 25648 7112 25704
rect 7168 25648 7236 25704
rect 7292 25648 7360 25704
rect 7416 25648 7426 25704
rect 6358 25638 7426 25648
rect 8741 26944 10553 26954
rect 8741 26888 8751 26944
rect 8807 26888 8875 26944
rect 8931 26888 8999 26944
rect 9055 26888 9123 26944
rect 9179 26888 9247 26944
rect 9303 26888 9371 26944
rect 9427 26888 9495 26944
rect 9551 26888 9619 26944
rect 9675 26888 9743 26944
rect 9799 26888 9867 26944
rect 9923 26888 9991 26944
rect 10047 26888 10115 26944
rect 10171 26888 10239 26944
rect 10295 26888 10363 26944
rect 10419 26888 10487 26944
rect 10543 26888 10553 26944
rect 8741 26820 10553 26888
rect 8741 26764 8751 26820
rect 8807 26764 8875 26820
rect 8931 26764 8999 26820
rect 9055 26764 9123 26820
rect 9179 26764 9247 26820
rect 9303 26764 9371 26820
rect 9427 26764 9495 26820
rect 9551 26764 9619 26820
rect 9675 26764 9743 26820
rect 9799 26764 9867 26820
rect 9923 26764 9991 26820
rect 10047 26764 10115 26820
rect 10171 26764 10239 26820
rect 10295 26764 10363 26820
rect 10419 26764 10487 26820
rect 10543 26764 10553 26820
rect 8741 26696 10553 26764
rect 8741 26640 8751 26696
rect 8807 26640 8875 26696
rect 8931 26640 8999 26696
rect 9055 26640 9123 26696
rect 9179 26640 9247 26696
rect 9303 26640 9371 26696
rect 9427 26640 9495 26696
rect 9551 26640 9619 26696
rect 9675 26640 9743 26696
rect 9799 26640 9867 26696
rect 9923 26640 9991 26696
rect 10047 26640 10115 26696
rect 10171 26640 10239 26696
rect 10295 26640 10363 26696
rect 10419 26640 10487 26696
rect 10543 26640 10553 26696
rect 8741 26572 10553 26640
rect 8741 26516 8751 26572
rect 8807 26516 8875 26572
rect 8931 26516 8999 26572
rect 9055 26516 9123 26572
rect 9179 26516 9247 26572
rect 9303 26516 9371 26572
rect 9427 26516 9495 26572
rect 9551 26516 9619 26572
rect 9675 26516 9743 26572
rect 9799 26516 9867 26572
rect 9923 26516 9991 26572
rect 10047 26516 10115 26572
rect 10171 26516 10239 26572
rect 10295 26516 10363 26572
rect 10419 26516 10487 26572
rect 10543 26516 10553 26572
rect 8741 26448 10553 26516
rect 8741 26392 8751 26448
rect 8807 26392 8875 26448
rect 8931 26392 8999 26448
rect 9055 26392 9123 26448
rect 9179 26392 9247 26448
rect 9303 26392 9371 26448
rect 9427 26392 9495 26448
rect 9551 26392 9619 26448
rect 9675 26392 9743 26448
rect 9799 26392 9867 26448
rect 9923 26392 9991 26448
rect 10047 26392 10115 26448
rect 10171 26392 10239 26448
rect 10295 26392 10363 26448
rect 10419 26392 10487 26448
rect 10543 26392 10553 26448
rect 8741 26324 10553 26392
rect 8741 26268 8751 26324
rect 8807 26268 8875 26324
rect 8931 26268 8999 26324
rect 9055 26268 9123 26324
rect 9179 26268 9247 26324
rect 9303 26268 9371 26324
rect 9427 26268 9495 26324
rect 9551 26268 9619 26324
rect 9675 26268 9743 26324
rect 9799 26268 9867 26324
rect 9923 26268 9991 26324
rect 10047 26268 10115 26324
rect 10171 26268 10239 26324
rect 10295 26268 10363 26324
rect 10419 26268 10487 26324
rect 10543 26268 10553 26324
rect 8741 26200 10553 26268
rect 8741 26144 8751 26200
rect 8807 26144 8875 26200
rect 8931 26144 8999 26200
rect 9055 26144 9123 26200
rect 9179 26144 9247 26200
rect 9303 26144 9371 26200
rect 9427 26144 9495 26200
rect 9551 26144 9619 26200
rect 9675 26144 9743 26200
rect 9799 26144 9867 26200
rect 9923 26144 9991 26200
rect 10047 26144 10115 26200
rect 10171 26144 10239 26200
rect 10295 26144 10363 26200
rect 10419 26144 10487 26200
rect 10543 26144 10553 26200
rect 8741 26076 10553 26144
rect 8741 26020 8751 26076
rect 8807 26020 8875 26076
rect 8931 26020 8999 26076
rect 9055 26020 9123 26076
rect 9179 26020 9247 26076
rect 9303 26020 9371 26076
rect 9427 26020 9495 26076
rect 9551 26020 9619 26076
rect 9675 26020 9743 26076
rect 9799 26020 9867 26076
rect 9923 26020 9991 26076
rect 10047 26020 10115 26076
rect 10171 26020 10239 26076
rect 10295 26020 10363 26076
rect 10419 26020 10487 26076
rect 10543 26020 10553 26076
rect 8741 25952 10553 26020
rect 8741 25896 8751 25952
rect 8807 25896 8875 25952
rect 8931 25896 8999 25952
rect 9055 25896 9123 25952
rect 9179 25896 9247 25952
rect 9303 25896 9371 25952
rect 9427 25896 9495 25952
rect 9551 25896 9619 25952
rect 9675 25896 9743 25952
rect 9799 25896 9867 25952
rect 9923 25896 9991 25952
rect 10047 25896 10115 25952
rect 10171 25896 10239 25952
rect 10295 25896 10363 25952
rect 10419 25896 10487 25952
rect 10543 25896 10553 25952
rect 8741 25828 10553 25896
rect 8741 25772 8751 25828
rect 8807 25772 8875 25828
rect 8931 25772 8999 25828
rect 9055 25772 9123 25828
rect 9179 25772 9247 25828
rect 9303 25772 9371 25828
rect 9427 25772 9495 25828
rect 9551 25772 9619 25828
rect 9675 25772 9743 25828
rect 9799 25772 9867 25828
rect 9923 25772 9991 25828
rect 10047 25772 10115 25828
rect 10171 25772 10239 25828
rect 10295 25772 10363 25828
rect 10419 25772 10487 25828
rect 10543 25772 10553 25828
rect 8741 25704 10553 25772
rect 8741 25648 8751 25704
rect 8807 25648 8875 25704
rect 8931 25648 8999 25704
rect 9055 25648 9123 25704
rect 9179 25648 9247 25704
rect 9303 25648 9371 25704
rect 9427 25648 9495 25704
rect 9551 25648 9619 25704
rect 9675 25648 9743 25704
rect 9799 25648 9867 25704
rect 9923 25648 9991 25704
rect 10047 25648 10115 25704
rect 10171 25648 10239 25704
rect 10295 25648 10363 25704
rect 10419 25648 10487 25704
rect 10543 25648 10553 25704
rect 8741 25638 10553 25648
rect 12842 26944 13910 26954
rect 12842 26888 12852 26944
rect 12908 26888 12976 26944
rect 13032 26888 13100 26944
rect 13156 26888 13224 26944
rect 13280 26888 13348 26944
rect 13404 26888 13472 26944
rect 13528 26888 13596 26944
rect 13652 26888 13720 26944
rect 13776 26888 13844 26944
rect 13900 26888 13910 26944
rect 12842 26820 13910 26888
rect 12842 26764 12852 26820
rect 12908 26764 12976 26820
rect 13032 26764 13100 26820
rect 13156 26764 13224 26820
rect 13280 26764 13348 26820
rect 13404 26764 13472 26820
rect 13528 26764 13596 26820
rect 13652 26764 13720 26820
rect 13776 26764 13844 26820
rect 13900 26764 13910 26820
rect 12842 26696 13910 26764
rect 12842 26640 12852 26696
rect 12908 26640 12976 26696
rect 13032 26640 13100 26696
rect 13156 26640 13224 26696
rect 13280 26640 13348 26696
rect 13404 26640 13472 26696
rect 13528 26640 13596 26696
rect 13652 26640 13720 26696
rect 13776 26640 13844 26696
rect 13900 26640 13910 26696
rect 12842 26572 13910 26640
rect 12842 26516 12852 26572
rect 12908 26516 12976 26572
rect 13032 26516 13100 26572
rect 13156 26516 13224 26572
rect 13280 26516 13348 26572
rect 13404 26516 13472 26572
rect 13528 26516 13596 26572
rect 13652 26516 13720 26572
rect 13776 26516 13844 26572
rect 13900 26516 13910 26572
rect 12842 26448 13910 26516
rect 12842 26392 12852 26448
rect 12908 26392 12976 26448
rect 13032 26392 13100 26448
rect 13156 26392 13224 26448
rect 13280 26392 13348 26448
rect 13404 26392 13472 26448
rect 13528 26392 13596 26448
rect 13652 26392 13720 26448
rect 13776 26392 13844 26448
rect 13900 26392 13910 26448
rect 12842 26324 13910 26392
rect 12842 26268 12852 26324
rect 12908 26268 12976 26324
rect 13032 26268 13100 26324
rect 13156 26268 13224 26324
rect 13280 26268 13348 26324
rect 13404 26268 13472 26324
rect 13528 26268 13596 26324
rect 13652 26268 13720 26324
rect 13776 26268 13844 26324
rect 13900 26268 13910 26324
rect 12842 26200 13910 26268
rect 12842 26144 12852 26200
rect 12908 26144 12976 26200
rect 13032 26144 13100 26200
rect 13156 26144 13224 26200
rect 13280 26144 13348 26200
rect 13404 26144 13472 26200
rect 13528 26144 13596 26200
rect 13652 26144 13720 26200
rect 13776 26144 13844 26200
rect 13900 26144 13910 26200
rect 12842 26076 13910 26144
rect 12842 26020 12852 26076
rect 12908 26020 12976 26076
rect 13032 26020 13100 26076
rect 13156 26020 13224 26076
rect 13280 26020 13348 26076
rect 13404 26020 13472 26076
rect 13528 26020 13596 26076
rect 13652 26020 13720 26076
rect 13776 26020 13844 26076
rect 13900 26020 13910 26076
rect 12842 25952 13910 26020
rect 12842 25896 12852 25952
rect 12908 25896 12976 25952
rect 13032 25896 13100 25952
rect 13156 25896 13224 25952
rect 13280 25896 13348 25952
rect 13404 25896 13472 25952
rect 13528 25896 13596 25952
rect 13652 25896 13720 25952
rect 13776 25896 13844 25952
rect 13900 25896 13910 25952
rect 12842 25828 13910 25896
rect 12842 25772 12852 25828
rect 12908 25772 12976 25828
rect 13032 25772 13100 25828
rect 13156 25772 13224 25828
rect 13280 25772 13348 25828
rect 13404 25772 13472 25828
rect 13528 25772 13596 25828
rect 13652 25772 13720 25828
rect 13776 25772 13844 25828
rect 13900 25772 13910 25828
rect 12842 25704 13910 25772
rect 12842 25648 12852 25704
rect 12908 25648 12976 25704
rect 13032 25648 13100 25704
rect 13156 25648 13224 25704
rect 13280 25648 13348 25704
rect 13404 25648 13472 25704
rect 13528 25648 13596 25704
rect 13652 25648 13720 25704
rect 13776 25648 13844 25704
rect 13900 25648 13910 25704
rect 12842 25638 13910 25648
rect 1068 25350 2136 25360
rect 1068 25294 1078 25350
rect 1134 25294 1202 25350
rect 1258 25294 1326 25350
rect 1382 25294 1450 25350
rect 1506 25294 1574 25350
rect 1630 25294 1698 25350
rect 1754 25294 1822 25350
rect 1878 25294 1946 25350
rect 2002 25294 2070 25350
rect 2126 25294 2136 25350
rect 1068 25226 2136 25294
rect 1068 25170 1078 25226
rect 1134 25170 1202 25226
rect 1258 25170 1326 25226
rect 1382 25170 1450 25226
rect 1506 25170 1574 25226
rect 1630 25170 1698 25226
rect 1754 25170 1822 25226
rect 1878 25170 1946 25226
rect 2002 25170 2070 25226
rect 2126 25170 2136 25226
rect 1068 25102 2136 25170
rect 1068 25046 1078 25102
rect 1134 25046 1202 25102
rect 1258 25046 1326 25102
rect 1382 25046 1450 25102
rect 1506 25046 1574 25102
rect 1630 25046 1698 25102
rect 1754 25046 1822 25102
rect 1878 25046 1946 25102
rect 2002 25046 2070 25102
rect 2126 25046 2136 25102
rect 1068 24978 2136 25046
rect 1068 24922 1078 24978
rect 1134 24922 1202 24978
rect 1258 24922 1326 24978
rect 1382 24922 1450 24978
rect 1506 24922 1574 24978
rect 1630 24922 1698 24978
rect 1754 24922 1822 24978
rect 1878 24922 1946 24978
rect 2002 24922 2070 24978
rect 2126 24922 2136 24978
rect 1068 24854 2136 24922
rect 1068 24798 1078 24854
rect 1134 24798 1202 24854
rect 1258 24798 1326 24854
rect 1382 24798 1450 24854
rect 1506 24798 1574 24854
rect 1630 24798 1698 24854
rect 1754 24798 1822 24854
rect 1878 24798 1946 24854
rect 2002 24798 2070 24854
rect 2126 24798 2136 24854
rect 1068 24730 2136 24798
rect 1068 24674 1078 24730
rect 1134 24674 1202 24730
rect 1258 24674 1326 24730
rect 1382 24674 1450 24730
rect 1506 24674 1574 24730
rect 1630 24674 1698 24730
rect 1754 24674 1822 24730
rect 1878 24674 1946 24730
rect 2002 24674 2070 24730
rect 2126 24674 2136 24730
rect 1068 24606 2136 24674
rect 1068 24550 1078 24606
rect 1134 24550 1202 24606
rect 1258 24550 1326 24606
rect 1382 24550 1450 24606
rect 1506 24550 1574 24606
rect 1630 24550 1698 24606
rect 1754 24550 1822 24606
rect 1878 24550 1946 24606
rect 2002 24550 2070 24606
rect 2126 24550 2136 24606
rect 1068 24482 2136 24550
rect 1068 24426 1078 24482
rect 1134 24426 1202 24482
rect 1258 24426 1326 24482
rect 1382 24426 1450 24482
rect 1506 24426 1574 24482
rect 1630 24426 1698 24482
rect 1754 24426 1822 24482
rect 1878 24426 1946 24482
rect 2002 24426 2070 24482
rect 2126 24426 2136 24482
rect 1068 24358 2136 24426
rect 1068 24302 1078 24358
rect 1134 24302 1202 24358
rect 1258 24302 1326 24358
rect 1382 24302 1450 24358
rect 1506 24302 1574 24358
rect 1630 24302 1698 24358
rect 1754 24302 1822 24358
rect 1878 24302 1946 24358
rect 2002 24302 2070 24358
rect 2126 24302 2136 24358
rect 1068 24234 2136 24302
rect 1068 24178 1078 24234
rect 1134 24178 1202 24234
rect 1258 24178 1326 24234
rect 1382 24178 1450 24234
rect 1506 24178 1574 24234
rect 1630 24178 1698 24234
rect 1754 24178 1822 24234
rect 1878 24178 1946 24234
rect 2002 24178 2070 24234
rect 2126 24178 2136 24234
rect 1068 24110 2136 24178
rect 1068 24054 1078 24110
rect 1134 24054 1202 24110
rect 1258 24054 1326 24110
rect 1382 24054 1450 24110
rect 1506 24054 1574 24110
rect 1630 24054 1698 24110
rect 1754 24054 1822 24110
rect 1878 24054 1946 24110
rect 2002 24054 2070 24110
rect 2126 24054 2136 24110
rect 1068 23986 2136 24054
rect 1068 23930 1078 23986
rect 1134 23930 1202 23986
rect 1258 23930 1326 23986
rect 1382 23930 1450 23986
rect 1506 23930 1574 23986
rect 1630 23930 1698 23986
rect 1754 23930 1822 23986
rect 1878 23930 1946 23986
rect 2002 23930 2070 23986
rect 2126 23930 2136 23986
rect 1068 23862 2136 23930
rect 1068 23806 1078 23862
rect 1134 23806 1202 23862
rect 1258 23806 1326 23862
rect 1382 23806 1450 23862
rect 1506 23806 1574 23862
rect 1630 23806 1698 23862
rect 1754 23806 1822 23862
rect 1878 23806 1946 23862
rect 2002 23806 2070 23862
rect 2126 23806 2136 23862
rect 1068 23738 2136 23806
rect 1068 23682 1078 23738
rect 1134 23682 1202 23738
rect 1258 23682 1326 23738
rect 1382 23682 1450 23738
rect 1506 23682 1574 23738
rect 1630 23682 1698 23738
rect 1754 23682 1822 23738
rect 1878 23682 1946 23738
rect 2002 23682 2070 23738
rect 2126 23682 2136 23738
rect 1068 23614 2136 23682
rect 1068 23558 1078 23614
rect 1134 23558 1202 23614
rect 1258 23558 1326 23614
rect 1382 23558 1450 23614
rect 1506 23558 1574 23614
rect 1630 23558 1698 23614
rect 1754 23558 1822 23614
rect 1878 23558 1946 23614
rect 2002 23558 2070 23614
rect 2126 23558 2136 23614
rect 1068 23490 2136 23558
rect 1068 23434 1078 23490
rect 1134 23434 1202 23490
rect 1258 23434 1326 23490
rect 1382 23434 1450 23490
rect 1506 23434 1574 23490
rect 1630 23434 1698 23490
rect 1754 23434 1822 23490
rect 1878 23434 1946 23490
rect 2002 23434 2070 23490
rect 2126 23434 2136 23490
rect 1068 23366 2136 23434
rect 1068 23310 1078 23366
rect 1134 23310 1202 23366
rect 1258 23310 1326 23366
rect 1382 23310 1450 23366
rect 1506 23310 1574 23366
rect 1630 23310 1698 23366
rect 1754 23310 1822 23366
rect 1878 23310 1946 23366
rect 2002 23310 2070 23366
rect 2126 23310 2136 23366
rect 1068 23242 2136 23310
rect 1068 23186 1078 23242
rect 1134 23186 1202 23242
rect 1258 23186 1326 23242
rect 1382 23186 1450 23242
rect 1506 23186 1574 23242
rect 1630 23186 1698 23242
rect 1754 23186 1822 23242
rect 1878 23186 1946 23242
rect 2002 23186 2070 23242
rect 2126 23186 2136 23242
rect 1068 23118 2136 23186
rect 1068 23062 1078 23118
rect 1134 23062 1202 23118
rect 1258 23062 1326 23118
rect 1382 23062 1450 23118
rect 1506 23062 1574 23118
rect 1630 23062 1698 23118
rect 1754 23062 1822 23118
rect 1878 23062 1946 23118
rect 2002 23062 2070 23118
rect 2126 23062 2136 23118
rect 1068 22994 2136 23062
rect 1068 22938 1078 22994
rect 1134 22938 1202 22994
rect 1258 22938 1326 22994
rect 1382 22938 1450 22994
rect 1506 22938 1574 22994
rect 1630 22938 1698 22994
rect 1754 22938 1822 22994
rect 1878 22938 1946 22994
rect 2002 22938 2070 22994
rect 2126 22938 2136 22994
rect 1068 22870 2136 22938
rect 1068 22814 1078 22870
rect 1134 22814 1202 22870
rect 1258 22814 1326 22870
rect 1382 22814 1450 22870
rect 1506 22814 1574 22870
rect 1630 22814 1698 22870
rect 1754 22814 1822 22870
rect 1878 22814 1946 22870
rect 2002 22814 2070 22870
rect 2126 22814 2136 22870
rect 1068 22746 2136 22814
rect 1068 22690 1078 22746
rect 1134 22690 1202 22746
rect 1258 22690 1326 22746
rect 1382 22690 1450 22746
rect 1506 22690 1574 22746
rect 1630 22690 1698 22746
rect 1754 22690 1822 22746
rect 1878 22690 1946 22746
rect 2002 22690 2070 22746
rect 2126 22690 2136 22746
rect 1068 22622 2136 22690
rect 1068 22566 1078 22622
rect 1134 22566 1202 22622
rect 1258 22566 1326 22622
rect 1382 22566 1450 22622
rect 1506 22566 1574 22622
rect 1630 22566 1698 22622
rect 1754 22566 1822 22622
rect 1878 22566 1946 22622
rect 2002 22566 2070 22622
rect 2126 22566 2136 22622
rect 1068 22498 2136 22566
rect 1068 22442 1078 22498
rect 1134 22442 1202 22498
rect 1258 22442 1326 22498
rect 1382 22442 1450 22498
rect 1506 22442 1574 22498
rect 1630 22442 1698 22498
rect 1754 22442 1822 22498
rect 1878 22442 1946 22498
rect 2002 22442 2070 22498
rect 2126 22442 2136 22498
rect 1068 22432 2136 22442
rect 4425 25350 6237 25360
rect 4425 25294 4435 25350
rect 4491 25294 4559 25350
rect 4615 25294 4683 25350
rect 4739 25294 4807 25350
rect 4863 25294 4931 25350
rect 4987 25294 5055 25350
rect 5111 25294 5179 25350
rect 5235 25294 5303 25350
rect 5359 25294 5427 25350
rect 5483 25294 5551 25350
rect 5607 25294 5675 25350
rect 5731 25294 5799 25350
rect 5855 25294 5923 25350
rect 5979 25294 6047 25350
rect 6103 25294 6171 25350
rect 6227 25294 6237 25350
rect 4425 25226 6237 25294
rect 4425 25170 4435 25226
rect 4491 25170 4559 25226
rect 4615 25170 4683 25226
rect 4739 25170 4807 25226
rect 4863 25170 4931 25226
rect 4987 25170 5055 25226
rect 5111 25170 5179 25226
rect 5235 25170 5303 25226
rect 5359 25170 5427 25226
rect 5483 25170 5551 25226
rect 5607 25170 5675 25226
rect 5731 25170 5799 25226
rect 5855 25170 5923 25226
rect 5979 25170 6047 25226
rect 6103 25170 6171 25226
rect 6227 25170 6237 25226
rect 4425 25102 6237 25170
rect 4425 25046 4435 25102
rect 4491 25046 4559 25102
rect 4615 25046 4683 25102
rect 4739 25046 4807 25102
rect 4863 25046 4931 25102
rect 4987 25046 5055 25102
rect 5111 25046 5179 25102
rect 5235 25046 5303 25102
rect 5359 25046 5427 25102
rect 5483 25046 5551 25102
rect 5607 25046 5675 25102
rect 5731 25046 5799 25102
rect 5855 25046 5923 25102
rect 5979 25046 6047 25102
rect 6103 25046 6171 25102
rect 6227 25046 6237 25102
rect 4425 24978 6237 25046
rect 4425 24922 4435 24978
rect 4491 24922 4559 24978
rect 4615 24922 4683 24978
rect 4739 24922 4807 24978
rect 4863 24922 4931 24978
rect 4987 24922 5055 24978
rect 5111 24922 5179 24978
rect 5235 24922 5303 24978
rect 5359 24922 5427 24978
rect 5483 24922 5551 24978
rect 5607 24922 5675 24978
rect 5731 24922 5799 24978
rect 5855 24922 5923 24978
rect 5979 24922 6047 24978
rect 6103 24922 6171 24978
rect 6227 24922 6237 24978
rect 4425 24854 6237 24922
rect 4425 24798 4435 24854
rect 4491 24798 4559 24854
rect 4615 24798 4683 24854
rect 4739 24798 4807 24854
rect 4863 24798 4931 24854
rect 4987 24798 5055 24854
rect 5111 24798 5179 24854
rect 5235 24798 5303 24854
rect 5359 24798 5427 24854
rect 5483 24798 5551 24854
rect 5607 24798 5675 24854
rect 5731 24798 5799 24854
rect 5855 24798 5923 24854
rect 5979 24798 6047 24854
rect 6103 24798 6171 24854
rect 6227 24798 6237 24854
rect 4425 24730 6237 24798
rect 4425 24674 4435 24730
rect 4491 24674 4559 24730
rect 4615 24674 4683 24730
rect 4739 24674 4807 24730
rect 4863 24674 4931 24730
rect 4987 24674 5055 24730
rect 5111 24674 5179 24730
rect 5235 24674 5303 24730
rect 5359 24674 5427 24730
rect 5483 24674 5551 24730
rect 5607 24674 5675 24730
rect 5731 24674 5799 24730
rect 5855 24674 5923 24730
rect 5979 24674 6047 24730
rect 6103 24674 6171 24730
rect 6227 24674 6237 24730
rect 4425 24606 6237 24674
rect 4425 24550 4435 24606
rect 4491 24550 4559 24606
rect 4615 24550 4683 24606
rect 4739 24550 4807 24606
rect 4863 24550 4931 24606
rect 4987 24550 5055 24606
rect 5111 24550 5179 24606
rect 5235 24550 5303 24606
rect 5359 24550 5427 24606
rect 5483 24550 5551 24606
rect 5607 24550 5675 24606
rect 5731 24550 5799 24606
rect 5855 24550 5923 24606
rect 5979 24550 6047 24606
rect 6103 24550 6171 24606
rect 6227 24550 6237 24606
rect 4425 24482 6237 24550
rect 4425 24426 4435 24482
rect 4491 24426 4559 24482
rect 4615 24426 4683 24482
rect 4739 24426 4807 24482
rect 4863 24426 4931 24482
rect 4987 24426 5055 24482
rect 5111 24426 5179 24482
rect 5235 24426 5303 24482
rect 5359 24426 5427 24482
rect 5483 24426 5551 24482
rect 5607 24426 5675 24482
rect 5731 24426 5799 24482
rect 5855 24426 5923 24482
rect 5979 24426 6047 24482
rect 6103 24426 6171 24482
rect 6227 24426 6237 24482
rect 4425 24358 6237 24426
rect 4425 24302 4435 24358
rect 4491 24302 4559 24358
rect 4615 24302 4683 24358
rect 4739 24302 4807 24358
rect 4863 24302 4931 24358
rect 4987 24302 5055 24358
rect 5111 24302 5179 24358
rect 5235 24302 5303 24358
rect 5359 24302 5427 24358
rect 5483 24302 5551 24358
rect 5607 24302 5675 24358
rect 5731 24302 5799 24358
rect 5855 24302 5923 24358
rect 5979 24302 6047 24358
rect 6103 24302 6171 24358
rect 6227 24302 6237 24358
rect 4425 24234 6237 24302
rect 4425 24178 4435 24234
rect 4491 24178 4559 24234
rect 4615 24178 4683 24234
rect 4739 24178 4807 24234
rect 4863 24178 4931 24234
rect 4987 24178 5055 24234
rect 5111 24178 5179 24234
rect 5235 24178 5303 24234
rect 5359 24178 5427 24234
rect 5483 24178 5551 24234
rect 5607 24178 5675 24234
rect 5731 24178 5799 24234
rect 5855 24178 5923 24234
rect 5979 24178 6047 24234
rect 6103 24178 6171 24234
rect 6227 24178 6237 24234
rect 4425 24110 6237 24178
rect 4425 24054 4435 24110
rect 4491 24054 4559 24110
rect 4615 24054 4683 24110
rect 4739 24054 4807 24110
rect 4863 24054 4931 24110
rect 4987 24054 5055 24110
rect 5111 24054 5179 24110
rect 5235 24054 5303 24110
rect 5359 24054 5427 24110
rect 5483 24054 5551 24110
rect 5607 24054 5675 24110
rect 5731 24054 5799 24110
rect 5855 24054 5923 24110
rect 5979 24054 6047 24110
rect 6103 24054 6171 24110
rect 6227 24054 6237 24110
rect 4425 23986 6237 24054
rect 4425 23930 4435 23986
rect 4491 23930 4559 23986
rect 4615 23930 4683 23986
rect 4739 23930 4807 23986
rect 4863 23930 4931 23986
rect 4987 23930 5055 23986
rect 5111 23930 5179 23986
rect 5235 23930 5303 23986
rect 5359 23930 5427 23986
rect 5483 23930 5551 23986
rect 5607 23930 5675 23986
rect 5731 23930 5799 23986
rect 5855 23930 5923 23986
rect 5979 23930 6047 23986
rect 6103 23930 6171 23986
rect 6227 23930 6237 23986
rect 4425 23862 6237 23930
rect 4425 23806 4435 23862
rect 4491 23806 4559 23862
rect 4615 23806 4683 23862
rect 4739 23806 4807 23862
rect 4863 23806 4931 23862
rect 4987 23806 5055 23862
rect 5111 23806 5179 23862
rect 5235 23806 5303 23862
rect 5359 23806 5427 23862
rect 5483 23806 5551 23862
rect 5607 23806 5675 23862
rect 5731 23806 5799 23862
rect 5855 23806 5923 23862
rect 5979 23806 6047 23862
rect 6103 23806 6171 23862
rect 6227 23806 6237 23862
rect 4425 23738 6237 23806
rect 4425 23682 4435 23738
rect 4491 23682 4559 23738
rect 4615 23682 4683 23738
rect 4739 23682 4807 23738
rect 4863 23682 4931 23738
rect 4987 23682 5055 23738
rect 5111 23682 5179 23738
rect 5235 23682 5303 23738
rect 5359 23682 5427 23738
rect 5483 23682 5551 23738
rect 5607 23682 5675 23738
rect 5731 23682 5799 23738
rect 5855 23682 5923 23738
rect 5979 23682 6047 23738
rect 6103 23682 6171 23738
rect 6227 23682 6237 23738
rect 4425 23614 6237 23682
rect 4425 23558 4435 23614
rect 4491 23558 4559 23614
rect 4615 23558 4683 23614
rect 4739 23558 4807 23614
rect 4863 23558 4931 23614
rect 4987 23558 5055 23614
rect 5111 23558 5179 23614
rect 5235 23558 5303 23614
rect 5359 23558 5427 23614
rect 5483 23558 5551 23614
rect 5607 23558 5675 23614
rect 5731 23558 5799 23614
rect 5855 23558 5923 23614
rect 5979 23558 6047 23614
rect 6103 23558 6171 23614
rect 6227 23558 6237 23614
rect 4425 23490 6237 23558
rect 4425 23434 4435 23490
rect 4491 23434 4559 23490
rect 4615 23434 4683 23490
rect 4739 23434 4807 23490
rect 4863 23434 4931 23490
rect 4987 23434 5055 23490
rect 5111 23434 5179 23490
rect 5235 23434 5303 23490
rect 5359 23434 5427 23490
rect 5483 23434 5551 23490
rect 5607 23434 5675 23490
rect 5731 23434 5799 23490
rect 5855 23434 5923 23490
rect 5979 23434 6047 23490
rect 6103 23434 6171 23490
rect 6227 23434 6237 23490
rect 4425 23366 6237 23434
rect 4425 23310 4435 23366
rect 4491 23310 4559 23366
rect 4615 23310 4683 23366
rect 4739 23310 4807 23366
rect 4863 23310 4931 23366
rect 4987 23310 5055 23366
rect 5111 23310 5179 23366
rect 5235 23310 5303 23366
rect 5359 23310 5427 23366
rect 5483 23310 5551 23366
rect 5607 23310 5675 23366
rect 5731 23310 5799 23366
rect 5855 23310 5923 23366
rect 5979 23310 6047 23366
rect 6103 23310 6171 23366
rect 6227 23310 6237 23366
rect 4425 23242 6237 23310
rect 4425 23186 4435 23242
rect 4491 23186 4559 23242
rect 4615 23186 4683 23242
rect 4739 23186 4807 23242
rect 4863 23186 4931 23242
rect 4987 23186 5055 23242
rect 5111 23186 5179 23242
rect 5235 23186 5303 23242
rect 5359 23186 5427 23242
rect 5483 23186 5551 23242
rect 5607 23186 5675 23242
rect 5731 23186 5799 23242
rect 5855 23186 5923 23242
rect 5979 23186 6047 23242
rect 6103 23186 6171 23242
rect 6227 23186 6237 23242
rect 4425 23118 6237 23186
rect 4425 23062 4435 23118
rect 4491 23062 4559 23118
rect 4615 23062 4683 23118
rect 4739 23062 4807 23118
rect 4863 23062 4931 23118
rect 4987 23062 5055 23118
rect 5111 23062 5179 23118
rect 5235 23062 5303 23118
rect 5359 23062 5427 23118
rect 5483 23062 5551 23118
rect 5607 23062 5675 23118
rect 5731 23062 5799 23118
rect 5855 23062 5923 23118
rect 5979 23062 6047 23118
rect 6103 23062 6171 23118
rect 6227 23062 6237 23118
rect 4425 22994 6237 23062
rect 4425 22938 4435 22994
rect 4491 22938 4559 22994
rect 4615 22938 4683 22994
rect 4739 22938 4807 22994
rect 4863 22938 4931 22994
rect 4987 22938 5055 22994
rect 5111 22938 5179 22994
rect 5235 22938 5303 22994
rect 5359 22938 5427 22994
rect 5483 22938 5551 22994
rect 5607 22938 5675 22994
rect 5731 22938 5799 22994
rect 5855 22938 5923 22994
rect 5979 22938 6047 22994
rect 6103 22938 6171 22994
rect 6227 22938 6237 22994
rect 4425 22870 6237 22938
rect 4425 22814 4435 22870
rect 4491 22814 4559 22870
rect 4615 22814 4683 22870
rect 4739 22814 4807 22870
rect 4863 22814 4931 22870
rect 4987 22814 5055 22870
rect 5111 22814 5179 22870
rect 5235 22814 5303 22870
rect 5359 22814 5427 22870
rect 5483 22814 5551 22870
rect 5607 22814 5675 22870
rect 5731 22814 5799 22870
rect 5855 22814 5923 22870
rect 5979 22814 6047 22870
rect 6103 22814 6171 22870
rect 6227 22814 6237 22870
rect 4425 22746 6237 22814
rect 4425 22690 4435 22746
rect 4491 22690 4559 22746
rect 4615 22690 4683 22746
rect 4739 22690 4807 22746
rect 4863 22690 4931 22746
rect 4987 22690 5055 22746
rect 5111 22690 5179 22746
rect 5235 22690 5303 22746
rect 5359 22690 5427 22746
rect 5483 22690 5551 22746
rect 5607 22690 5675 22746
rect 5731 22690 5799 22746
rect 5855 22690 5923 22746
rect 5979 22690 6047 22746
rect 6103 22690 6171 22746
rect 6227 22690 6237 22746
rect 4425 22622 6237 22690
rect 4425 22566 4435 22622
rect 4491 22566 4559 22622
rect 4615 22566 4683 22622
rect 4739 22566 4807 22622
rect 4863 22566 4931 22622
rect 4987 22566 5055 22622
rect 5111 22566 5179 22622
rect 5235 22566 5303 22622
rect 5359 22566 5427 22622
rect 5483 22566 5551 22622
rect 5607 22566 5675 22622
rect 5731 22566 5799 22622
rect 5855 22566 5923 22622
rect 5979 22566 6047 22622
rect 6103 22566 6171 22622
rect 6227 22566 6237 22622
rect 4425 22498 6237 22566
rect 4425 22442 4435 22498
rect 4491 22442 4559 22498
rect 4615 22442 4683 22498
rect 4739 22442 4807 22498
rect 4863 22442 4931 22498
rect 4987 22442 5055 22498
rect 5111 22442 5179 22498
rect 5235 22442 5303 22498
rect 5359 22442 5427 22498
rect 5483 22442 5551 22498
rect 5607 22442 5675 22498
rect 5731 22442 5799 22498
rect 5855 22442 5923 22498
rect 5979 22442 6047 22498
rect 6103 22442 6171 22498
rect 6227 22442 6237 22498
rect 4425 22432 6237 22442
rect 7552 25350 8620 25360
rect 7552 25294 7562 25350
rect 7618 25294 7686 25350
rect 7742 25294 7810 25350
rect 7866 25294 7934 25350
rect 7990 25294 8058 25350
rect 8114 25294 8182 25350
rect 8238 25294 8306 25350
rect 8362 25294 8430 25350
rect 8486 25294 8554 25350
rect 8610 25294 8620 25350
rect 7552 25226 8620 25294
rect 7552 25170 7562 25226
rect 7618 25170 7686 25226
rect 7742 25170 7810 25226
rect 7866 25170 7934 25226
rect 7990 25170 8058 25226
rect 8114 25170 8182 25226
rect 8238 25170 8306 25226
rect 8362 25170 8430 25226
rect 8486 25170 8554 25226
rect 8610 25170 8620 25226
rect 7552 25102 8620 25170
rect 7552 25046 7562 25102
rect 7618 25046 7686 25102
rect 7742 25046 7810 25102
rect 7866 25046 7934 25102
rect 7990 25046 8058 25102
rect 8114 25046 8182 25102
rect 8238 25046 8306 25102
rect 8362 25046 8430 25102
rect 8486 25046 8554 25102
rect 8610 25046 8620 25102
rect 7552 24978 8620 25046
rect 7552 24922 7562 24978
rect 7618 24922 7686 24978
rect 7742 24922 7810 24978
rect 7866 24922 7934 24978
rect 7990 24922 8058 24978
rect 8114 24922 8182 24978
rect 8238 24922 8306 24978
rect 8362 24922 8430 24978
rect 8486 24922 8554 24978
rect 8610 24922 8620 24978
rect 7552 24854 8620 24922
rect 7552 24798 7562 24854
rect 7618 24798 7686 24854
rect 7742 24798 7810 24854
rect 7866 24798 7934 24854
rect 7990 24798 8058 24854
rect 8114 24798 8182 24854
rect 8238 24798 8306 24854
rect 8362 24798 8430 24854
rect 8486 24798 8554 24854
rect 8610 24798 8620 24854
rect 7552 24730 8620 24798
rect 7552 24674 7562 24730
rect 7618 24674 7686 24730
rect 7742 24674 7810 24730
rect 7866 24674 7934 24730
rect 7990 24674 8058 24730
rect 8114 24674 8182 24730
rect 8238 24674 8306 24730
rect 8362 24674 8430 24730
rect 8486 24674 8554 24730
rect 8610 24674 8620 24730
rect 7552 24606 8620 24674
rect 7552 24550 7562 24606
rect 7618 24550 7686 24606
rect 7742 24550 7810 24606
rect 7866 24550 7934 24606
rect 7990 24550 8058 24606
rect 8114 24550 8182 24606
rect 8238 24550 8306 24606
rect 8362 24550 8430 24606
rect 8486 24550 8554 24606
rect 8610 24550 8620 24606
rect 7552 24482 8620 24550
rect 7552 24426 7562 24482
rect 7618 24426 7686 24482
rect 7742 24426 7810 24482
rect 7866 24426 7934 24482
rect 7990 24426 8058 24482
rect 8114 24426 8182 24482
rect 8238 24426 8306 24482
rect 8362 24426 8430 24482
rect 8486 24426 8554 24482
rect 8610 24426 8620 24482
rect 7552 24358 8620 24426
rect 7552 24302 7562 24358
rect 7618 24302 7686 24358
rect 7742 24302 7810 24358
rect 7866 24302 7934 24358
rect 7990 24302 8058 24358
rect 8114 24302 8182 24358
rect 8238 24302 8306 24358
rect 8362 24302 8430 24358
rect 8486 24302 8554 24358
rect 8610 24302 8620 24358
rect 7552 24234 8620 24302
rect 7552 24178 7562 24234
rect 7618 24178 7686 24234
rect 7742 24178 7810 24234
rect 7866 24178 7934 24234
rect 7990 24178 8058 24234
rect 8114 24178 8182 24234
rect 8238 24178 8306 24234
rect 8362 24178 8430 24234
rect 8486 24178 8554 24234
rect 8610 24178 8620 24234
rect 7552 24110 8620 24178
rect 7552 24054 7562 24110
rect 7618 24054 7686 24110
rect 7742 24054 7810 24110
rect 7866 24054 7934 24110
rect 7990 24054 8058 24110
rect 8114 24054 8182 24110
rect 8238 24054 8306 24110
rect 8362 24054 8430 24110
rect 8486 24054 8554 24110
rect 8610 24054 8620 24110
rect 7552 23986 8620 24054
rect 7552 23930 7562 23986
rect 7618 23930 7686 23986
rect 7742 23930 7810 23986
rect 7866 23930 7934 23986
rect 7990 23930 8058 23986
rect 8114 23930 8182 23986
rect 8238 23930 8306 23986
rect 8362 23930 8430 23986
rect 8486 23930 8554 23986
rect 8610 23930 8620 23986
rect 7552 23862 8620 23930
rect 7552 23806 7562 23862
rect 7618 23806 7686 23862
rect 7742 23806 7810 23862
rect 7866 23806 7934 23862
rect 7990 23806 8058 23862
rect 8114 23806 8182 23862
rect 8238 23806 8306 23862
rect 8362 23806 8430 23862
rect 8486 23806 8554 23862
rect 8610 23806 8620 23862
rect 7552 23738 8620 23806
rect 7552 23682 7562 23738
rect 7618 23682 7686 23738
rect 7742 23682 7810 23738
rect 7866 23682 7934 23738
rect 7990 23682 8058 23738
rect 8114 23682 8182 23738
rect 8238 23682 8306 23738
rect 8362 23682 8430 23738
rect 8486 23682 8554 23738
rect 8610 23682 8620 23738
rect 7552 23614 8620 23682
rect 7552 23558 7562 23614
rect 7618 23558 7686 23614
rect 7742 23558 7810 23614
rect 7866 23558 7934 23614
rect 7990 23558 8058 23614
rect 8114 23558 8182 23614
rect 8238 23558 8306 23614
rect 8362 23558 8430 23614
rect 8486 23558 8554 23614
rect 8610 23558 8620 23614
rect 7552 23490 8620 23558
rect 7552 23434 7562 23490
rect 7618 23434 7686 23490
rect 7742 23434 7810 23490
rect 7866 23434 7934 23490
rect 7990 23434 8058 23490
rect 8114 23434 8182 23490
rect 8238 23434 8306 23490
rect 8362 23434 8430 23490
rect 8486 23434 8554 23490
rect 8610 23434 8620 23490
rect 7552 23366 8620 23434
rect 7552 23310 7562 23366
rect 7618 23310 7686 23366
rect 7742 23310 7810 23366
rect 7866 23310 7934 23366
rect 7990 23310 8058 23366
rect 8114 23310 8182 23366
rect 8238 23310 8306 23366
rect 8362 23310 8430 23366
rect 8486 23310 8554 23366
rect 8610 23310 8620 23366
rect 7552 23242 8620 23310
rect 7552 23186 7562 23242
rect 7618 23186 7686 23242
rect 7742 23186 7810 23242
rect 7866 23186 7934 23242
rect 7990 23186 8058 23242
rect 8114 23186 8182 23242
rect 8238 23186 8306 23242
rect 8362 23186 8430 23242
rect 8486 23186 8554 23242
rect 8610 23186 8620 23242
rect 7552 23118 8620 23186
rect 7552 23062 7562 23118
rect 7618 23062 7686 23118
rect 7742 23062 7810 23118
rect 7866 23062 7934 23118
rect 7990 23062 8058 23118
rect 8114 23062 8182 23118
rect 8238 23062 8306 23118
rect 8362 23062 8430 23118
rect 8486 23062 8554 23118
rect 8610 23062 8620 23118
rect 7552 22994 8620 23062
rect 7552 22938 7562 22994
rect 7618 22938 7686 22994
rect 7742 22938 7810 22994
rect 7866 22938 7934 22994
rect 7990 22938 8058 22994
rect 8114 22938 8182 22994
rect 8238 22938 8306 22994
rect 8362 22938 8430 22994
rect 8486 22938 8554 22994
rect 8610 22938 8620 22994
rect 7552 22870 8620 22938
rect 7552 22814 7562 22870
rect 7618 22814 7686 22870
rect 7742 22814 7810 22870
rect 7866 22814 7934 22870
rect 7990 22814 8058 22870
rect 8114 22814 8182 22870
rect 8238 22814 8306 22870
rect 8362 22814 8430 22870
rect 8486 22814 8554 22870
rect 8610 22814 8620 22870
rect 7552 22746 8620 22814
rect 7552 22690 7562 22746
rect 7618 22690 7686 22746
rect 7742 22690 7810 22746
rect 7866 22690 7934 22746
rect 7990 22690 8058 22746
rect 8114 22690 8182 22746
rect 8238 22690 8306 22746
rect 8362 22690 8430 22746
rect 8486 22690 8554 22746
rect 8610 22690 8620 22746
rect 7552 22622 8620 22690
rect 7552 22566 7562 22622
rect 7618 22566 7686 22622
rect 7742 22566 7810 22622
rect 7866 22566 7934 22622
rect 7990 22566 8058 22622
rect 8114 22566 8182 22622
rect 8238 22566 8306 22622
rect 8362 22566 8430 22622
rect 8486 22566 8554 22622
rect 8610 22566 8620 22622
rect 7552 22498 8620 22566
rect 7552 22442 7562 22498
rect 7618 22442 7686 22498
rect 7742 22442 7810 22498
rect 7866 22442 7934 22498
rect 7990 22442 8058 22498
rect 8114 22442 8182 22498
rect 8238 22442 8306 22498
rect 8362 22442 8430 22498
rect 8486 22442 8554 22498
rect 8610 22442 8620 22498
rect 7552 22432 8620 22442
rect 10669 25350 12481 25360
rect 10669 25294 10679 25350
rect 10735 25294 10803 25350
rect 10859 25294 10927 25350
rect 10983 25294 11051 25350
rect 11107 25294 11175 25350
rect 11231 25294 11299 25350
rect 11355 25294 11423 25350
rect 11479 25294 11547 25350
rect 11603 25294 11671 25350
rect 11727 25294 11795 25350
rect 11851 25294 11919 25350
rect 11975 25294 12043 25350
rect 12099 25294 12167 25350
rect 12223 25294 12291 25350
rect 12347 25294 12415 25350
rect 12471 25294 12481 25350
rect 10669 25226 12481 25294
rect 10669 25170 10679 25226
rect 10735 25170 10803 25226
rect 10859 25170 10927 25226
rect 10983 25170 11051 25226
rect 11107 25170 11175 25226
rect 11231 25170 11299 25226
rect 11355 25170 11423 25226
rect 11479 25170 11547 25226
rect 11603 25170 11671 25226
rect 11727 25170 11795 25226
rect 11851 25170 11919 25226
rect 11975 25170 12043 25226
rect 12099 25170 12167 25226
rect 12223 25170 12291 25226
rect 12347 25170 12415 25226
rect 12471 25170 12481 25226
rect 10669 25102 12481 25170
rect 10669 25046 10679 25102
rect 10735 25046 10803 25102
rect 10859 25046 10927 25102
rect 10983 25046 11051 25102
rect 11107 25046 11175 25102
rect 11231 25046 11299 25102
rect 11355 25046 11423 25102
rect 11479 25046 11547 25102
rect 11603 25046 11671 25102
rect 11727 25046 11795 25102
rect 11851 25046 11919 25102
rect 11975 25046 12043 25102
rect 12099 25046 12167 25102
rect 12223 25046 12291 25102
rect 12347 25046 12415 25102
rect 12471 25046 12481 25102
rect 10669 24978 12481 25046
rect 10669 24922 10679 24978
rect 10735 24922 10803 24978
rect 10859 24922 10927 24978
rect 10983 24922 11051 24978
rect 11107 24922 11175 24978
rect 11231 24922 11299 24978
rect 11355 24922 11423 24978
rect 11479 24922 11547 24978
rect 11603 24922 11671 24978
rect 11727 24922 11795 24978
rect 11851 24922 11919 24978
rect 11975 24922 12043 24978
rect 12099 24922 12167 24978
rect 12223 24922 12291 24978
rect 12347 24922 12415 24978
rect 12471 24922 12481 24978
rect 10669 24854 12481 24922
rect 10669 24798 10679 24854
rect 10735 24798 10803 24854
rect 10859 24798 10927 24854
rect 10983 24798 11051 24854
rect 11107 24798 11175 24854
rect 11231 24798 11299 24854
rect 11355 24798 11423 24854
rect 11479 24798 11547 24854
rect 11603 24798 11671 24854
rect 11727 24798 11795 24854
rect 11851 24798 11919 24854
rect 11975 24798 12043 24854
rect 12099 24798 12167 24854
rect 12223 24798 12291 24854
rect 12347 24798 12415 24854
rect 12471 24798 12481 24854
rect 10669 24730 12481 24798
rect 10669 24674 10679 24730
rect 10735 24674 10803 24730
rect 10859 24674 10927 24730
rect 10983 24674 11051 24730
rect 11107 24674 11175 24730
rect 11231 24674 11299 24730
rect 11355 24674 11423 24730
rect 11479 24674 11547 24730
rect 11603 24674 11671 24730
rect 11727 24674 11795 24730
rect 11851 24674 11919 24730
rect 11975 24674 12043 24730
rect 12099 24674 12167 24730
rect 12223 24674 12291 24730
rect 12347 24674 12415 24730
rect 12471 24674 12481 24730
rect 10669 24606 12481 24674
rect 10669 24550 10679 24606
rect 10735 24550 10803 24606
rect 10859 24550 10927 24606
rect 10983 24550 11051 24606
rect 11107 24550 11175 24606
rect 11231 24550 11299 24606
rect 11355 24550 11423 24606
rect 11479 24550 11547 24606
rect 11603 24550 11671 24606
rect 11727 24550 11795 24606
rect 11851 24550 11919 24606
rect 11975 24550 12043 24606
rect 12099 24550 12167 24606
rect 12223 24550 12291 24606
rect 12347 24550 12415 24606
rect 12471 24550 12481 24606
rect 10669 24482 12481 24550
rect 10669 24426 10679 24482
rect 10735 24426 10803 24482
rect 10859 24426 10927 24482
rect 10983 24426 11051 24482
rect 11107 24426 11175 24482
rect 11231 24426 11299 24482
rect 11355 24426 11423 24482
rect 11479 24426 11547 24482
rect 11603 24426 11671 24482
rect 11727 24426 11795 24482
rect 11851 24426 11919 24482
rect 11975 24426 12043 24482
rect 12099 24426 12167 24482
rect 12223 24426 12291 24482
rect 12347 24426 12415 24482
rect 12471 24426 12481 24482
rect 10669 24358 12481 24426
rect 10669 24302 10679 24358
rect 10735 24302 10803 24358
rect 10859 24302 10927 24358
rect 10983 24302 11051 24358
rect 11107 24302 11175 24358
rect 11231 24302 11299 24358
rect 11355 24302 11423 24358
rect 11479 24302 11547 24358
rect 11603 24302 11671 24358
rect 11727 24302 11795 24358
rect 11851 24302 11919 24358
rect 11975 24302 12043 24358
rect 12099 24302 12167 24358
rect 12223 24302 12291 24358
rect 12347 24302 12415 24358
rect 12471 24302 12481 24358
rect 10669 24234 12481 24302
rect 10669 24178 10679 24234
rect 10735 24178 10803 24234
rect 10859 24178 10927 24234
rect 10983 24178 11051 24234
rect 11107 24178 11175 24234
rect 11231 24178 11299 24234
rect 11355 24178 11423 24234
rect 11479 24178 11547 24234
rect 11603 24178 11671 24234
rect 11727 24178 11795 24234
rect 11851 24178 11919 24234
rect 11975 24178 12043 24234
rect 12099 24178 12167 24234
rect 12223 24178 12291 24234
rect 12347 24178 12415 24234
rect 12471 24178 12481 24234
rect 10669 24110 12481 24178
rect 10669 24054 10679 24110
rect 10735 24054 10803 24110
rect 10859 24054 10927 24110
rect 10983 24054 11051 24110
rect 11107 24054 11175 24110
rect 11231 24054 11299 24110
rect 11355 24054 11423 24110
rect 11479 24054 11547 24110
rect 11603 24054 11671 24110
rect 11727 24054 11795 24110
rect 11851 24054 11919 24110
rect 11975 24054 12043 24110
rect 12099 24054 12167 24110
rect 12223 24054 12291 24110
rect 12347 24054 12415 24110
rect 12471 24054 12481 24110
rect 10669 23986 12481 24054
rect 10669 23930 10679 23986
rect 10735 23930 10803 23986
rect 10859 23930 10927 23986
rect 10983 23930 11051 23986
rect 11107 23930 11175 23986
rect 11231 23930 11299 23986
rect 11355 23930 11423 23986
rect 11479 23930 11547 23986
rect 11603 23930 11671 23986
rect 11727 23930 11795 23986
rect 11851 23930 11919 23986
rect 11975 23930 12043 23986
rect 12099 23930 12167 23986
rect 12223 23930 12291 23986
rect 12347 23930 12415 23986
rect 12471 23930 12481 23986
rect 10669 23862 12481 23930
rect 10669 23806 10679 23862
rect 10735 23806 10803 23862
rect 10859 23806 10927 23862
rect 10983 23806 11051 23862
rect 11107 23806 11175 23862
rect 11231 23806 11299 23862
rect 11355 23806 11423 23862
rect 11479 23806 11547 23862
rect 11603 23806 11671 23862
rect 11727 23806 11795 23862
rect 11851 23806 11919 23862
rect 11975 23806 12043 23862
rect 12099 23806 12167 23862
rect 12223 23806 12291 23862
rect 12347 23806 12415 23862
rect 12471 23806 12481 23862
rect 10669 23738 12481 23806
rect 10669 23682 10679 23738
rect 10735 23682 10803 23738
rect 10859 23682 10927 23738
rect 10983 23682 11051 23738
rect 11107 23682 11175 23738
rect 11231 23682 11299 23738
rect 11355 23682 11423 23738
rect 11479 23682 11547 23738
rect 11603 23682 11671 23738
rect 11727 23682 11795 23738
rect 11851 23682 11919 23738
rect 11975 23682 12043 23738
rect 12099 23682 12167 23738
rect 12223 23682 12291 23738
rect 12347 23682 12415 23738
rect 12471 23682 12481 23738
rect 10669 23614 12481 23682
rect 10669 23558 10679 23614
rect 10735 23558 10803 23614
rect 10859 23558 10927 23614
rect 10983 23558 11051 23614
rect 11107 23558 11175 23614
rect 11231 23558 11299 23614
rect 11355 23558 11423 23614
rect 11479 23558 11547 23614
rect 11603 23558 11671 23614
rect 11727 23558 11795 23614
rect 11851 23558 11919 23614
rect 11975 23558 12043 23614
rect 12099 23558 12167 23614
rect 12223 23558 12291 23614
rect 12347 23558 12415 23614
rect 12471 23558 12481 23614
rect 10669 23490 12481 23558
rect 10669 23434 10679 23490
rect 10735 23434 10803 23490
rect 10859 23434 10927 23490
rect 10983 23434 11051 23490
rect 11107 23434 11175 23490
rect 11231 23434 11299 23490
rect 11355 23434 11423 23490
rect 11479 23434 11547 23490
rect 11603 23434 11671 23490
rect 11727 23434 11795 23490
rect 11851 23434 11919 23490
rect 11975 23434 12043 23490
rect 12099 23434 12167 23490
rect 12223 23434 12291 23490
rect 12347 23434 12415 23490
rect 12471 23434 12481 23490
rect 10669 23366 12481 23434
rect 10669 23310 10679 23366
rect 10735 23310 10803 23366
rect 10859 23310 10927 23366
rect 10983 23310 11051 23366
rect 11107 23310 11175 23366
rect 11231 23310 11299 23366
rect 11355 23310 11423 23366
rect 11479 23310 11547 23366
rect 11603 23310 11671 23366
rect 11727 23310 11795 23366
rect 11851 23310 11919 23366
rect 11975 23310 12043 23366
rect 12099 23310 12167 23366
rect 12223 23310 12291 23366
rect 12347 23310 12415 23366
rect 12471 23310 12481 23366
rect 10669 23242 12481 23310
rect 10669 23186 10679 23242
rect 10735 23186 10803 23242
rect 10859 23186 10927 23242
rect 10983 23186 11051 23242
rect 11107 23186 11175 23242
rect 11231 23186 11299 23242
rect 11355 23186 11423 23242
rect 11479 23186 11547 23242
rect 11603 23186 11671 23242
rect 11727 23186 11795 23242
rect 11851 23186 11919 23242
rect 11975 23186 12043 23242
rect 12099 23186 12167 23242
rect 12223 23186 12291 23242
rect 12347 23186 12415 23242
rect 12471 23186 12481 23242
rect 10669 23118 12481 23186
rect 10669 23062 10679 23118
rect 10735 23062 10803 23118
rect 10859 23062 10927 23118
rect 10983 23062 11051 23118
rect 11107 23062 11175 23118
rect 11231 23062 11299 23118
rect 11355 23062 11423 23118
rect 11479 23062 11547 23118
rect 11603 23062 11671 23118
rect 11727 23062 11795 23118
rect 11851 23062 11919 23118
rect 11975 23062 12043 23118
rect 12099 23062 12167 23118
rect 12223 23062 12291 23118
rect 12347 23062 12415 23118
rect 12471 23062 12481 23118
rect 10669 22994 12481 23062
rect 10669 22938 10679 22994
rect 10735 22938 10803 22994
rect 10859 22938 10927 22994
rect 10983 22938 11051 22994
rect 11107 22938 11175 22994
rect 11231 22938 11299 22994
rect 11355 22938 11423 22994
rect 11479 22938 11547 22994
rect 11603 22938 11671 22994
rect 11727 22938 11795 22994
rect 11851 22938 11919 22994
rect 11975 22938 12043 22994
rect 12099 22938 12167 22994
rect 12223 22938 12291 22994
rect 12347 22938 12415 22994
rect 12471 22938 12481 22994
rect 10669 22870 12481 22938
rect 10669 22814 10679 22870
rect 10735 22814 10803 22870
rect 10859 22814 10927 22870
rect 10983 22814 11051 22870
rect 11107 22814 11175 22870
rect 11231 22814 11299 22870
rect 11355 22814 11423 22870
rect 11479 22814 11547 22870
rect 11603 22814 11671 22870
rect 11727 22814 11795 22870
rect 11851 22814 11919 22870
rect 11975 22814 12043 22870
rect 12099 22814 12167 22870
rect 12223 22814 12291 22870
rect 12347 22814 12415 22870
rect 12471 22814 12481 22870
rect 10669 22746 12481 22814
rect 10669 22690 10679 22746
rect 10735 22690 10803 22746
rect 10859 22690 10927 22746
rect 10983 22690 11051 22746
rect 11107 22690 11175 22746
rect 11231 22690 11299 22746
rect 11355 22690 11423 22746
rect 11479 22690 11547 22746
rect 11603 22690 11671 22746
rect 11727 22690 11795 22746
rect 11851 22690 11919 22746
rect 11975 22690 12043 22746
rect 12099 22690 12167 22746
rect 12223 22690 12291 22746
rect 12347 22690 12415 22746
rect 12471 22690 12481 22746
rect 10669 22622 12481 22690
rect 10669 22566 10679 22622
rect 10735 22566 10803 22622
rect 10859 22566 10927 22622
rect 10983 22566 11051 22622
rect 11107 22566 11175 22622
rect 11231 22566 11299 22622
rect 11355 22566 11423 22622
rect 11479 22566 11547 22622
rect 11603 22566 11671 22622
rect 11727 22566 11795 22622
rect 11851 22566 11919 22622
rect 11975 22566 12043 22622
rect 12099 22566 12167 22622
rect 12223 22566 12291 22622
rect 12347 22566 12415 22622
rect 12471 22566 12481 22622
rect 10669 22498 12481 22566
rect 10669 22442 10679 22498
rect 10735 22442 10803 22498
rect 10859 22442 10927 22498
rect 10983 22442 11051 22498
rect 11107 22442 11175 22498
rect 11231 22442 11299 22498
rect 11355 22442 11423 22498
rect 11479 22442 11547 22498
rect 11603 22442 11671 22498
rect 11727 22442 11795 22498
rect 11851 22442 11919 22498
rect 11975 22442 12043 22498
rect 12099 22442 12167 22498
rect 12223 22442 12291 22498
rect 12347 22442 12415 22498
rect 12471 22442 12481 22498
rect 10669 22432 12481 22442
rect 1068 22150 2136 22160
rect 1068 22094 1078 22150
rect 1134 22094 1202 22150
rect 1258 22094 1326 22150
rect 1382 22094 1450 22150
rect 1506 22094 1574 22150
rect 1630 22094 1698 22150
rect 1754 22094 1822 22150
rect 1878 22094 1946 22150
rect 2002 22094 2070 22150
rect 2126 22094 2136 22150
rect 1068 22026 2136 22094
rect 1068 21970 1078 22026
rect 1134 21970 1202 22026
rect 1258 21970 1326 22026
rect 1382 21970 1450 22026
rect 1506 21970 1574 22026
rect 1630 21970 1698 22026
rect 1754 21970 1822 22026
rect 1878 21970 1946 22026
rect 2002 21970 2070 22026
rect 2126 21970 2136 22026
rect 1068 21902 2136 21970
rect 1068 21846 1078 21902
rect 1134 21846 1202 21902
rect 1258 21846 1326 21902
rect 1382 21846 1450 21902
rect 1506 21846 1574 21902
rect 1630 21846 1698 21902
rect 1754 21846 1822 21902
rect 1878 21846 1946 21902
rect 2002 21846 2070 21902
rect 2126 21846 2136 21902
rect 1068 21778 2136 21846
rect 1068 21722 1078 21778
rect 1134 21722 1202 21778
rect 1258 21722 1326 21778
rect 1382 21722 1450 21778
rect 1506 21722 1574 21778
rect 1630 21722 1698 21778
rect 1754 21722 1822 21778
rect 1878 21722 1946 21778
rect 2002 21722 2070 21778
rect 2126 21722 2136 21778
rect 1068 21654 2136 21722
rect 1068 21598 1078 21654
rect 1134 21598 1202 21654
rect 1258 21598 1326 21654
rect 1382 21598 1450 21654
rect 1506 21598 1574 21654
rect 1630 21598 1698 21654
rect 1754 21598 1822 21654
rect 1878 21598 1946 21654
rect 2002 21598 2070 21654
rect 2126 21598 2136 21654
rect 1068 21530 2136 21598
rect 1068 21474 1078 21530
rect 1134 21474 1202 21530
rect 1258 21474 1326 21530
rect 1382 21474 1450 21530
rect 1506 21474 1574 21530
rect 1630 21474 1698 21530
rect 1754 21474 1822 21530
rect 1878 21474 1946 21530
rect 2002 21474 2070 21530
rect 2126 21474 2136 21530
rect 1068 21406 2136 21474
rect 1068 21350 1078 21406
rect 1134 21350 1202 21406
rect 1258 21350 1326 21406
rect 1382 21350 1450 21406
rect 1506 21350 1574 21406
rect 1630 21350 1698 21406
rect 1754 21350 1822 21406
rect 1878 21350 1946 21406
rect 2002 21350 2070 21406
rect 2126 21350 2136 21406
rect 1068 21282 2136 21350
rect 1068 21226 1078 21282
rect 1134 21226 1202 21282
rect 1258 21226 1326 21282
rect 1382 21226 1450 21282
rect 1506 21226 1574 21282
rect 1630 21226 1698 21282
rect 1754 21226 1822 21282
rect 1878 21226 1946 21282
rect 2002 21226 2070 21282
rect 2126 21226 2136 21282
rect 1068 21158 2136 21226
rect 1068 21102 1078 21158
rect 1134 21102 1202 21158
rect 1258 21102 1326 21158
rect 1382 21102 1450 21158
rect 1506 21102 1574 21158
rect 1630 21102 1698 21158
rect 1754 21102 1822 21158
rect 1878 21102 1946 21158
rect 2002 21102 2070 21158
rect 2126 21102 2136 21158
rect 1068 21034 2136 21102
rect 1068 20978 1078 21034
rect 1134 20978 1202 21034
rect 1258 20978 1326 21034
rect 1382 20978 1450 21034
rect 1506 20978 1574 21034
rect 1630 20978 1698 21034
rect 1754 20978 1822 21034
rect 1878 20978 1946 21034
rect 2002 20978 2070 21034
rect 2126 20978 2136 21034
rect 1068 20910 2136 20978
rect 1068 20854 1078 20910
rect 1134 20854 1202 20910
rect 1258 20854 1326 20910
rect 1382 20854 1450 20910
rect 1506 20854 1574 20910
rect 1630 20854 1698 20910
rect 1754 20854 1822 20910
rect 1878 20854 1946 20910
rect 2002 20854 2070 20910
rect 2126 20854 2136 20910
rect 1068 20786 2136 20854
rect 1068 20730 1078 20786
rect 1134 20730 1202 20786
rect 1258 20730 1326 20786
rect 1382 20730 1450 20786
rect 1506 20730 1574 20786
rect 1630 20730 1698 20786
rect 1754 20730 1822 20786
rect 1878 20730 1946 20786
rect 2002 20730 2070 20786
rect 2126 20730 2136 20786
rect 1068 20662 2136 20730
rect 1068 20606 1078 20662
rect 1134 20606 1202 20662
rect 1258 20606 1326 20662
rect 1382 20606 1450 20662
rect 1506 20606 1574 20662
rect 1630 20606 1698 20662
rect 1754 20606 1822 20662
rect 1878 20606 1946 20662
rect 2002 20606 2070 20662
rect 2126 20606 2136 20662
rect 1068 20538 2136 20606
rect 1068 20482 1078 20538
rect 1134 20482 1202 20538
rect 1258 20482 1326 20538
rect 1382 20482 1450 20538
rect 1506 20482 1574 20538
rect 1630 20482 1698 20538
rect 1754 20482 1822 20538
rect 1878 20482 1946 20538
rect 2002 20482 2070 20538
rect 2126 20482 2136 20538
rect 1068 20414 2136 20482
rect 1068 20358 1078 20414
rect 1134 20358 1202 20414
rect 1258 20358 1326 20414
rect 1382 20358 1450 20414
rect 1506 20358 1574 20414
rect 1630 20358 1698 20414
rect 1754 20358 1822 20414
rect 1878 20358 1946 20414
rect 2002 20358 2070 20414
rect 2126 20358 2136 20414
rect 1068 20290 2136 20358
rect 1068 20234 1078 20290
rect 1134 20234 1202 20290
rect 1258 20234 1326 20290
rect 1382 20234 1450 20290
rect 1506 20234 1574 20290
rect 1630 20234 1698 20290
rect 1754 20234 1822 20290
rect 1878 20234 1946 20290
rect 2002 20234 2070 20290
rect 2126 20234 2136 20290
rect 1068 20166 2136 20234
rect 1068 20110 1078 20166
rect 1134 20110 1202 20166
rect 1258 20110 1326 20166
rect 1382 20110 1450 20166
rect 1506 20110 1574 20166
rect 1630 20110 1698 20166
rect 1754 20110 1822 20166
rect 1878 20110 1946 20166
rect 2002 20110 2070 20166
rect 2126 20110 2136 20166
rect 1068 20042 2136 20110
rect 1068 19986 1078 20042
rect 1134 19986 1202 20042
rect 1258 19986 1326 20042
rect 1382 19986 1450 20042
rect 1506 19986 1574 20042
rect 1630 19986 1698 20042
rect 1754 19986 1822 20042
rect 1878 19986 1946 20042
rect 2002 19986 2070 20042
rect 2126 19986 2136 20042
rect 1068 19918 2136 19986
rect 1068 19862 1078 19918
rect 1134 19862 1202 19918
rect 1258 19862 1326 19918
rect 1382 19862 1450 19918
rect 1506 19862 1574 19918
rect 1630 19862 1698 19918
rect 1754 19862 1822 19918
rect 1878 19862 1946 19918
rect 2002 19862 2070 19918
rect 2126 19862 2136 19918
rect 1068 19794 2136 19862
rect 1068 19738 1078 19794
rect 1134 19738 1202 19794
rect 1258 19738 1326 19794
rect 1382 19738 1450 19794
rect 1506 19738 1574 19794
rect 1630 19738 1698 19794
rect 1754 19738 1822 19794
rect 1878 19738 1946 19794
rect 2002 19738 2070 19794
rect 2126 19738 2136 19794
rect 1068 19670 2136 19738
rect 1068 19614 1078 19670
rect 1134 19614 1202 19670
rect 1258 19614 1326 19670
rect 1382 19614 1450 19670
rect 1506 19614 1574 19670
rect 1630 19614 1698 19670
rect 1754 19614 1822 19670
rect 1878 19614 1946 19670
rect 2002 19614 2070 19670
rect 2126 19614 2136 19670
rect 1068 19546 2136 19614
rect 1068 19490 1078 19546
rect 1134 19490 1202 19546
rect 1258 19490 1326 19546
rect 1382 19490 1450 19546
rect 1506 19490 1574 19546
rect 1630 19490 1698 19546
rect 1754 19490 1822 19546
rect 1878 19490 1946 19546
rect 2002 19490 2070 19546
rect 2126 19490 2136 19546
rect 1068 19422 2136 19490
rect 1068 19366 1078 19422
rect 1134 19366 1202 19422
rect 1258 19366 1326 19422
rect 1382 19366 1450 19422
rect 1506 19366 1574 19422
rect 1630 19366 1698 19422
rect 1754 19366 1822 19422
rect 1878 19366 1946 19422
rect 2002 19366 2070 19422
rect 2126 19366 2136 19422
rect 1068 19298 2136 19366
rect 1068 19242 1078 19298
rect 1134 19242 1202 19298
rect 1258 19242 1326 19298
rect 1382 19242 1450 19298
rect 1506 19242 1574 19298
rect 1630 19242 1698 19298
rect 1754 19242 1822 19298
rect 1878 19242 1946 19298
rect 2002 19242 2070 19298
rect 2126 19242 2136 19298
rect 1068 19232 2136 19242
rect 4425 22150 6237 22160
rect 4425 22094 4435 22150
rect 4491 22094 4559 22150
rect 4615 22094 4683 22150
rect 4739 22094 4807 22150
rect 4863 22094 4931 22150
rect 4987 22094 5055 22150
rect 5111 22094 5179 22150
rect 5235 22094 5303 22150
rect 5359 22094 5427 22150
rect 5483 22094 5551 22150
rect 5607 22094 5675 22150
rect 5731 22094 5799 22150
rect 5855 22094 5923 22150
rect 5979 22094 6047 22150
rect 6103 22094 6171 22150
rect 6227 22094 6237 22150
rect 4425 22026 6237 22094
rect 4425 21970 4435 22026
rect 4491 21970 4559 22026
rect 4615 21970 4683 22026
rect 4739 21970 4807 22026
rect 4863 21970 4931 22026
rect 4987 21970 5055 22026
rect 5111 21970 5179 22026
rect 5235 21970 5303 22026
rect 5359 21970 5427 22026
rect 5483 21970 5551 22026
rect 5607 21970 5675 22026
rect 5731 21970 5799 22026
rect 5855 21970 5923 22026
rect 5979 21970 6047 22026
rect 6103 21970 6171 22026
rect 6227 21970 6237 22026
rect 4425 21902 6237 21970
rect 4425 21846 4435 21902
rect 4491 21846 4559 21902
rect 4615 21846 4683 21902
rect 4739 21846 4807 21902
rect 4863 21846 4931 21902
rect 4987 21846 5055 21902
rect 5111 21846 5179 21902
rect 5235 21846 5303 21902
rect 5359 21846 5427 21902
rect 5483 21846 5551 21902
rect 5607 21846 5675 21902
rect 5731 21846 5799 21902
rect 5855 21846 5923 21902
rect 5979 21846 6047 21902
rect 6103 21846 6171 21902
rect 6227 21846 6237 21902
rect 4425 21778 6237 21846
rect 4425 21722 4435 21778
rect 4491 21722 4559 21778
rect 4615 21722 4683 21778
rect 4739 21722 4807 21778
rect 4863 21722 4931 21778
rect 4987 21722 5055 21778
rect 5111 21722 5179 21778
rect 5235 21722 5303 21778
rect 5359 21722 5427 21778
rect 5483 21722 5551 21778
rect 5607 21722 5675 21778
rect 5731 21722 5799 21778
rect 5855 21722 5923 21778
rect 5979 21722 6047 21778
rect 6103 21722 6171 21778
rect 6227 21722 6237 21778
rect 4425 21654 6237 21722
rect 4425 21598 4435 21654
rect 4491 21598 4559 21654
rect 4615 21598 4683 21654
rect 4739 21598 4807 21654
rect 4863 21598 4931 21654
rect 4987 21598 5055 21654
rect 5111 21598 5179 21654
rect 5235 21598 5303 21654
rect 5359 21598 5427 21654
rect 5483 21598 5551 21654
rect 5607 21598 5675 21654
rect 5731 21598 5799 21654
rect 5855 21598 5923 21654
rect 5979 21598 6047 21654
rect 6103 21598 6171 21654
rect 6227 21598 6237 21654
rect 4425 21530 6237 21598
rect 4425 21474 4435 21530
rect 4491 21474 4559 21530
rect 4615 21474 4683 21530
rect 4739 21474 4807 21530
rect 4863 21474 4931 21530
rect 4987 21474 5055 21530
rect 5111 21474 5179 21530
rect 5235 21474 5303 21530
rect 5359 21474 5427 21530
rect 5483 21474 5551 21530
rect 5607 21474 5675 21530
rect 5731 21474 5799 21530
rect 5855 21474 5923 21530
rect 5979 21474 6047 21530
rect 6103 21474 6171 21530
rect 6227 21474 6237 21530
rect 4425 21406 6237 21474
rect 4425 21350 4435 21406
rect 4491 21350 4559 21406
rect 4615 21350 4683 21406
rect 4739 21350 4807 21406
rect 4863 21350 4931 21406
rect 4987 21350 5055 21406
rect 5111 21350 5179 21406
rect 5235 21350 5303 21406
rect 5359 21350 5427 21406
rect 5483 21350 5551 21406
rect 5607 21350 5675 21406
rect 5731 21350 5799 21406
rect 5855 21350 5923 21406
rect 5979 21350 6047 21406
rect 6103 21350 6171 21406
rect 6227 21350 6237 21406
rect 4425 21282 6237 21350
rect 4425 21226 4435 21282
rect 4491 21226 4559 21282
rect 4615 21226 4683 21282
rect 4739 21226 4807 21282
rect 4863 21226 4931 21282
rect 4987 21226 5055 21282
rect 5111 21226 5179 21282
rect 5235 21226 5303 21282
rect 5359 21226 5427 21282
rect 5483 21226 5551 21282
rect 5607 21226 5675 21282
rect 5731 21226 5799 21282
rect 5855 21226 5923 21282
rect 5979 21226 6047 21282
rect 6103 21226 6171 21282
rect 6227 21226 6237 21282
rect 4425 21158 6237 21226
rect 4425 21102 4435 21158
rect 4491 21102 4559 21158
rect 4615 21102 4683 21158
rect 4739 21102 4807 21158
rect 4863 21102 4931 21158
rect 4987 21102 5055 21158
rect 5111 21102 5179 21158
rect 5235 21102 5303 21158
rect 5359 21102 5427 21158
rect 5483 21102 5551 21158
rect 5607 21102 5675 21158
rect 5731 21102 5799 21158
rect 5855 21102 5923 21158
rect 5979 21102 6047 21158
rect 6103 21102 6171 21158
rect 6227 21102 6237 21158
rect 4425 21034 6237 21102
rect 4425 20978 4435 21034
rect 4491 20978 4559 21034
rect 4615 20978 4683 21034
rect 4739 20978 4807 21034
rect 4863 20978 4931 21034
rect 4987 20978 5055 21034
rect 5111 20978 5179 21034
rect 5235 20978 5303 21034
rect 5359 20978 5427 21034
rect 5483 20978 5551 21034
rect 5607 20978 5675 21034
rect 5731 20978 5799 21034
rect 5855 20978 5923 21034
rect 5979 20978 6047 21034
rect 6103 20978 6171 21034
rect 6227 20978 6237 21034
rect 4425 20910 6237 20978
rect 4425 20854 4435 20910
rect 4491 20854 4559 20910
rect 4615 20854 4683 20910
rect 4739 20854 4807 20910
rect 4863 20854 4931 20910
rect 4987 20854 5055 20910
rect 5111 20854 5179 20910
rect 5235 20854 5303 20910
rect 5359 20854 5427 20910
rect 5483 20854 5551 20910
rect 5607 20854 5675 20910
rect 5731 20854 5799 20910
rect 5855 20854 5923 20910
rect 5979 20854 6047 20910
rect 6103 20854 6171 20910
rect 6227 20854 6237 20910
rect 4425 20786 6237 20854
rect 4425 20730 4435 20786
rect 4491 20730 4559 20786
rect 4615 20730 4683 20786
rect 4739 20730 4807 20786
rect 4863 20730 4931 20786
rect 4987 20730 5055 20786
rect 5111 20730 5179 20786
rect 5235 20730 5303 20786
rect 5359 20730 5427 20786
rect 5483 20730 5551 20786
rect 5607 20730 5675 20786
rect 5731 20730 5799 20786
rect 5855 20730 5923 20786
rect 5979 20730 6047 20786
rect 6103 20730 6171 20786
rect 6227 20730 6237 20786
rect 4425 20662 6237 20730
rect 4425 20606 4435 20662
rect 4491 20606 4559 20662
rect 4615 20606 4683 20662
rect 4739 20606 4807 20662
rect 4863 20606 4931 20662
rect 4987 20606 5055 20662
rect 5111 20606 5179 20662
rect 5235 20606 5303 20662
rect 5359 20606 5427 20662
rect 5483 20606 5551 20662
rect 5607 20606 5675 20662
rect 5731 20606 5799 20662
rect 5855 20606 5923 20662
rect 5979 20606 6047 20662
rect 6103 20606 6171 20662
rect 6227 20606 6237 20662
rect 4425 20538 6237 20606
rect 4425 20482 4435 20538
rect 4491 20482 4559 20538
rect 4615 20482 4683 20538
rect 4739 20482 4807 20538
rect 4863 20482 4931 20538
rect 4987 20482 5055 20538
rect 5111 20482 5179 20538
rect 5235 20482 5303 20538
rect 5359 20482 5427 20538
rect 5483 20482 5551 20538
rect 5607 20482 5675 20538
rect 5731 20482 5799 20538
rect 5855 20482 5923 20538
rect 5979 20482 6047 20538
rect 6103 20482 6171 20538
rect 6227 20482 6237 20538
rect 4425 20414 6237 20482
rect 4425 20358 4435 20414
rect 4491 20358 4559 20414
rect 4615 20358 4683 20414
rect 4739 20358 4807 20414
rect 4863 20358 4931 20414
rect 4987 20358 5055 20414
rect 5111 20358 5179 20414
rect 5235 20358 5303 20414
rect 5359 20358 5427 20414
rect 5483 20358 5551 20414
rect 5607 20358 5675 20414
rect 5731 20358 5799 20414
rect 5855 20358 5923 20414
rect 5979 20358 6047 20414
rect 6103 20358 6171 20414
rect 6227 20358 6237 20414
rect 4425 20290 6237 20358
rect 4425 20234 4435 20290
rect 4491 20234 4559 20290
rect 4615 20234 4683 20290
rect 4739 20234 4807 20290
rect 4863 20234 4931 20290
rect 4987 20234 5055 20290
rect 5111 20234 5179 20290
rect 5235 20234 5303 20290
rect 5359 20234 5427 20290
rect 5483 20234 5551 20290
rect 5607 20234 5675 20290
rect 5731 20234 5799 20290
rect 5855 20234 5923 20290
rect 5979 20234 6047 20290
rect 6103 20234 6171 20290
rect 6227 20234 6237 20290
rect 4425 20166 6237 20234
rect 4425 20110 4435 20166
rect 4491 20110 4559 20166
rect 4615 20110 4683 20166
rect 4739 20110 4807 20166
rect 4863 20110 4931 20166
rect 4987 20110 5055 20166
rect 5111 20110 5179 20166
rect 5235 20110 5303 20166
rect 5359 20110 5427 20166
rect 5483 20110 5551 20166
rect 5607 20110 5675 20166
rect 5731 20110 5799 20166
rect 5855 20110 5923 20166
rect 5979 20110 6047 20166
rect 6103 20110 6171 20166
rect 6227 20110 6237 20166
rect 4425 20042 6237 20110
rect 4425 19986 4435 20042
rect 4491 19986 4559 20042
rect 4615 19986 4683 20042
rect 4739 19986 4807 20042
rect 4863 19986 4931 20042
rect 4987 19986 5055 20042
rect 5111 19986 5179 20042
rect 5235 19986 5303 20042
rect 5359 19986 5427 20042
rect 5483 19986 5551 20042
rect 5607 19986 5675 20042
rect 5731 19986 5799 20042
rect 5855 19986 5923 20042
rect 5979 19986 6047 20042
rect 6103 19986 6171 20042
rect 6227 19986 6237 20042
rect 4425 19918 6237 19986
rect 4425 19862 4435 19918
rect 4491 19862 4559 19918
rect 4615 19862 4683 19918
rect 4739 19862 4807 19918
rect 4863 19862 4931 19918
rect 4987 19862 5055 19918
rect 5111 19862 5179 19918
rect 5235 19862 5303 19918
rect 5359 19862 5427 19918
rect 5483 19862 5551 19918
rect 5607 19862 5675 19918
rect 5731 19862 5799 19918
rect 5855 19862 5923 19918
rect 5979 19862 6047 19918
rect 6103 19862 6171 19918
rect 6227 19862 6237 19918
rect 4425 19794 6237 19862
rect 4425 19738 4435 19794
rect 4491 19738 4559 19794
rect 4615 19738 4683 19794
rect 4739 19738 4807 19794
rect 4863 19738 4931 19794
rect 4987 19738 5055 19794
rect 5111 19738 5179 19794
rect 5235 19738 5303 19794
rect 5359 19738 5427 19794
rect 5483 19738 5551 19794
rect 5607 19738 5675 19794
rect 5731 19738 5799 19794
rect 5855 19738 5923 19794
rect 5979 19738 6047 19794
rect 6103 19738 6171 19794
rect 6227 19738 6237 19794
rect 4425 19670 6237 19738
rect 4425 19614 4435 19670
rect 4491 19614 4559 19670
rect 4615 19614 4683 19670
rect 4739 19614 4807 19670
rect 4863 19614 4931 19670
rect 4987 19614 5055 19670
rect 5111 19614 5179 19670
rect 5235 19614 5303 19670
rect 5359 19614 5427 19670
rect 5483 19614 5551 19670
rect 5607 19614 5675 19670
rect 5731 19614 5799 19670
rect 5855 19614 5923 19670
rect 5979 19614 6047 19670
rect 6103 19614 6171 19670
rect 6227 19614 6237 19670
rect 4425 19546 6237 19614
rect 4425 19490 4435 19546
rect 4491 19490 4559 19546
rect 4615 19490 4683 19546
rect 4739 19490 4807 19546
rect 4863 19490 4931 19546
rect 4987 19490 5055 19546
rect 5111 19490 5179 19546
rect 5235 19490 5303 19546
rect 5359 19490 5427 19546
rect 5483 19490 5551 19546
rect 5607 19490 5675 19546
rect 5731 19490 5799 19546
rect 5855 19490 5923 19546
rect 5979 19490 6047 19546
rect 6103 19490 6171 19546
rect 6227 19490 6237 19546
rect 4425 19422 6237 19490
rect 4425 19366 4435 19422
rect 4491 19366 4559 19422
rect 4615 19366 4683 19422
rect 4739 19366 4807 19422
rect 4863 19366 4931 19422
rect 4987 19366 5055 19422
rect 5111 19366 5179 19422
rect 5235 19366 5303 19422
rect 5359 19366 5427 19422
rect 5483 19366 5551 19422
rect 5607 19366 5675 19422
rect 5731 19366 5799 19422
rect 5855 19366 5923 19422
rect 5979 19366 6047 19422
rect 6103 19366 6171 19422
rect 6227 19366 6237 19422
rect 4425 19298 6237 19366
rect 4425 19242 4435 19298
rect 4491 19242 4559 19298
rect 4615 19242 4683 19298
rect 4739 19242 4807 19298
rect 4863 19242 4931 19298
rect 4987 19242 5055 19298
rect 5111 19242 5179 19298
rect 5235 19242 5303 19298
rect 5359 19242 5427 19298
rect 5483 19242 5551 19298
rect 5607 19242 5675 19298
rect 5731 19242 5799 19298
rect 5855 19242 5923 19298
rect 5979 19242 6047 19298
rect 6103 19242 6171 19298
rect 6227 19242 6237 19298
rect 4425 19232 6237 19242
rect 7552 22150 8620 22160
rect 7552 22094 7562 22150
rect 7618 22094 7686 22150
rect 7742 22094 7810 22150
rect 7866 22094 7934 22150
rect 7990 22094 8058 22150
rect 8114 22094 8182 22150
rect 8238 22094 8306 22150
rect 8362 22094 8430 22150
rect 8486 22094 8554 22150
rect 8610 22094 8620 22150
rect 7552 22026 8620 22094
rect 7552 21970 7562 22026
rect 7618 21970 7686 22026
rect 7742 21970 7810 22026
rect 7866 21970 7934 22026
rect 7990 21970 8058 22026
rect 8114 21970 8182 22026
rect 8238 21970 8306 22026
rect 8362 21970 8430 22026
rect 8486 21970 8554 22026
rect 8610 21970 8620 22026
rect 7552 21902 8620 21970
rect 7552 21846 7562 21902
rect 7618 21846 7686 21902
rect 7742 21846 7810 21902
rect 7866 21846 7934 21902
rect 7990 21846 8058 21902
rect 8114 21846 8182 21902
rect 8238 21846 8306 21902
rect 8362 21846 8430 21902
rect 8486 21846 8554 21902
rect 8610 21846 8620 21902
rect 7552 21778 8620 21846
rect 7552 21722 7562 21778
rect 7618 21722 7686 21778
rect 7742 21722 7810 21778
rect 7866 21722 7934 21778
rect 7990 21722 8058 21778
rect 8114 21722 8182 21778
rect 8238 21722 8306 21778
rect 8362 21722 8430 21778
rect 8486 21722 8554 21778
rect 8610 21722 8620 21778
rect 7552 21654 8620 21722
rect 7552 21598 7562 21654
rect 7618 21598 7686 21654
rect 7742 21598 7810 21654
rect 7866 21598 7934 21654
rect 7990 21598 8058 21654
rect 8114 21598 8182 21654
rect 8238 21598 8306 21654
rect 8362 21598 8430 21654
rect 8486 21598 8554 21654
rect 8610 21598 8620 21654
rect 7552 21530 8620 21598
rect 7552 21474 7562 21530
rect 7618 21474 7686 21530
rect 7742 21474 7810 21530
rect 7866 21474 7934 21530
rect 7990 21474 8058 21530
rect 8114 21474 8182 21530
rect 8238 21474 8306 21530
rect 8362 21474 8430 21530
rect 8486 21474 8554 21530
rect 8610 21474 8620 21530
rect 7552 21406 8620 21474
rect 7552 21350 7562 21406
rect 7618 21350 7686 21406
rect 7742 21350 7810 21406
rect 7866 21350 7934 21406
rect 7990 21350 8058 21406
rect 8114 21350 8182 21406
rect 8238 21350 8306 21406
rect 8362 21350 8430 21406
rect 8486 21350 8554 21406
rect 8610 21350 8620 21406
rect 7552 21282 8620 21350
rect 7552 21226 7562 21282
rect 7618 21226 7686 21282
rect 7742 21226 7810 21282
rect 7866 21226 7934 21282
rect 7990 21226 8058 21282
rect 8114 21226 8182 21282
rect 8238 21226 8306 21282
rect 8362 21226 8430 21282
rect 8486 21226 8554 21282
rect 8610 21226 8620 21282
rect 7552 21158 8620 21226
rect 7552 21102 7562 21158
rect 7618 21102 7686 21158
rect 7742 21102 7810 21158
rect 7866 21102 7934 21158
rect 7990 21102 8058 21158
rect 8114 21102 8182 21158
rect 8238 21102 8306 21158
rect 8362 21102 8430 21158
rect 8486 21102 8554 21158
rect 8610 21102 8620 21158
rect 7552 21034 8620 21102
rect 7552 20978 7562 21034
rect 7618 20978 7686 21034
rect 7742 20978 7810 21034
rect 7866 20978 7934 21034
rect 7990 20978 8058 21034
rect 8114 20978 8182 21034
rect 8238 20978 8306 21034
rect 8362 20978 8430 21034
rect 8486 20978 8554 21034
rect 8610 20978 8620 21034
rect 7552 20910 8620 20978
rect 7552 20854 7562 20910
rect 7618 20854 7686 20910
rect 7742 20854 7810 20910
rect 7866 20854 7934 20910
rect 7990 20854 8058 20910
rect 8114 20854 8182 20910
rect 8238 20854 8306 20910
rect 8362 20854 8430 20910
rect 8486 20854 8554 20910
rect 8610 20854 8620 20910
rect 7552 20786 8620 20854
rect 7552 20730 7562 20786
rect 7618 20730 7686 20786
rect 7742 20730 7810 20786
rect 7866 20730 7934 20786
rect 7990 20730 8058 20786
rect 8114 20730 8182 20786
rect 8238 20730 8306 20786
rect 8362 20730 8430 20786
rect 8486 20730 8554 20786
rect 8610 20730 8620 20786
rect 7552 20662 8620 20730
rect 7552 20606 7562 20662
rect 7618 20606 7686 20662
rect 7742 20606 7810 20662
rect 7866 20606 7934 20662
rect 7990 20606 8058 20662
rect 8114 20606 8182 20662
rect 8238 20606 8306 20662
rect 8362 20606 8430 20662
rect 8486 20606 8554 20662
rect 8610 20606 8620 20662
rect 7552 20538 8620 20606
rect 7552 20482 7562 20538
rect 7618 20482 7686 20538
rect 7742 20482 7810 20538
rect 7866 20482 7934 20538
rect 7990 20482 8058 20538
rect 8114 20482 8182 20538
rect 8238 20482 8306 20538
rect 8362 20482 8430 20538
rect 8486 20482 8554 20538
rect 8610 20482 8620 20538
rect 7552 20414 8620 20482
rect 7552 20358 7562 20414
rect 7618 20358 7686 20414
rect 7742 20358 7810 20414
rect 7866 20358 7934 20414
rect 7990 20358 8058 20414
rect 8114 20358 8182 20414
rect 8238 20358 8306 20414
rect 8362 20358 8430 20414
rect 8486 20358 8554 20414
rect 8610 20358 8620 20414
rect 7552 20290 8620 20358
rect 7552 20234 7562 20290
rect 7618 20234 7686 20290
rect 7742 20234 7810 20290
rect 7866 20234 7934 20290
rect 7990 20234 8058 20290
rect 8114 20234 8182 20290
rect 8238 20234 8306 20290
rect 8362 20234 8430 20290
rect 8486 20234 8554 20290
rect 8610 20234 8620 20290
rect 7552 20166 8620 20234
rect 7552 20110 7562 20166
rect 7618 20110 7686 20166
rect 7742 20110 7810 20166
rect 7866 20110 7934 20166
rect 7990 20110 8058 20166
rect 8114 20110 8182 20166
rect 8238 20110 8306 20166
rect 8362 20110 8430 20166
rect 8486 20110 8554 20166
rect 8610 20110 8620 20166
rect 7552 20042 8620 20110
rect 7552 19986 7562 20042
rect 7618 19986 7686 20042
rect 7742 19986 7810 20042
rect 7866 19986 7934 20042
rect 7990 19986 8058 20042
rect 8114 19986 8182 20042
rect 8238 19986 8306 20042
rect 8362 19986 8430 20042
rect 8486 19986 8554 20042
rect 8610 19986 8620 20042
rect 7552 19918 8620 19986
rect 7552 19862 7562 19918
rect 7618 19862 7686 19918
rect 7742 19862 7810 19918
rect 7866 19862 7934 19918
rect 7990 19862 8058 19918
rect 8114 19862 8182 19918
rect 8238 19862 8306 19918
rect 8362 19862 8430 19918
rect 8486 19862 8554 19918
rect 8610 19862 8620 19918
rect 7552 19794 8620 19862
rect 7552 19738 7562 19794
rect 7618 19738 7686 19794
rect 7742 19738 7810 19794
rect 7866 19738 7934 19794
rect 7990 19738 8058 19794
rect 8114 19738 8182 19794
rect 8238 19738 8306 19794
rect 8362 19738 8430 19794
rect 8486 19738 8554 19794
rect 8610 19738 8620 19794
rect 7552 19670 8620 19738
rect 7552 19614 7562 19670
rect 7618 19614 7686 19670
rect 7742 19614 7810 19670
rect 7866 19614 7934 19670
rect 7990 19614 8058 19670
rect 8114 19614 8182 19670
rect 8238 19614 8306 19670
rect 8362 19614 8430 19670
rect 8486 19614 8554 19670
rect 8610 19614 8620 19670
rect 7552 19546 8620 19614
rect 7552 19490 7562 19546
rect 7618 19490 7686 19546
rect 7742 19490 7810 19546
rect 7866 19490 7934 19546
rect 7990 19490 8058 19546
rect 8114 19490 8182 19546
rect 8238 19490 8306 19546
rect 8362 19490 8430 19546
rect 8486 19490 8554 19546
rect 8610 19490 8620 19546
rect 7552 19422 8620 19490
rect 7552 19366 7562 19422
rect 7618 19366 7686 19422
rect 7742 19366 7810 19422
rect 7866 19366 7934 19422
rect 7990 19366 8058 19422
rect 8114 19366 8182 19422
rect 8238 19366 8306 19422
rect 8362 19366 8430 19422
rect 8486 19366 8554 19422
rect 8610 19366 8620 19422
rect 7552 19298 8620 19366
rect 7552 19242 7562 19298
rect 7618 19242 7686 19298
rect 7742 19242 7810 19298
rect 7866 19242 7934 19298
rect 7990 19242 8058 19298
rect 8114 19242 8182 19298
rect 8238 19242 8306 19298
rect 8362 19242 8430 19298
rect 8486 19242 8554 19298
rect 8610 19242 8620 19298
rect 7552 19232 8620 19242
rect 10669 22150 12481 22160
rect 10669 22094 10679 22150
rect 10735 22094 10803 22150
rect 10859 22094 10927 22150
rect 10983 22094 11051 22150
rect 11107 22094 11175 22150
rect 11231 22094 11299 22150
rect 11355 22094 11423 22150
rect 11479 22094 11547 22150
rect 11603 22094 11671 22150
rect 11727 22094 11795 22150
rect 11851 22094 11919 22150
rect 11975 22094 12043 22150
rect 12099 22094 12167 22150
rect 12223 22094 12291 22150
rect 12347 22094 12415 22150
rect 12471 22094 12481 22150
rect 10669 22026 12481 22094
rect 10669 21970 10679 22026
rect 10735 21970 10803 22026
rect 10859 21970 10927 22026
rect 10983 21970 11051 22026
rect 11107 21970 11175 22026
rect 11231 21970 11299 22026
rect 11355 21970 11423 22026
rect 11479 21970 11547 22026
rect 11603 21970 11671 22026
rect 11727 21970 11795 22026
rect 11851 21970 11919 22026
rect 11975 21970 12043 22026
rect 12099 21970 12167 22026
rect 12223 21970 12291 22026
rect 12347 21970 12415 22026
rect 12471 21970 12481 22026
rect 10669 21902 12481 21970
rect 10669 21846 10679 21902
rect 10735 21846 10803 21902
rect 10859 21846 10927 21902
rect 10983 21846 11051 21902
rect 11107 21846 11175 21902
rect 11231 21846 11299 21902
rect 11355 21846 11423 21902
rect 11479 21846 11547 21902
rect 11603 21846 11671 21902
rect 11727 21846 11795 21902
rect 11851 21846 11919 21902
rect 11975 21846 12043 21902
rect 12099 21846 12167 21902
rect 12223 21846 12291 21902
rect 12347 21846 12415 21902
rect 12471 21846 12481 21902
rect 10669 21778 12481 21846
rect 10669 21722 10679 21778
rect 10735 21722 10803 21778
rect 10859 21722 10927 21778
rect 10983 21722 11051 21778
rect 11107 21722 11175 21778
rect 11231 21722 11299 21778
rect 11355 21722 11423 21778
rect 11479 21722 11547 21778
rect 11603 21722 11671 21778
rect 11727 21722 11795 21778
rect 11851 21722 11919 21778
rect 11975 21722 12043 21778
rect 12099 21722 12167 21778
rect 12223 21722 12291 21778
rect 12347 21722 12415 21778
rect 12471 21722 12481 21778
rect 10669 21654 12481 21722
rect 10669 21598 10679 21654
rect 10735 21598 10803 21654
rect 10859 21598 10927 21654
rect 10983 21598 11051 21654
rect 11107 21598 11175 21654
rect 11231 21598 11299 21654
rect 11355 21598 11423 21654
rect 11479 21598 11547 21654
rect 11603 21598 11671 21654
rect 11727 21598 11795 21654
rect 11851 21598 11919 21654
rect 11975 21598 12043 21654
rect 12099 21598 12167 21654
rect 12223 21598 12291 21654
rect 12347 21598 12415 21654
rect 12471 21598 12481 21654
rect 10669 21530 12481 21598
rect 10669 21474 10679 21530
rect 10735 21474 10803 21530
rect 10859 21474 10927 21530
rect 10983 21474 11051 21530
rect 11107 21474 11175 21530
rect 11231 21474 11299 21530
rect 11355 21474 11423 21530
rect 11479 21474 11547 21530
rect 11603 21474 11671 21530
rect 11727 21474 11795 21530
rect 11851 21474 11919 21530
rect 11975 21474 12043 21530
rect 12099 21474 12167 21530
rect 12223 21474 12291 21530
rect 12347 21474 12415 21530
rect 12471 21474 12481 21530
rect 10669 21406 12481 21474
rect 10669 21350 10679 21406
rect 10735 21350 10803 21406
rect 10859 21350 10927 21406
rect 10983 21350 11051 21406
rect 11107 21350 11175 21406
rect 11231 21350 11299 21406
rect 11355 21350 11423 21406
rect 11479 21350 11547 21406
rect 11603 21350 11671 21406
rect 11727 21350 11795 21406
rect 11851 21350 11919 21406
rect 11975 21350 12043 21406
rect 12099 21350 12167 21406
rect 12223 21350 12291 21406
rect 12347 21350 12415 21406
rect 12471 21350 12481 21406
rect 10669 21282 12481 21350
rect 10669 21226 10679 21282
rect 10735 21226 10803 21282
rect 10859 21226 10927 21282
rect 10983 21226 11051 21282
rect 11107 21226 11175 21282
rect 11231 21226 11299 21282
rect 11355 21226 11423 21282
rect 11479 21226 11547 21282
rect 11603 21226 11671 21282
rect 11727 21226 11795 21282
rect 11851 21226 11919 21282
rect 11975 21226 12043 21282
rect 12099 21226 12167 21282
rect 12223 21226 12291 21282
rect 12347 21226 12415 21282
rect 12471 21226 12481 21282
rect 10669 21158 12481 21226
rect 10669 21102 10679 21158
rect 10735 21102 10803 21158
rect 10859 21102 10927 21158
rect 10983 21102 11051 21158
rect 11107 21102 11175 21158
rect 11231 21102 11299 21158
rect 11355 21102 11423 21158
rect 11479 21102 11547 21158
rect 11603 21102 11671 21158
rect 11727 21102 11795 21158
rect 11851 21102 11919 21158
rect 11975 21102 12043 21158
rect 12099 21102 12167 21158
rect 12223 21102 12291 21158
rect 12347 21102 12415 21158
rect 12471 21102 12481 21158
rect 10669 21034 12481 21102
rect 10669 20978 10679 21034
rect 10735 20978 10803 21034
rect 10859 20978 10927 21034
rect 10983 20978 11051 21034
rect 11107 20978 11175 21034
rect 11231 20978 11299 21034
rect 11355 20978 11423 21034
rect 11479 20978 11547 21034
rect 11603 20978 11671 21034
rect 11727 20978 11795 21034
rect 11851 20978 11919 21034
rect 11975 20978 12043 21034
rect 12099 20978 12167 21034
rect 12223 20978 12291 21034
rect 12347 20978 12415 21034
rect 12471 20978 12481 21034
rect 10669 20910 12481 20978
rect 10669 20854 10679 20910
rect 10735 20854 10803 20910
rect 10859 20854 10927 20910
rect 10983 20854 11051 20910
rect 11107 20854 11175 20910
rect 11231 20854 11299 20910
rect 11355 20854 11423 20910
rect 11479 20854 11547 20910
rect 11603 20854 11671 20910
rect 11727 20854 11795 20910
rect 11851 20854 11919 20910
rect 11975 20854 12043 20910
rect 12099 20854 12167 20910
rect 12223 20854 12291 20910
rect 12347 20854 12415 20910
rect 12471 20854 12481 20910
rect 10669 20786 12481 20854
rect 10669 20730 10679 20786
rect 10735 20730 10803 20786
rect 10859 20730 10927 20786
rect 10983 20730 11051 20786
rect 11107 20730 11175 20786
rect 11231 20730 11299 20786
rect 11355 20730 11423 20786
rect 11479 20730 11547 20786
rect 11603 20730 11671 20786
rect 11727 20730 11795 20786
rect 11851 20730 11919 20786
rect 11975 20730 12043 20786
rect 12099 20730 12167 20786
rect 12223 20730 12291 20786
rect 12347 20730 12415 20786
rect 12471 20730 12481 20786
rect 10669 20662 12481 20730
rect 10669 20606 10679 20662
rect 10735 20606 10803 20662
rect 10859 20606 10927 20662
rect 10983 20606 11051 20662
rect 11107 20606 11175 20662
rect 11231 20606 11299 20662
rect 11355 20606 11423 20662
rect 11479 20606 11547 20662
rect 11603 20606 11671 20662
rect 11727 20606 11795 20662
rect 11851 20606 11919 20662
rect 11975 20606 12043 20662
rect 12099 20606 12167 20662
rect 12223 20606 12291 20662
rect 12347 20606 12415 20662
rect 12471 20606 12481 20662
rect 10669 20538 12481 20606
rect 10669 20482 10679 20538
rect 10735 20482 10803 20538
rect 10859 20482 10927 20538
rect 10983 20482 11051 20538
rect 11107 20482 11175 20538
rect 11231 20482 11299 20538
rect 11355 20482 11423 20538
rect 11479 20482 11547 20538
rect 11603 20482 11671 20538
rect 11727 20482 11795 20538
rect 11851 20482 11919 20538
rect 11975 20482 12043 20538
rect 12099 20482 12167 20538
rect 12223 20482 12291 20538
rect 12347 20482 12415 20538
rect 12471 20482 12481 20538
rect 10669 20414 12481 20482
rect 10669 20358 10679 20414
rect 10735 20358 10803 20414
rect 10859 20358 10927 20414
rect 10983 20358 11051 20414
rect 11107 20358 11175 20414
rect 11231 20358 11299 20414
rect 11355 20358 11423 20414
rect 11479 20358 11547 20414
rect 11603 20358 11671 20414
rect 11727 20358 11795 20414
rect 11851 20358 11919 20414
rect 11975 20358 12043 20414
rect 12099 20358 12167 20414
rect 12223 20358 12291 20414
rect 12347 20358 12415 20414
rect 12471 20358 12481 20414
rect 10669 20290 12481 20358
rect 10669 20234 10679 20290
rect 10735 20234 10803 20290
rect 10859 20234 10927 20290
rect 10983 20234 11051 20290
rect 11107 20234 11175 20290
rect 11231 20234 11299 20290
rect 11355 20234 11423 20290
rect 11479 20234 11547 20290
rect 11603 20234 11671 20290
rect 11727 20234 11795 20290
rect 11851 20234 11919 20290
rect 11975 20234 12043 20290
rect 12099 20234 12167 20290
rect 12223 20234 12291 20290
rect 12347 20234 12415 20290
rect 12471 20234 12481 20290
rect 10669 20166 12481 20234
rect 10669 20110 10679 20166
rect 10735 20110 10803 20166
rect 10859 20110 10927 20166
rect 10983 20110 11051 20166
rect 11107 20110 11175 20166
rect 11231 20110 11299 20166
rect 11355 20110 11423 20166
rect 11479 20110 11547 20166
rect 11603 20110 11671 20166
rect 11727 20110 11795 20166
rect 11851 20110 11919 20166
rect 11975 20110 12043 20166
rect 12099 20110 12167 20166
rect 12223 20110 12291 20166
rect 12347 20110 12415 20166
rect 12471 20110 12481 20166
rect 10669 20042 12481 20110
rect 10669 19986 10679 20042
rect 10735 19986 10803 20042
rect 10859 19986 10927 20042
rect 10983 19986 11051 20042
rect 11107 19986 11175 20042
rect 11231 19986 11299 20042
rect 11355 19986 11423 20042
rect 11479 19986 11547 20042
rect 11603 19986 11671 20042
rect 11727 19986 11795 20042
rect 11851 19986 11919 20042
rect 11975 19986 12043 20042
rect 12099 19986 12167 20042
rect 12223 19986 12291 20042
rect 12347 19986 12415 20042
rect 12471 19986 12481 20042
rect 10669 19918 12481 19986
rect 10669 19862 10679 19918
rect 10735 19862 10803 19918
rect 10859 19862 10927 19918
rect 10983 19862 11051 19918
rect 11107 19862 11175 19918
rect 11231 19862 11299 19918
rect 11355 19862 11423 19918
rect 11479 19862 11547 19918
rect 11603 19862 11671 19918
rect 11727 19862 11795 19918
rect 11851 19862 11919 19918
rect 11975 19862 12043 19918
rect 12099 19862 12167 19918
rect 12223 19862 12291 19918
rect 12347 19862 12415 19918
rect 12471 19862 12481 19918
rect 10669 19794 12481 19862
rect 10669 19738 10679 19794
rect 10735 19738 10803 19794
rect 10859 19738 10927 19794
rect 10983 19738 11051 19794
rect 11107 19738 11175 19794
rect 11231 19738 11299 19794
rect 11355 19738 11423 19794
rect 11479 19738 11547 19794
rect 11603 19738 11671 19794
rect 11727 19738 11795 19794
rect 11851 19738 11919 19794
rect 11975 19738 12043 19794
rect 12099 19738 12167 19794
rect 12223 19738 12291 19794
rect 12347 19738 12415 19794
rect 12471 19738 12481 19794
rect 10669 19670 12481 19738
rect 10669 19614 10679 19670
rect 10735 19614 10803 19670
rect 10859 19614 10927 19670
rect 10983 19614 11051 19670
rect 11107 19614 11175 19670
rect 11231 19614 11299 19670
rect 11355 19614 11423 19670
rect 11479 19614 11547 19670
rect 11603 19614 11671 19670
rect 11727 19614 11795 19670
rect 11851 19614 11919 19670
rect 11975 19614 12043 19670
rect 12099 19614 12167 19670
rect 12223 19614 12291 19670
rect 12347 19614 12415 19670
rect 12471 19614 12481 19670
rect 10669 19546 12481 19614
rect 10669 19490 10679 19546
rect 10735 19490 10803 19546
rect 10859 19490 10927 19546
rect 10983 19490 11051 19546
rect 11107 19490 11175 19546
rect 11231 19490 11299 19546
rect 11355 19490 11423 19546
rect 11479 19490 11547 19546
rect 11603 19490 11671 19546
rect 11727 19490 11795 19546
rect 11851 19490 11919 19546
rect 11975 19490 12043 19546
rect 12099 19490 12167 19546
rect 12223 19490 12291 19546
rect 12347 19490 12415 19546
rect 12471 19490 12481 19546
rect 10669 19422 12481 19490
rect 10669 19366 10679 19422
rect 10735 19366 10803 19422
rect 10859 19366 10927 19422
rect 10983 19366 11051 19422
rect 11107 19366 11175 19422
rect 11231 19366 11299 19422
rect 11355 19366 11423 19422
rect 11479 19366 11547 19422
rect 11603 19366 11671 19422
rect 11727 19366 11795 19422
rect 11851 19366 11919 19422
rect 11975 19366 12043 19422
rect 12099 19366 12167 19422
rect 12223 19366 12291 19422
rect 12347 19366 12415 19422
rect 12471 19366 12481 19422
rect 10669 19298 12481 19366
rect 10669 19242 10679 19298
rect 10735 19242 10803 19298
rect 10859 19242 10927 19298
rect 10983 19242 11051 19298
rect 11107 19242 11175 19298
rect 11231 19242 11299 19298
rect 11355 19242 11423 19298
rect 11479 19242 11547 19298
rect 11603 19242 11671 19298
rect 11727 19242 11795 19298
rect 11851 19242 11919 19298
rect 11975 19242 12043 19298
rect 12099 19242 12167 19298
rect 12223 19242 12291 19298
rect 12347 19242 12415 19298
rect 12471 19242 12481 19298
rect 10669 19232 12481 19242
rect 1068 18950 2136 18960
rect 1068 18894 1078 18950
rect 1134 18894 1202 18950
rect 1258 18894 1326 18950
rect 1382 18894 1450 18950
rect 1506 18894 1574 18950
rect 1630 18894 1698 18950
rect 1754 18894 1822 18950
rect 1878 18894 1946 18950
rect 2002 18894 2070 18950
rect 2126 18894 2136 18950
rect 1068 18826 2136 18894
rect 1068 18770 1078 18826
rect 1134 18770 1202 18826
rect 1258 18770 1326 18826
rect 1382 18770 1450 18826
rect 1506 18770 1574 18826
rect 1630 18770 1698 18826
rect 1754 18770 1822 18826
rect 1878 18770 1946 18826
rect 2002 18770 2070 18826
rect 2126 18770 2136 18826
rect 1068 18702 2136 18770
rect 1068 18646 1078 18702
rect 1134 18646 1202 18702
rect 1258 18646 1326 18702
rect 1382 18646 1450 18702
rect 1506 18646 1574 18702
rect 1630 18646 1698 18702
rect 1754 18646 1822 18702
rect 1878 18646 1946 18702
rect 2002 18646 2070 18702
rect 2126 18646 2136 18702
rect 1068 18578 2136 18646
rect 1068 18522 1078 18578
rect 1134 18522 1202 18578
rect 1258 18522 1326 18578
rect 1382 18522 1450 18578
rect 1506 18522 1574 18578
rect 1630 18522 1698 18578
rect 1754 18522 1822 18578
rect 1878 18522 1946 18578
rect 2002 18522 2070 18578
rect 2126 18522 2136 18578
rect 1068 18454 2136 18522
rect 1068 18398 1078 18454
rect 1134 18398 1202 18454
rect 1258 18398 1326 18454
rect 1382 18398 1450 18454
rect 1506 18398 1574 18454
rect 1630 18398 1698 18454
rect 1754 18398 1822 18454
rect 1878 18398 1946 18454
rect 2002 18398 2070 18454
rect 2126 18398 2136 18454
rect 1068 18330 2136 18398
rect 1068 18274 1078 18330
rect 1134 18274 1202 18330
rect 1258 18274 1326 18330
rect 1382 18274 1450 18330
rect 1506 18274 1574 18330
rect 1630 18274 1698 18330
rect 1754 18274 1822 18330
rect 1878 18274 1946 18330
rect 2002 18274 2070 18330
rect 2126 18274 2136 18330
rect 1068 18206 2136 18274
rect 1068 18150 1078 18206
rect 1134 18150 1202 18206
rect 1258 18150 1326 18206
rect 1382 18150 1450 18206
rect 1506 18150 1574 18206
rect 1630 18150 1698 18206
rect 1754 18150 1822 18206
rect 1878 18150 1946 18206
rect 2002 18150 2070 18206
rect 2126 18150 2136 18206
rect 1068 18082 2136 18150
rect 1068 18026 1078 18082
rect 1134 18026 1202 18082
rect 1258 18026 1326 18082
rect 1382 18026 1450 18082
rect 1506 18026 1574 18082
rect 1630 18026 1698 18082
rect 1754 18026 1822 18082
rect 1878 18026 1946 18082
rect 2002 18026 2070 18082
rect 2126 18026 2136 18082
rect 1068 17958 2136 18026
rect 1068 17902 1078 17958
rect 1134 17902 1202 17958
rect 1258 17902 1326 17958
rect 1382 17902 1450 17958
rect 1506 17902 1574 17958
rect 1630 17902 1698 17958
rect 1754 17902 1822 17958
rect 1878 17902 1946 17958
rect 2002 17902 2070 17958
rect 2126 17902 2136 17958
rect 1068 17834 2136 17902
rect 1068 17778 1078 17834
rect 1134 17778 1202 17834
rect 1258 17778 1326 17834
rect 1382 17778 1450 17834
rect 1506 17778 1574 17834
rect 1630 17778 1698 17834
rect 1754 17778 1822 17834
rect 1878 17778 1946 17834
rect 2002 17778 2070 17834
rect 2126 17778 2136 17834
rect 1068 17710 2136 17778
rect 1068 17654 1078 17710
rect 1134 17654 1202 17710
rect 1258 17654 1326 17710
rect 1382 17654 1450 17710
rect 1506 17654 1574 17710
rect 1630 17654 1698 17710
rect 1754 17654 1822 17710
rect 1878 17654 1946 17710
rect 2002 17654 2070 17710
rect 2126 17654 2136 17710
rect 1068 17586 2136 17654
rect 1068 17530 1078 17586
rect 1134 17530 1202 17586
rect 1258 17530 1326 17586
rect 1382 17530 1450 17586
rect 1506 17530 1574 17586
rect 1630 17530 1698 17586
rect 1754 17530 1822 17586
rect 1878 17530 1946 17586
rect 2002 17530 2070 17586
rect 2126 17530 2136 17586
rect 1068 17462 2136 17530
rect 1068 17406 1078 17462
rect 1134 17406 1202 17462
rect 1258 17406 1326 17462
rect 1382 17406 1450 17462
rect 1506 17406 1574 17462
rect 1630 17406 1698 17462
rect 1754 17406 1822 17462
rect 1878 17406 1946 17462
rect 2002 17406 2070 17462
rect 2126 17406 2136 17462
rect 1068 17338 2136 17406
rect 1068 17282 1078 17338
rect 1134 17282 1202 17338
rect 1258 17282 1326 17338
rect 1382 17282 1450 17338
rect 1506 17282 1574 17338
rect 1630 17282 1698 17338
rect 1754 17282 1822 17338
rect 1878 17282 1946 17338
rect 2002 17282 2070 17338
rect 2126 17282 2136 17338
rect 1068 17214 2136 17282
rect 1068 17158 1078 17214
rect 1134 17158 1202 17214
rect 1258 17158 1326 17214
rect 1382 17158 1450 17214
rect 1506 17158 1574 17214
rect 1630 17158 1698 17214
rect 1754 17158 1822 17214
rect 1878 17158 1946 17214
rect 2002 17158 2070 17214
rect 2126 17158 2136 17214
rect 1068 17090 2136 17158
rect 1068 17034 1078 17090
rect 1134 17034 1202 17090
rect 1258 17034 1326 17090
rect 1382 17034 1450 17090
rect 1506 17034 1574 17090
rect 1630 17034 1698 17090
rect 1754 17034 1822 17090
rect 1878 17034 1946 17090
rect 2002 17034 2070 17090
rect 2126 17034 2136 17090
rect 1068 16966 2136 17034
rect 1068 16910 1078 16966
rect 1134 16910 1202 16966
rect 1258 16910 1326 16966
rect 1382 16910 1450 16966
rect 1506 16910 1574 16966
rect 1630 16910 1698 16966
rect 1754 16910 1822 16966
rect 1878 16910 1946 16966
rect 2002 16910 2070 16966
rect 2126 16910 2136 16966
rect 1068 16842 2136 16910
rect 1068 16786 1078 16842
rect 1134 16786 1202 16842
rect 1258 16786 1326 16842
rect 1382 16786 1450 16842
rect 1506 16786 1574 16842
rect 1630 16786 1698 16842
rect 1754 16786 1822 16842
rect 1878 16786 1946 16842
rect 2002 16786 2070 16842
rect 2126 16786 2136 16842
rect 1068 16718 2136 16786
rect 1068 16662 1078 16718
rect 1134 16662 1202 16718
rect 1258 16662 1326 16718
rect 1382 16662 1450 16718
rect 1506 16662 1574 16718
rect 1630 16662 1698 16718
rect 1754 16662 1822 16718
rect 1878 16662 1946 16718
rect 2002 16662 2070 16718
rect 2126 16662 2136 16718
rect 1068 16594 2136 16662
rect 1068 16538 1078 16594
rect 1134 16538 1202 16594
rect 1258 16538 1326 16594
rect 1382 16538 1450 16594
rect 1506 16538 1574 16594
rect 1630 16538 1698 16594
rect 1754 16538 1822 16594
rect 1878 16538 1946 16594
rect 2002 16538 2070 16594
rect 2126 16538 2136 16594
rect 1068 16470 2136 16538
rect 1068 16414 1078 16470
rect 1134 16414 1202 16470
rect 1258 16414 1326 16470
rect 1382 16414 1450 16470
rect 1506 16414 1574 16470
rect 1630 16414 1698 16470
rect 1754 16414 1822 16470
rect 1878 16414 1946 16470
rect 2002 16414 2070 16470
rect 2126 16414 2136 16470
rect 1068 16346 2136 16414
rect 1068 16290 1078 16346
rect 1134 16290 1202 16346
rect 1258 16290 1326 16346
rect 1382 16290 1450 16346
rect 1506 16290 1574 16346
rect 1630 16290 1698 16346
rect 1754 16290 1822 16346
rect 1878 16290 1946 16346
rect 2002 16290 2070 16346
rect 2126 16290 2136 16346
rect 1068 16222 2136 16290
rect 1068 16166 1078 16222
rect 1134 16166 1202 16222
rect 1258 16166 1326 16222
rect 1382 16166 1450 16222
rect 1506 16166 1574 16222
rect 1630 16166 1698 16222
rect 1754 16166 1822 16222
rect 1878 16166 1946 16222
rect 2002 16166 2070 16222
rect 2126 16166 2136 16222
rect 1068 16098 2136 16166
rect 1068 16042 1078 16098
rect 1134 16042 1202 16098
rect 1258 16042 1326 16098
rect 1382 16042 1450 16098
rect 1506 16042 1574 16098
rect 1630 16042 1698 16098
rect 1754 16042 1822 16098
rect 1878 16042 1946 16098
rect 2002 16042 2070 16098
rect 2126 16042 2136 16098
rect 1068 16032 2136 16042
rect 4425 18950 6237 18960
rect 4425 18894 4435 18950
rect 4491 18894 4559 18950
rect 4615 18894 4683 18950
rect 4739 18894 4807 18950
rect 4863 18894 4931 18950
rect 4987 18894 5055 18950
rect 5111 18894 5179 18950
rect 5235 18894 5303 18950
rect 5359 18894 5427 18950
rect 5483 18894 5551 18950
rect 5607 18894 5675 18950
rect 5731 18894 5799 18950
rect 5855 18894 5923 18950
rect 5979 18894 6047 18950
rect 6103 18894 6171 18950
rect 6227 18894 6237 18950
rect 4425 18826 6237 18894
rect 4425 18770 4435 18826
rect 4491 18770 4559 18826
rect 4615 18770 4683 18826
rect 4739 18770 4807 18826
rect 4863 18770 4931 18826
rect 4987 18770 5055 18826
rect 5111 18770 5179 18826
rect 5235 18770 5303 18826
rect 5359 18770 5427 18826
rect 5483 18770 5551 18826
rect 5607 18770 5675 18826
rect 5731 18770 5799 18826
rect 5855 18770 5923 18826
rect 5979 18770 6047 18826
rect 6103 18770 6171 18826
rect 6227 18770 6237 18826
rect 4425 18702 6237 18770
rect 4425 18646 4435 18702
rect 4491 18646 4559 18702
rect 4615 18646 4683 18702
rect 4739 18646 4807 18702
rect 4863 18646 4931 18702
rect 4987 18646 5055 18702
rect 5111 18646 5179 18702
rect 5235 18646 5303 18702
rect 5359 18646 5427 18702
rect 5483 18646 5551 18702
rect 5607 18646 5675 18702
rect 5731 18646 5799 18702
rect 5855 18646 5923 18702
rect 5979 18646 6047 18702
rect 6103 18646 6171 18702
rect 6227 18646 6237 18702
rect 4425 18578 6237 18646
rect 4425 18522 4435 18578
rect 4491 18522 4559 18578
rect 4615 18522 4683 18578
rect 4739 18522 4807 18578
rect 4863 18522 4931 18578
rect 4987 18522 5055 18578
rect 5111 18522 5179 18578
rect 5235 18522 5303 18578
rect 5359 18522 5427 18578
rect 5483 18522 5551 18578
rect 5607 18522 5675 18578
rect 5731 18522 5799 18578
rect 5855 18522 5923 18578
rect 5979 18522 6047 18578
rect 6103 18522 6171 18578
rect 6227 18522 6237 18578
rect 4425 18454 6237 18522
rect 4425 18398 4435 18454
rect 4491 18398 4559 18454
rect 4615 18398 4683 18454
rect 4739 18398 4807 18454
rect 4863 18398 4931 18454
rect 4987 18398 5055 18454
rect 5111 18398 5179 18454
rect 5235 18398 5303 18454
rect 5359 18398 5427 18454
rect 5483 18398 5551 18454
rect 5607 18398 5675 18454
rect 5731 18398 5799 18454
rect 5855 18398 5923 18454
rect 5979 18398 6047 18454
rect 6103 18398 6171 18454
rect 6227 18398 6237 18454
rect 4425 18330 6237 18398
rect 4425 18274 4435 18330
rect 4491 18274 4559 18330
rect 4615 18274 4683 18330
rect 4739 18274 4807 18330
rect 4863 18274 4931 18330
rect 4987 18274 5055 18330
rect 5111 18274 5179 18330
rect 5235 18274 5303 18330
rect 5359 18274 5427 18330
rect 5483 18274 5551 18330
rect 5607 18274 5675 18330
rect 5731 18274 5799 18330
rect 5855 18274 5923 18330
rect 5979 18274 6047 18330
rect 6103 18274 6171 18330
rect 6227 18274 6237 18330
rect 4425 18206 6237 18274
rect 4425 18150 4435 18206
rect 4491 18150 4559 18206
rect 4615 18150 4683 18206
rect 4739 18150 4807 18206
rect 4863 18150 4931 18206
rect 4987 18150 5055 18206
rect 5111 18150 5179 18206
rect 5235 18150 5303 18206
rect 5359 18150 5427 18206
rect 5483 18150 5551 18206
rect 5607 18150 5675 18206
rect 5731 18150 5799 18206
rect 5855 18150 5923 18206
rect 5979 18150 6047 18206
rect 6103 18150 6171 18206
rect 6227 18150 6237 18206
rect 4425 18082 6237 18150
rect 4425 18026 4435 18082
rect 4491 18026 4559 18082
rect 4615 18026 4683 18082
rect 4739 18026 4807 18082
rect 4863 18026 4931 18082
rect 4987 18026 5055 18082
rect 5111 18026 5179 18082
rect 5235 18026 5303 18082
rect 5359 18026 5427 18082
rect 5483 18026 5551 18082
rect 5607 18026 5675 18082
rect 5731 18026 5799 18082
rect 5855 18026 5923 18082
rect 5979 18026 6047 18082
rect 6103 18026 6171 18082
rect 6227 18026 6237 18082
rect 4425 17958 6237 18026
rect 4425 17902 4435 17958
rect 4491 17902 4559 17958
rect 4615 17902 4683 17958
rect 4739 17902 4807 17958
rect 4863 17902 4931 17958
rect 4987 17902 5055 17958
rect 5111 17902 5179 17958
rect 5235 17902 5303 17958
rect 5359 17902 5427 17958
rect 5483 17902 5551 17958
rect 5607 17902 5675 17958
rect 5731 17902 5799 17958
rect 5855 17902 5923 17958
rect 5979 17902 6047 17958
rect 6103 17902 6171 17958
rect 6227 17902 6237 17958
rect 4425 17834 6237 17902
rect 4425 17778 4435 17834
rect 4491 17778 4559 17834
rect 4615 17778 4683 17834
rect 4739 17778 4807 17834
rect 4863 17778 4931 17834
rect 4987 17778 5055 17834
rect 5111 17778 5179 17834
rect 5235 17778 5303 17834
rect 5359 17778 5427 17834
rect 5483 17778 5551 17834
rect 5607 17778 5675 17834
rect 5731 17778 5799 17834
rect 5855 17778 5923 17834
rect 5979 17778 6047 17834
rect 6103 17778 6171 17834
rect 6227 17778 6237 17834
rect 4425 17710 6237 17778
rect 4425 17654 4435 17710
rect 4491 17654 4559 17710
rect 4615 17654 4683 17710
rect 4739 17654 4807 17710
rect 4863 17654 4931 17710
rect 4987 17654 5055 17710
rect 5111 17654 5179 17710
rect 5235 17654 5303 17710
rect 5359 17654 5427 17710
rect 5483 17654 5551 17710
rect 5607 17654 5675 17710
rect 5731 17654 5799 17710
rect 5855 17654 5923 17710
rect 5979 17654 6047 17710
rect 6103 17654 6171 17710
rect 6227 17654 6237 17710
rect 4425 17586 6237 17654
rect 4425 17530 4435 17586
rect 4491 17530 4559 17586
rect 4615 17530 4683 17586
rect 4739 17530 4807 17586
rect 4863 17530 4931 17586
rect 4987 17530 5055 17586
rect 5111 17530 5179 17586
rect 5235 17530 5303 17586
rect 5359 17530 5427 17586
rect 5483 17530 5551 17586
rect 5607 17530 5675 17586
rect 5731 17530 5799 17586
rect 5855 17530 5923 17586
rect 5979 17530 6047 17586
rect 6103 17530 6171 17586
rect 6227 17530 6237 17586
rect 4425 17462 6237 17530
rect 4425 17406 4435 17462
rect 4491 17406 4559 17462
rect 4615 17406 4683 17462
rect 4739 17406 4807 17462
rect 4863 17406 4931 17462
rect 4987 17406 5055 17462
rect 5111 17406 5179 17462
rect 5235 17406 5303 17462
rect 5359 17406 5427 17462
rect 5483 17406 5551 17462
rect 5607 17406 5675 17462
rect 5731 17406 5799 17462
rect 5855 17406 5923 17462
rect 5979 17406 6047 17462
rect 6103 17406 6171 17462
rect 6227 17406 6237 17462
rect 4425 17338 6237 17406
rect 4425 17282 4435 17338
rect 4491 17282 4559 17338
rect 4615 17282 4683 17338
rect 4739 17282 4807 17338
rect 4863 17282 4931 17338
rect 4987 17282 5055 17338
rect 5111 17282 5179 17338
rect 5235 17282 5303 17338
rect 5359 17282 5427 17338
rect 5483 17282 5551 17338
rect 5607 17282 5675 17338
rect 5731 17282 5799 17338
rect 5855 17282 5923 17338
rect 5979 17282 6047 17338
rect 6103 17282 6171 17338
rect 6227 17282 6237 17338
rect 4425 17214 6237 17282
rect 4425 17158 4435 17214
rect 4491 17158 4559 17214
rect 4615 17158 4683 17214
rect 4739 17158 4807 17214
rect 4863 17158 4931 17214
rect 4987 17158 5055 17214
rect 5111 17158 5179 17214
rect 5235 17158 5303 17214
rect 5359 17158 5427 17214
rect 5483 17158 5551 17214
rect 5607 17158 5675 17214
rect 5731 17158 5799 17214
rect 5855 17158 5923 17214
rect 5979 17158 6047 17214
rect 6103 17158 6171 17214
rect 6227 17158 6237 17214
rect 4425 17090 6237 17158
rect 4425 17034 4435 17090
rect 4491 17034 4559 17090
rect 4615 17034 4683 17090
rect 4739 17034 4807 17090
rect 4863 17034 4931 17090
rect 4987 17034 5055 17090
rect 5111 17034 5179 17090
rect 5235 17034 5303 17090
rect 5359 17034 5427 17090
rect 5483 17034 5551 17090
rect 5607 17034 5675 17090
rect 5731 17034 5799 17090
rect 5855 17034 5923 17090
rect 5979 17034 6047 17090
rect 6103 17034 6171 17090
rect 6227 17034 6237 17090
rect 4425 16966 6237 17034
rect 4425 16910 4435 16966
rect 4491 16910 4559 16966
rect 4615 16910 4683 16966
rect 4739 16910 4807 16966
rect 4863 16910 4931 16966
rect 4987 16910 5055 16966
rect 5111 16910 5179 16966
rect 5235 16910 5303 16966
rect 5359 16910 5427 16966
rect 5483 16910 5551 16966
rect 5607 16910 5675 16966
rect 5731 16910 5799 16966
rect 5855 16910 5923 16966
rect 5979 16910 6047 16966
rect 6103 16910 6171 16966
rect 6227 16910 6237 16966
rect 4425 16842 6237 16910
rect 4425 16786 4435 16842
rect 4491 16786 4559 16842
rect 4615 16786 4683 16842
rect 4739 16786 4807 16842
rect 4863 16786 4931 16842
rect 4987 16786 5055 16842
rect 5111 16786 5179 16842
rect 5235 16786 5303 16842
rect 5359 16786 5427 16842
rect 5483 16786 5551 16842
rect 5607 16786 5675 16842
rect 5731 16786 5799 16842
rect 5855 16786 5923 16842
rect 5979 16786 6047 16842
rect 6103 16786 6171 16842
rect 6227 16786 6237 16842
rect 4425 16718 6237 16786
rect 4425 16662 4435 16718
rect 4491 16662 4559 16718
rect 4615 16662 4683 16718
rect 4739 16662 4807 16718
rect 4863 16662 4931 16718
rect 4987 16662 5055 16718
rect 5111 16662 5179 16718
rect 5235 16662 5303 16718
rect 5359 16662 5427 16718
rect 5483 16662 5551 16718
rect 5607 16662 5675 16718
rect 5731 16662 5799 16718
rect 5855 16662 5923 16718
rect 5979 16662 6047 16718
rect 6103 16662 6171 16718
rect 6227 16662 6237 16718
rect 4425 16594 6237 16662
rect 4425 16538 4435 16594
rect 4491 16538 4559 16594
rect 4615 16538 4683 16594
rect 4739 16538 4807 16594
rect 4863 16538 4931 16594
rect 4987 16538 5055 16594
rect 5111 16538 5179 16594
rect 5235 16538 5303 16594
rect 5359 16538 5427 16594
rect 5483 16538 5551 16594
rect 5607 16538 5675 16594
rect 5731 16538 5799 16594
rect 5855 16538 5923 16594
rect 5979 16538 6047 16594
rect 6103 16538 6171 16594
rect 6227 16538 6237 16594
rect 4425 16470 6237 16538
rect 4425 16414 4435 16470
rect 4491 16414 4559 16470
rect 4615 16414 4683 16470
rect 4739 16414 4807 16470
rect 4863 16414 4931 16470
rect 4987 16414 5055 16470
rect 5111 16414 5179 16470
rect 5235 16414 5303 16470
rect 5359 16414 5427 16470
rect 5483 16414 5551 16470
rect 5607 16414 5675 16470
rect 5731 16414 5799 16470
rect 5855 16414 5923 16470
rect 5979 16414 6047 16470
rect 6103 16414 6171 16470
rect 6227 16414 6237 16470
rect 4425 16346 6237 16414
rect 4425 16290 4435 16346
rect 4491 16290 4559 16346
rect 4615 16290 4683 16346
rect 4739 16290 4807 16346
rect 4863 16290 4931 16346
rect 4987 16290 5055 16346
rect 5111 16290 5179 16346
rect 5235 16290 5303 16346
rect 5359 16290 5427 16346
rect 5483 16290 5551 16346
rect 5607 16290 5675 16346
rect 5731 16290 5799 16346
rect 5855 16290 5923 16346
rect 5979 16290 6047 16346
rect 6103 16290 6171 16346
rect 6227 16290 6237 16346
rect 4425 16222 6237 16290
rect 4425 16166 4435 16222
rect 4491 16166 4559 16222
rect 4615 16166 4683 16222
rect 4739 16166 4807 16222
rect 4863 16166 4931 16222
rect 4987 16166 5055 16222
rect 5111 16166 5179 16222
rect 5235 16166 5303 16222
rect 5359 16166 5427 16222
rect 5483 16166 5551 16222
rect 5607 16166 5675 16222
rect 5731 16166 5799 16222
rect 5855 16166 5923 16222
rect 5979 16166 6047 16222
rect 6103 16166 6171 16222
rect 6227 16166 6237 16222
rect 4425 16098 6237 16166
rect 4425 16042 4435 16098
rect 4491 16042 4559 16098
rect 4615 16042 4683 16098
rect 4739 16042 4807 16098
rect 4863 16042 4931 16098
rect 4987 16042 5055 16098
rect 5111 16042 5179 16098
rect 5235 16042 5303 16098
rect 5359 16042 5427 16098
rect 5483 16042 5551 16098
rect 5607 16042 5675 16098
rect 5731 16042 5799 16098
rect 5855 16042 5923 16098
rect 5979 16042 6047 16098
rect 6103 16042 6171 16098
rect 6227 16042 6237 16098
rect 4425 16032 6237 16042
rect 7552 18950 8620 18960
rect 7552 18894 7562 18950
rect 7618 18894 7686 18950
rect 7742 18894 7810 18950
rect 7866 18894 7934 18950
rect 7990 18894 8058 18950
rect 8114 18894 8182 18950
rect 8238 18894 8306 18950
rect 8362 18894 8430 18950
rect 8486 18894 8554 18950
rect 8610 18894 8620 18950
rect 7552 18826 8620 18894
rect 7552 18770 7562 18826
rect 7618 18770 7686 18826
rect 7742 18770 7810 18826
rect 7866 18770 7934 18826
rect 7990 18770 8058 18826
rect 8114 18770 8182 18826
rect 8238 18770 8306 18826
rect 8362 18770 8430 18826
rect 8486 18770 8554 18826
rect 8610 18770 8620 18826
rect 7552 18702 8620 18770
rect 7552 18646 7562 18702
rect 7618 18646 7686 18702
rect 7742 18646 7810 18702
rect 7866 18646 7934 18702
rect 7990 18646 8058 18702
rect 8114 18646 8182 18702
rect 8238 18646 8306 18702
rect 8362 18646 8430 18702
rect 8486 18646 8554 18702
rect 8610 18646 8620 18702
rect 7552 18578 8620 18646
rect 7552 18522 7562 18578
rect 7618 18522 7686 18578
rect 7742 18522 7810 18578
rect 7866 18522 7934 18578
rect 7990 18522 8058 18578
rect 8114 18522 8182 18578
rect 8238 18522 8306 18578
rect 8362 18522 8430 18578
rect 8486 18522 8554 18578
rect 8610 18522 8620 18578
rect 7552 18454 8620 18522
rect 7552 18398 7562 18454
rect 7618 18398 7686 18454
rect 7742 18398 7810 18454
rect 7866 18398 7934 18454
rect 7990 18398 8058 18454
rect 8114 18398 8182 18454
rect 8238 18398 8306 18454
rect 8362 18398 8430 18454
rect 8486 18398 8554 18454
rect 8610 18398 8620 18454
rect 7552 18330 8620 18398
rect 7552 18274 7562 18330
rect 7618 18274 7686 18330
rect 7742 18274 7810 18330
rect 7866 18274 7934 18330
rect 7990 18274 8058 18330
rect 8114 18274 8182 18330
rect 8238 18274 8306 18330
rect 8362 18274 8430 18330
rect 8486 18274 8554 18330
rect 8610 18274 8620 18330
rect 7552 18206 8620 18274
rect 7552 18150 7562 18206
rect 7618 18150 7686 18206
rect 7742 18150 7810 18206
rect 7866 18150 7934 18206
rect 7990 18150 8058 18206
rect 8114 18150 8182 18206
rect 8238 18150 8306 18206
rect 8362 18150 8430 18206
rect 8486 18150 8554 18206
rect 8610 18150 8620 18206
rect 7552 18082 8620 18150
rect 7552 18026 7562 18082
rect 7618 18026 7686 18082
rect 7742 18026 7810 18082
rect 7866 18026 7934 18082
rect 7990 18026 8058 18082
rect 8114 18026 8182 18082
rect 8238 18026 8306 18082
rect 8362 18026 8430 18082
rect 8486 18026 8554 18082
rect 8610 18026 8620 18082
rect 7552 17958 8620 18026
rect 7552 17902 7562 17958
rect 7618 17902 7686 17958
rect 7742 17902 7810 17958
rect 7866 17902 7934 17958
rect 7990 17902 8058 17958
rect 8114 17902 8182 17958
rect 8238 17902 8306 17958
rect 8362 17902 8430 17958
rect 8486 17902 8554 17958
rect 8610 17902 8620 17958
rect 7552 17834 8620 17902
rect 7552 17778 7562 17834
rect 7618 17778 7686 17834
rect 7742 17778 7810 17834
rect 7866 17778 7934 17834
rect 7990 17778 8058 17834
rect 8114 17778 8182 17834
rect 8238 17778 8306 17834
rect 8362 17778 8430 17834
rect 8486 17778 8554 17834
rect 8610 17778 8620 17834
rect 7552 17710 8620 17778
rect 7552 17654 7562 17710
rect 7618 17654 7686 17710
rect 7742 17654 7810 17710
rect 7866 17654 7934 17710
rect 7990 17654 8058 17710
rect 8114 17654 8182 17710
rect 8238 17654 8306 17710
rect 8362 17654 8430 17710
rect 8486 17654 8554 17710
rect 8610 17654 8620 17710
rect 7552 17586 8620 17654
rect 7552 17530 7562 17586
rect 7618 17530 7686 17586
rect 7742 17530 7810 17586
rect 7866 17530 7934 17586
rect 7990 17530 8058 17586
rect 8114 17530 8182 17586
rect 8238 17530 8306 17586
rect 8362 17530 8430 17586
rect 8486 17530 8554 17586
rect 8610 17530 8620 17586
rect 7552 17462 8620 17530
rect 7552 17406 7562 17462
rect 7618 17406 7686 17462
rect 7742 17406 7810 17462
rect 7866 17406 7934 17462
rect 7990 17406 8058 17462
rect 8114 17406 8182 17462
rect 8238 17406 8306 17462
rect 8362 17406 8430 17462
rect 8486 17406 8554 17462
rect 8610 17406 8620 17462
rect 7552 17338 8620 17406
rect 7552 17282 7562 17338
rect 7618 17282 7686 17338
rect 7742 17282 7810 17338
rect 7866 17282 7934 17338
rect 7990 17282 8058 17338
rect 8114 17282 8182 17338
rect 8238 17282 8306 17338
rect 8362 17282 8430 17338
rect 8486 17282 8554 17338
rect 8610 17282 8620 17338
rect 7552 17214 8620 17282
rect 7552 17158 7562 17214
rect 7618 17158 7686 17214
rect 7742 17158 7810 17214
rect 7866 17158 7934 17214
rect 7990 17158 8058 17214
rect 8114 17158 8182 17214
rect 8238 17158 8306 17214
rect 8362 17158 8430 17214
rect 8486 17158 8554 17214
rect 8610 17158 8620 17214
rect 7552 17090 8620 17158
rect 7552 17034 7562 17090
rect 7618 17034 7686 17090
rect 7742 17034 7810 17090
rect 7866 17034 7934 17090
rect 7990 17034 8058 17090
rect 8114 17034 8182 17090
rect 8238 17034 8306 17090
rect 8362 17034 8430 17090
rect 8486 17034 8554 17090
rect 8610 17034 8620 17090
rect 7552 16966 8620 17034
rect 7552 16910 7562 16966
rect 7618 16910 7686 16966
rect 7742 16910 7810 16966
rect 7866 16910 7934 16966
rect 7990 16910 8058 16966
rect 8114 16910 8182 16966
rect 8238 16910 8306 16966
rect 8362 16910 8430 16966
rect 8486 16910 8554 16966
rect 8610 16910 8620 16966
rect 7552 16842 8620 16910
rect 7552 16786 7562 16842
rect 7618 16786 7686 16842
rect 7742 16786 7810 16842
rect 7866 16786 7934 16842
rect 7990 16786 8058 16842
rect 8114 16786 8182 16842
rect 8238 16786 8306 16842
rect 8362 16786 8430 16842
rect 8486 16786 8554 16842
rect 8610 16786 8620 16842
rect 7552 16718 8620 16786
rect 7552 16662 7562 16718
rect 7618 16662 7686 16718
rect 7742 16662 7810 16718
rect 7866 16662 7934 16718
rect 7990 16662 8058 16718
rect 8114 16662 8182 16718
rect 8238 16662 8306 16718
rect 8362 16662 8430 16718
rect 8486 16662 8554 16718
rect 8610 16662 8620 16718
rect 7552 16594 8620 16662
rect 7552 16538 7562 16594
rect 7618 16538 7686 16594
rect 7742 16538 7810 16594
rect 7866 16538 7934 16594
rect 7990 16538 8058 16594
rect 8114 16538 8182 16594
rect 8238 16538 8306 16594
rect 8362 16538 8430 16594
rect 8486 16538 8554 16594
rect 8610 16538 8620 16594
rect 7552 16470 8620 16538
rect 7552 16414 7562 16470
rect 7618 16414 7686 16470
rect 7742 16414 7810 16470
rect 7866 16414 7934 16470
rect 7990 16414 8058 16470
rect 8114 16414 8182 16470
rect 8238 16414 8306 16470
rect 8362 16414 8430 16470
rect 8486 16414 8554 16470
rect 8610 16414 8620 16470
rect 7552 16346 8620 16414
rect 7552 16290 7562 16346
rect 7618 16290 7686 16346
rect 7742 16290 7810 16346
rect 7866 16290 7934 16346
rect 7990 16290 8058 16346
rect 8114 16290 8182 16346
rect 8238 16290 8306 16346
rect 8362 16290 8430 16346
rect 8486 16290 8554 16346
rect 8610 16290 8620 16346
rect 7552 16222 8620 16290
rect 7552 16166 7562 16222
rect 7618 16166 7686 16222
rect 7742 16166 7810 16222
rect 7866 16166 7934 16222
rect 7990 16166 8058 16222
rect 8114 16166 8182 16222
rect 8238 16166 8306 16222
rect 8362 16166 8430 16222
rect 8486 16166 8554 16222
rect 8610 16166 8620 16222
rect 7552 16098 8620 16166
rect 7552 16042 7562 16098
rect 7618 16042 7686 16098
rect 7742 16042 7810 16098
rect 7866 16042 7934 16098
rect 7990 16042 8058 16098
rect 8114 16042 8182 16098
rect 8238 16042 8306 16098
rect 8362 16042 8430 16098
rect 8486 16042 8554 16098
rect 8610 16042 8620 16098
rect 7552 16032 8620 16042
rect 10669 18950 12481 18960
rect 10669 18894 10679 18950
rect 10735 18894 10803 18950
rect 10859 18894 10927 18950
rect 10983 18894 11051 18950
rect 11107 18894 11175 18950
rect 11231 18894 11299 18950
rect 11355 18894 11423 18950
rect 11479 18894 11547 18950
rect 11603 18894 11671 18950
rect 11727 18894 11795 18950
rect 11851 18894 11919 18950
rect 11975 18894 12043 18950
rect 12099 18894 12167 18950
rect 12223 18894 12291 18950
rect 12347 18894 12415 18950
rect 12471 18894 12481 18950
rect 10669 18826 12481 18894
rect 10669 18770 10679 18826
rect 10735 18770 10803 18826
rect 10859 18770 10927 18826
rect 10983 18770 11051 18826
rect 11107 18770 11175 18826
rect 11231 18770 11299 18826
rect 11355 18770 11423 18826
rect 11479 18770 11547 18826
rect 11603 18770 11671 18826
rect 11727 18770 11795 18826
rect 11851 18770 11919 18826
rect 11975 18770 12043 18826
rect 12099 18770 12167 18826
rect 12223 18770 12291 18826
rect 12347 18770 12415 18826
rect 12471 18770 12481 18826
rect 10669 18702 12481 18770
rect 10669 18646 10679 18702
rect 10735 18646 10803 18702
rect 10859 18646 10927 18702
rect 10983 18646 11051 18702
rect 11107 18646 11175 18702
rect 11231 18646 11299 18702
rect 11355 18646 11423 18702
rect 11479 18646 11547 18702
rect 11603 18646 11671 18702
rect 11727 18646 11795 18702
rect 11851 18646 11919 18702
rect 11975 18646 12043 18702
rect 12099 18646 12167 18702
rect 12223 18646 12291 18702
rect 12347 18646 12415 18702
rect 12471 18646 12481 18702
rect 10669 18578 12481 18646
rect 10669 18522 10679 18578
rect 10735 18522 10803 18578
rect 10859 18522 10927 18578
rect 10983 18522 11051 18578
rect 11107 18522 11175 18578
rect 11231 18522 11299 18578
rect 11355 18522 11423 18578
rect 11479 18522 11547 18578
rect 11603 18522 11671 18578
rect 11727 18522 11795 18578
rect 11851 18522 11919 18578
rect 11975 18522 12043 18578
rect 12099 18522 12167 18578
rect 12223 18522 12291 18578
rect 12347 18522 12415 18578
rect 12471 18522 12481 18578
rect 10669 18454 12481 18522
rect 10669 18398 10679 18454
rect 10735 18398 10803 18454
rect 10859 18398 10927 18454
rect 10983 18398 11051 18454
rect 11107 18398 11175 18454
rect 11231 18398 11299 18454
rect 11355 18398 11423 18454
rect 11479 18398 11547 18454
rect 11603 18398 11671 18454
rect 11727 18398 11795 18454
rect 11851 18398 11919 18454
rect 11975 18398 12043 18454
rect 12099 18398 12167 18454
rect 12223 18398 12291 18454
rect 12347 18398 12415 18454
rect 12471 18398 12481 18454
rect 10669 18330 12481 18398
rect 10669 18274 10679 18330
rect 10735 18274 10803 18330
rect 10859 18274 10927 18330
rect 10983 18274 11051 18330
rect 11107 18274 11175 18330
rect 11231 18274 11299 18330
rect 11355 18274 11423 18330
rect 11479 18274 11547 18330
rect 11603 18274 11671 18330
rect 11727 18274 11795 18330
rect 11851 18274 11919 18330
rect 11975 18274 12043 18330
rect 12099 18274 12167 18330
rect 12223 18274 12291 18330
rect 12347 18274 12415 18330
rect 12471 18274 12481 18330
rect 10669 18206 12481 18274
rect 10669 18150 10679 18206
rect 10735 18150 10803 18206
rect 10859 18150 10927 18206
rect 10983 18150 11051 18206
rect 11107 18150 11175 18206
rect 11231 18150 11299 18206
rect 11355 18150 11423 18206
rect 11479 18150 11547 18206
rect 11603 18150 11671 18206
rect 11727 18150 11795 18206
rect 11851 18150 11919 18206
rect 11975 18150 12043 18206
rect 12099 18150 12167 18206
rect 12223 18150 12291 18206
rect 12347 18150 12415 18206
rect 12471 18150 12481 18206
rect 10669 18082 12481 18150
rect 10669 18026 10679 18082
rect 10735 18026 10803 18082
rect 10859 18026 10927 18082
rect 10983 18026 11051 18082
rect 11107 18026 11175 18082
rect 11231 18026 11299 18082
rect 11355 18026 11423 18082
rect 11479 18026 11547 18082
rect 11603 18026 11671 18082
rect 11727 18026 11795 18082
rect 11851 18026 11919 18082
rect 11975 18026 12043 18082
rect 12099 18026 12167 18082
rect 12223 18026 12291 18082
rect 12347 18026 12415 18082
rect 12471 18026 12481 18082
rect 10669 17958 12481 18026
rect 10669 17902 10679 17958
rect 10735 17902 10803 17958
rect 10859 17902 10927 17958
rect 10983 17902 11051 17958
rect 11107 17902 11175 17958
rect 11231 17902 11299 17958
rect 11355 17902 11423 17958
rect 11479 17902 11547 17958
rect 11603 17902 11671 17958
rect 11727 17902 11795 17958
rect 11851 17902 11919 17958
rect 11975 17902 12043 17958
rect 12099 17902 12167 17958
rect 12223 17902 12291 17958
rect 12347 17902 12415 17958
rect 12471 17902 12481 17958
rect 10669 17834 12481 17902
rect 10669 17778 10679 17834
rect 10735 17778 10803 17834
rect 10859 17778 10927 17834
rect 10983 17778 11051 17834
rect 11107 17778 11175 17834
rect 11231 17778 11299 17834
rect 11355 17778 11423 17834
rect 11479 17778 11547 17834
rect 11603 17778 11671 17834
rect 11727 17778 11795 17834
rect 11851 17778 11919 17834
rect 11975 17778 12043 17834
rect 12099 17778 12167 17834
rect 12223 17778 12291 17834
rect 12347 17778 12415 17834
rect 12471 17778 12481 17834
rect 10669 17710 12481 17778
rect 10669 17654 10679 17710
rect 10735 17654 10803 17710
rect 10859 17654 10927 17710
rect 10983 17654 11051 17710
rect 11107 17654 11175 17710
rect 11231 17654 11299 17710
rect 11355 17654 11423 17710
rect 11479 17654 11547 17710
rect 11603 17654 11671 17710
rect 11727 17654 11795 17710
rect 11851 17654 11919 17710
rect 11975 17654 12043 17710
rect 12099 17654 12167 17710
rect 12223 17654 12291 17710
rect 12347 17654 12415 17710
rect 12471 17654 12481 17710
rect 10669 17586 12481 17654
rect 10669 17530 10679 17586
rect 10735 17530 10803 17586
rect 10859 17530 10927 17586
rect 10983 17530 11051 17586
rect 11107 17530 11175 17586
rect 11231 17530 11299 17586
rect 11355 17530 11423 17586
rect 11479 17530 11547 17586
rect 11603 17530 11671 17586
rect 11727 17530 11795 17586
rect 11851 17530 11919 17586
rect 11975 17530 12043 17586
rect 12099 17530 12167 17586
rect 12223 17530 12291 17586
rect 12347 17530 12415 17586
rect 12471 17530 12481 17586
rect 10669 17462 12481 17530
rect 10669 17406 10679 17462
rect 10735 17406 10803 17462
rect 10859 17406 10927 17462
rect 10983 17406 11051 17462
rect 11107 17406 11175 17462
rect 11231 17406 11299 17462
rect 11355 17406 11423 17462
rect 11479 17406 11547 17462
rect 11603 17406 11671 17462
rect 11727 17406 11795 17462
rect 11851 17406 11919 17462
rect 11975 17406 12043 17462
rect 12099 17406 12167 17462
rect 12223 17406 12291 17462
rect 12347 17406 12415 17462
rect 12471 17406 12481 17462
rect 10669 17338 12481 17406
rect 10669 17282 10679 17338
rect 10735 17282 10803 17338
rect 10859 17282 10927 17338
rect 10983 17282 11051 17338
rect 11107 17282 11175 17338
rect 11231 17282 11299 17338
rect 11355 17282 11423 17338
rect 11479 17282 11547 17338
rect 11603 17282 11671 17338
rect 11727 17282 11795 17338
rect 11851 17282 11919 17338
rect 11975 17282 12043 17338
rect 12099 17282 12167 17338
rect 12223 17282 12291 17338
rect 12347 17282 12415 17338
rect 12471 17282 12481 17338
rect 10669 17214 12481 17282
rect 10669 17158 10679 17214
rect 10735 17158 10803 17214
rect 10859 17158 10927 17214
rect 10983 17158 11051 17214
rect 11107 17158 11175 17214
rect 11231 17158 11299 17214
rect 11355 17158 11423 17214
rect 11479 17158 11547 17214
rect 11603 17158 11671 17214
rect 11727 17158 11795 17214
rect 11851 17158 11919 17214
rect 11975 17158 12043 17214
rect 12099 17158 12167 17214
rect 12223 17158 12291 17214
rect 12347 17158 12415 17214
rect 12471 17158 12481 17214
rect 10669 17090 12481 17158
rect 10669 17034 10679 17090
rect 10735 17034 10803 17090
rect 10859 17034 10927 17090
rect 10983 17034 11051 17090
rect 11107 17034 11175 17090
rect 11231 17034 11299 17090
rect 11355 17034 11423 17090
rect 11479 17034 11547 17090
rect 11603 17034 11671 17090
rect 11727 17034 11795 17090
rect 11851 17034 11919 17090
rect 11975 17034 12043 17090
rect 12099 17034 12167 17090
rect 12223 17034 12291 17090
rect 12347 17034 12415 17090
rect 12471 17034 12481 17090
rect 10669 16966 12481 17034
rect 10669 16910 10679 16966
rect 10735 16910 10803 16966
rect 10859 16910 10927 16966
rect 10983 16910 11051 16966
rect 11107 16910 11175 16966
rect 11231 16910 11299 16966
rect 11355 16910 11423 16966
rect 11479 16910 11547 16966
rect 11603 16910 11671 16966
rect 11727 16910 11795 16966
rect 11851 16910 11919 16966
rect 11975 16910 12043 16966
rect 12099 16910 12167 16966
rect 12223 16910 12291 16966
rect 12347 16910 12415 16966
rect 12471 16910 12481 16966
rect 10669 16842 12481 16910
rect 10669 16786 10679 16842
rect 10735 16786 10803 16842
rect 10859 16786 10927 16842
rect 10983 16786 11051 16842
rect 11107 16786 11175 16842
rect 11231 16786 11299 16842
rect 11355 16786 11423 16842
rect 11479 16786 11547 16842
rect 11603 16786 11671 16842
rect 11727 16786 11795 16842
rect 11851 16786 11919 16842
rect 11975 16786 12043 16842
rect 12099 16786 12167 16842
rect 12223 16786 12291 16842
rect 12347 16786 12415 16842
rect 12471 16786 12481 16842
rect 10669 16718 12481 16786
rect 10669 16662 10679 16718
rect 10735 16662 10803 16718
rect 10859 16662 10927 16718
rect 10983 16662 11051 16718
rect 11107 16662 11175 16718
rect 11231 16662 11299 16718
rect 11355 16662 11423 16718
rect 11479 16662 11547 16718
rect 11603 16662 11671 16718
rect 11727 16662 11795 16718
rect 11851 16662 11919 16718
rect 11975 16662 12043 16718
rect 12099 16662 12167 16718
rect 12223 16662 12291 16718
rect 12347 16662 12415 16718
rect 12471 16662 12481 16718
rect 10669 16594 12481 16662
rect 10669 16538 10679 16594
rect 10735 16538 10803 16594
rect 10859 16538 10927 16594
rect 10983 16538 11051 16594
rect 11107 16538 11175 16594
rect 11231 16538 11299 16594
rect 11355 16538 11423 16594
rect 11479 16538 11547 16594
rect 11603 16538 11671 16594
rect 11727 16538 11795 16594
rect 11851 16538 11919 16594
rect 11975 16538 12043 16594
rect 12099 16538 12167 16594
rect 12223 16538 12291 16594
rect 12347 16538 12415 16594
rect 12471 16538 12481 16594
rect 10669 16470 12481 16538
rect 10669 16414 10679 16470
rect 10735 16414 10803 16470
rect 10859 16414 10927 16470
rect 10983 16414 11051 16470
rect 11107 16414 11175 16470
rect 11231 16414 11299 16470
rect 11355 16414 11423 16470
rect 11479 16414 11547 16470
rect 11603 16414 11671 16470
rect 11727 16414 11795 16470
rect 11851 16414 11919 16470
rect 11975 16414 12043 16470
rect 12099 16414 12167 16470
rect 12223 16414 12291 16470
rect 12347 16414 12415 16470
rect 12471 16414 12481 16470
rect 10669 16346 12481 16414
rect 10669 16290 10679 16346
rect 10735 16290 10803 16346
rect 10859 16290 10927 16346
rect 10983 16290 11051 16346
rect 11107 16290 11175 16346
rect 11231 16290 11299 16346
rect 11355 16290 11423 16346
rect 11479 16290 11547 16346
rect 11603 16290 11671 16346
rect 11727 16290 11795 16346
rect 11851 16290 11919 16346
rect 11975 16290 12043 16346
rect 12099 16290 12167 16346
rect 12223 16290 12291 16346
rect 12347 16290 12415 16346
rect 12471 16290 12481 16346
rect 10669 16222 12481 16290
rect 10669 16166 10679 16222
rect 10735 16166 10803 16222
rect 10859 16166 10927 16222
rect 10983 16166 11051 16222
rect 11107 16166 11175 16222
rect 11231 16166 11299 16222
rect 11355 16166 11423 16222
rect 11479 16166 11547 16222
rect 11603 16166 11671 16222
rect 11727 16166 11795 16222
rect 11851 16166 11919 16222
rect 11975 16166 12043 16222
rect 12099 16166 12167 16222
rect 12223 16166 12291 16222
rect 12347 16166 12415 16222
rect 12471 16166 12481 16222
rect 10669 16098 12481 16166
rect 10669 16042 10679 16098
rect 10735 16042 10803 16098
rect 10859 16042 10927 16098
rect 10983 16042 11051 16098
rect 11107 16042 11175 16098
rect 11231 16042 11299 16098
rect 11355 16042 11423 16098
rect 11479 16042 11547 16098
rect 11603 16042 11671 16098
rect 11727 16042 11795 16098
rect 11851 16042 11919 16098
rect 11975 16042 12043 16098
rect 12099 16042 12167 16098
rect 12223 16042 12291 16098
rect 12347 16042 12415 16098
rect 12471 16042 12481 16098
rect 10669 16032 12481 16042
rect 1068 15750 2136 15760
rect 1068 15694 1078 15750
rect 1134 15694 1202 15750
rect 1258 15694 1326 15750
rect 1382 15694 1450 15750
rect 1506 15694 1574 15750
rect 1630 15694 1698 15750
rect 1754 15694 1822 15750
rect 1878 15694 1946 15750
rect 2002 15694 2070 15750
rect 2126 15694 2136 15750
rect 1068 15626 2136 15694
rect 1068 15570 1078 15626
rect 1134 15570 1202 15626
rect 1258 15570 1326 15626
rect 1382 15570 1450 15626
rect 1506 15570 1574 15626
rect 1630 15570 1698 15626
rect 1754 15570 1822 15626
rect 1878 15570 1946 15626
rect 2002 15570 2070 15626
rect 2126 15570 2136 15626
rect 1068 15502 2136 15570
rect 1068 15446 1078 15502
rect 1134 15446 1202 15502
rect 1258 15446 1326 15502
rect 1382 15446 1450 15502
rect 1506 15446 1574 15502
rect 1630 15446 1698 15502
rect 1754 15446 1822 15502
rect 1878 15446 1946 15502
rect 2002 15446 2070 15502
rect 2126 15446 2136 15502
rect 1068 15378 2136 15446
rect 1068 15322 1078 15378
rect 1134 15322 1202 15378
rect 1258 15322 1326 15378
rect 1382 15322 1450 15378
rect 1506 15322 1574 15378
rect 1630 15322 1698 15378
rect 1754 15322 1822 15378
rect 1878 15322 1946 15378
rect 2002 15322 2070 15378
rect 2126 15322 2136 15378
rect 1068 15254 2136 15322
rect 1068 15198 1078 15254
rect 1134 15198 1202 15254
rect 1258 15198 1326 15254
rect 1382 15198 1450 15254
rect 1506 15198 1574 15254
rect 1630 15198 1698 15254
rect 1754 15198 1822 15254
rect 1878 15198 1946 15254
rect 2002 15198 2070 15254
rect 2126 15198 2136 15254
rect 1068 15130 2136 15198
rect 1068 15074 1078 15130
rect 1134 15074 1202 15130
rect 1258 15074 1326 15130
rect 1382 15074 1450 15130
rect 1506 15074 1574 15130
rect 1630 15074 1698 15130
rect 1754 15074 1822 15130
rect 1878 15074 1946 15130
rect 2002 15074 2070 15130
rect 2126 15074 2136 15130
rect 1068 15006 2136 15074
rect 1068 14950 1078 15006
rect 1134 14950 1202 15006
rect 1258 14950 1326 15006
rect 1382 14950 1450 15006
rect 1506 14950 1574 15006
rect 1630 14950 1698 15006
rect 1754 14950 1822 15006
rect 1878 14950 1946 15006
rect 2002 14950 2070 15006
rect 2126 14950 2136 15006
rect 1068 14882 2136 14950
rect 1068 14826 1078 14882
rect 1134 14826 1202 14882
rect 1258 14826 1326 14882
rect 1382 14826 1450 14882
rect 1506 14826 1574 14882
rect 1630 14826 1698 14882
rect 1754 14826 1822 14882
rect 1878 14826 1946 14882
rect 2002 14826 2070 14882
rect 2126 14826 2136 14882
rect 1068 14758 2136 14826
rect 1068 14702 1078 14758
rect 1134 14702 1202 14758
rect 1258 14702 1326 14758
rect 1382 14702 1450 14758
rect 1506 14702 1574 14758
rect 1630 14702 1698 14758
rect 1754 14702 1822 14758
rect 1878 14702 1946 14758
rect 2002 14702 2070 14758
rect 2126 14702 2136 14758
rect 1068 14634 2136 14702
rect 1068 14578 1078 14634
rect 1134 14578 1202 14634
rect 1258 14578 1326 14634
rect 1382 14578 1450 14634
rect 1506 14578 1574 14634
rect 1630 14578 1698 14634
rect 1754 14578 1822 14634
rect 1878 14578 1946 14634
rect 2002 14578 2070 14634
rect 2126 14578 2136 14634
rect 1068 14510 2136 14578
rect 1068 14454 1078 14510
rect 1134 14454 1202 14510
rect 1258 14454 1326 14510
rect 1382 14454 1450 14510
rect 1506 14454 1574 14510
rect 1630 14454 1698 14510
rect 1754 14454 1822 14510
rect 1878 14454 1946 14510
rect 2002 14454 2070 14510
rect 2126 14454 2136 14510
rect 1068 14386 2136 14454
rect 1068 14330 1078 14386
rect 1134 14330 1202 14386
rect 1258 14330 1326 14386
rect 1382 14330 1450 14386
rect 1506 14330 1574 14386
rect 1630 14330 1698 14386
rect 1754 14330 1822 14386
rect 1878 14330 1946 14386
rect 2002 14330 2070 14386
rect 2126 14330 2136 14386
rect 1068 14262 2136 14330
rect 1068 14206 1078 14262
rect 1134 14206 1202 14262
rect 1258 14206 1326 14262
rect 1382 14206 1450 14262
rect 1506 14206 1574 14262
rect 1630 14206 1698 14262
rect 1754 14206 1822 14262
rect 1878 14206 1946 14262
rect 2002 14206 2070 14262
rect 2126 14206 2136 14262
rect 1068 14138 2136 14206
rect 1068 14082 1078 14138
rect 1134 14082 1202 14138
rect 1258 14082 1326 14138
rect 1382 14082 1450 14138
rect 1506 14082 1574 14138
rect 1630 14082 1698 14138
rect 1754 14082 1822 14138
rect 1878 14082 1946 14138
rect 2002 14082 2070 14138
rect 2126 14082 2136 14138
rect 1068 14014 2136 14082
rect 1068 13958 1078 14014
rect 1134 13958 1202 14014
rect 1258 13958 1326 14014
rect 1382 13958 1450 14014
rect 1506 13958 1574 14014
rect 1630 13958 1698 14014
rect 1754 13958 1822 14014
rect 1878 13958 1946 14014
rect 2002 13958 2070 14014
rect 2126 13958 2136 14014
rect 1068 13890 2136 13958
rect 1068 13834 1078 13890
rect 1134 13834 1202 13890
rect 1258 13834 1326 13890
rect 1382 13834 1450 13890
rect 1506 13834 1574 13890
rect 1630 13834 1698 13890
rect 1754 13834 1822 13890
rect 1878 13834 1946 13890
rect 2002 13834 2070 13890
rect 2126 13834 2136 13890
rect 1068 13766 2136 13834
rect 1068 13710 1078 13766
rect 1134 13710 1202 13766
rect 1258 13710 1326 13766
rect 1382 13710 1450 13766
rect 1506 13710 1574 13766
rect 1630 13710 1698 13766
rect 1754 13710 1822 13766
rect 1878 13710 1946 13766
rect 2002 13710 2070 13766
rect 2126 13710 2136 13766
rect 1068 13642 2136 13710
rect 1068 13586 1078 13642
rect 1134 13586 1202 13642
rect 1258 13586 1326 13642
rect 1382 13586 1450 13642
rect 1506 13586 1574 13642
rect 1630 13586 1698 13642
rect 1754 13586 1822 13642
rect 1878 13586 1946 13642
rect 2002 13586 2070 13642
rect 2126 13586 2136 13642
rect 1068 13518 2136 13586
rect 1068 13462 1078 13518
rect 1134 13462 1202 13518
rect 1258 13462 1326 13518
rect 1382 13462 1450 13518
rect 1506 13462 1574 13518
rect 1630 13462 1698 13518
rect 1754 13462 1822 13518
rect 1878 13462 1946 13518
rect 2002 13462 2070 13518
rect 2126 13462 2136 13518
rect 1068 13394 2136 13462
rect 1068 13338 1078 13394
rect 1134 13338 1202 13394
rect 1258 13338 1326 13394
rect 1382 13338 1450 13394
rect 1506 13338 1574 13394
rect 1630 13338 1698 13394
rect 1754 13338 1822 13394
rect 1878 13338 1946 13394
rect 2002 13338 2070 13394
rect 2126 13338 2136 13394
rect 1068 13270 2136 13338
rect 1068 13214 1078 13270
rect 1134 13214 1202 13270
rect 1258 13214 1326 13270
rect 1382 13214 1450 13270
rect 1506 13214 1574 13270
rect 1630 13214 1698 13270
rect 1754 13214 1822 13270
rect 1878 13214 1946 13270
rect 2002 13214 2070 13270
rect 2126 13214 2136 13270
rect 1068 13146 2136 13214
rect 1068 13090 1078 13146
rect 1134 13090 1202 13146
rect 1258 13090 1326 13146
rect 1382 13090 1450 13146
rect 1506 13090 1574 13146
rect 1630 13090 1698 13146
rect 1754 13090 1822 13146
rect 1878 13090 1946 13146
rect 2002 13090 2070 13146
rect 2126 13090 2136 13146
rect 1068 13022 2136 13090
rect 1068 12966 1078 13022
rect 1134 12966 1202 13022
rect 1258 12966 1326 13022
rect 1382 12966 1450 13022
rect 1506 12966 1574 13022
rect 1630 12966 1698 13022
rect 1754 12966 1822 13022
rect 1878 12966 1946 13022
rect 2002 12966 2070 13022
rect 2126 12966 2136 13022
rect 1068 12898 2136 12966
rect 1068 12842 1078 12898
rect 1134 12842 1202 12898
rect 1258 12842 1326 12898
rect 1382 12842 1450 12898
rect 1506 12842 1574 12898
rect 1630 12842 1698 12898
rect 1754 12842 1822 12898
rect 1878 12842 1946 12898
rect 2002 12842 2070 12898
rect 2126 12842 2136 12898
rect 1068 12832 2136 12842
rect 4425 15750 6237 15760
rect 4425 15694 4435 15750
rect 4491 15694 4559 15750
rect 4615 15694 4683 15750
rect 4739 15694 4807 15750
rect 4863 15694 4931 15750
rect 4987 15694 5055 15750
rect 5111 15694 5179 15750
rect 5235 15694 5303 15750
rect 5359 15694 5427 15750
rect 5483 15694 5551 15750
rect 5607 15694 5675 15750
rect 5731 15694 5799 15750
rect 5855 15694 5923 15750
rect 5979 15694 6047 15750
rect 6103 15694 6171 15750
rect 6227 15694 6237 15750
rect 4425 15626 6237 15694
rect 4425 15570 4435 15626
rect 4491 15570 4559 15626
rect 4615 15570 4683 15626
rect 4739 15570 4807 15626
rect 4863 15570 4931 15626
rect 4987 15570 5055 15626
rect 5111 15570 5179 15626
rect 5235 15570 5303 15626
rect 5359 15570 5427 15626
rect 5483 15570 5551 15626
rect 5607 15570 5675 15626
rect 5731 15570 5799 15626
rect 5855 15570 5923 15626
rect 5979 15570 6047 15626
rect 6103 15570 6171 15626
rect 6227 15570 6237 15626
rect 4425 15502 6237 15570
rect 4425 15446 4435 15502
rect 4491 15446 4559 15502
rect 4615 15446 4683 15502
rect 4739 15446 4807 15502
rect 4863 15446 4931 15502
rect 4987 15446 5055 15502
rect 5111 15446 5179 15502
rect 5235 15446 5303 15502
rect 5359 15446 5427 15502
rect 5483 15446 5551 15502
rect 5607 15446 5675 15502
rect 5731 15446 5799 15502
rect 5855 15446 5923 15502
rect 5979 15446 6047 15502
rect 6103 15446 6171 15502
rect 6227 15446 6237 15502
rect 4425 15378 6237 15446
rect 4425 15322 4435 15378
rect 4491 15322 4559 15378
rect 4615 15322 4683 15378
rect 4739 15322 4807 15378
rect 4863 15322 4931 15378
rect 4987 15322 5055 15378
rect 5111 15322 5179 15378
rect 5235 15322 5303 15378
rect 5359 15322 5427 15378
rect 5483 15322 5551 15378
rect 5607 15322 5675 15378
rect 5731 15322 5799 15378
rect 5855 15322 5923 15378
rect 5979 15322 6047 15378
rect 6103 15322 6171 15378
rect 6227 15322 6237 15378
rect 4425 15254 6237 15322
rect 4425 15198 4435 15254
rect 4491 15198 4559 15254
rect 4615 15198 4683 15254
rect 4739 15198 4807 15254
rect 4863 15198 4931 15254
rect 4987 15198 5055 15254
rect 5111 15198 5179 15254
rect 5235 15198 5303 15254
rect 5359 15198 5427 15254
rect 5483 15198 5551 15254
rect 5607 15198 5675 15254
rect 5731 15198 5799 15254
rect 5855 15198 5923 15254
rect 5979 15198 6047 15254
rect 6103 15198 6171 15254
rect 6227 15198 6237 15254
rect 4425 15130 6237 15198
rect 4425 15074 4435 15130
rect 4491 15074 4559 15130
rect 4615 15074 4683 15130
rect 4739 15074 4807 15130
rect 4863 15074 4931 15130
rect 4987 15074 5055 15130
rect 5111 15074 5179 15130
rect 5235 15074 5303 15130
rect 5359 15074 5427 15130
rect 5483 15074 5551 15130
rect 5607 15074 5675 15130
rect 5731 15074 5799 15130
rect 5855 15074 5923 15130
rect 5979 15074 6047 15130
rect 6103 15074 6171 15130
rect 6227 15074 6237 15130
rect 4425 15006 6237 15074
rect 4425 14950 4435 15006
rect 4491 14950 4559 15006
rect 4615 14950 4683 15006
rect 4739 14950 4807 15006
rect 4863 14950 4931 15006
rect 4987 14950 5055 15006
rect 5111 14950 5179 15006
rect 5235 14950 5303 15006
rect 5359 14950 5427 15006
rect 5483 14950 5551 15006
rect 5607 14950 5675 15006
rect 5731 14950 5799 15006
rect 5855 14950 5923 15006
rect 5979 14950 6047 15006
rect 6103 14950 6171 15006
rect 6227 14950 6237 15006
rect 4425 14882 6237 14950
rect 4425 14826 4435 14882
rect 4491 14826 4559 14882
rect 4615 14826 4683 14882
rect 4739 14826 4807 14882
rect 4863 14826 4931 14882
rect 4987 14826 5055 14882
rect 5111 14826 5179 14882
rect 5235 14826 5303 14882
rect 5359 14826 5427 14882
rect 5483 14826 5551 14882
rect 5607 14826 5675 14882
rect 5731 14826 5799 14882
rect 5855 14826 5923 14882
rect 5979 14826 6047 14882
rect 6103 14826 6171 14882
rect 6227 14826 6237 14882
rect 4425 14758 6237 14826
rect 4425 14702 4435 14758
rect 4491 14702 4559 14758
rect 4615 14702 4683 14758
rect 4739 14702 4807 14758
rect 4863 14702 4931 14758
rect 4987 14702 5055 14758
rect 5111 14702 5179 14758
rect 5235 14702 5303 14758
rect 5359 14702 5427 14758
rect 5483 14702 5551 14758
rect 5607 14702 5675 14758
rect 5731 14702 5799 14758
rect 5855 14702 5923 14758
rect 5979 14702 6047 14758
rect 6103 14702 6171 14758
rect 6227 14702 6237 14758
rect 4425 14634 6237 14702
rect 4425 14578 4435 14634
rect 4491 14578 4559 14634
rect 4615 14578 4683 14634
rect 4739 14578 4807 14634
rect 4863 14578 4931 14634
rect 4987 14578 5055 14634
rect 5111 14578 5179 14634
rect 5235 14578 5303 14634
rect 5359 14578 5427 14634
rect 5483 14578 5551 14634
rect 5607 14578 5675 14634
rect 5731 14578 5799 14634
rect 5855 14578 5923 14634
rect 5979 14578 6047 14634
rect 6103 14578 6171 14634
rect 6227 14578 6237 14634
rect 4425 14510 6237 14578
rect 4425 14454 4435 14510
rect 4491 14454 4559 14510
rect 4615 14454 4683 14510
rect 4739 14454 4807 14510
rect 4863 14454 4931 14510
rect 4987 14454 5055 14510
rect 5111 14454 5179 14510
rect 5235 14454 5303 14510
rect 5359 14454 5427 14510
rect 5483 14454 5551 14510
rect 5607 14454 5675 14510
rect 5731 14454 5799 14510
rect 5855 14454 5923 14510
rect 5979 14454 6047 14510
rect 6103 14454 6171 14510
rect 6227 14454 6237 14510
rect 4425 14386 6237 14454
rect 4425 14330 4435 14386
rect 4491 14330 4559 14386
rect 4615 14330 4683 14386
rect 4739 14330 4807 14386
rect 4863 14330 4931 14386
rect 4987 14330 5055 14386
rect 5111 14330 5179 14386
rect 5235 14330 5303 14386
rect 5359 14330 5427 14386
rect 5483 14330 5551 14386
rect 5607 14330 5675 14386
rect 5731 14330 5799 14386
rect 5855 14330 5923 14386
rect 5979 14330 6047 14386
rect 6103 14330 6171 14386
rect 6227 14330 6237 14386
rect 4425 14262 6237 14330
rect 4425 14206 4435 14262
rect 4491 14206 4559 14262
rect 4615 14206 4683 14262
rect 4739 14206 4807 14262
rect 4863 14206 4931 14262
rect 4987 14206 5055 14262
rect 5111 14206 5179 14262
rect 5235 14206 5303 14262
rect 5359 14206 5427 14262
rect 5483 14206 5551 14262
rect 5607 14206 5675 14262
rect 5731 14206 5799 14262
rect 5855 14206 5923 14262
rect 5979 14206 6047 14262
rect 6103 14206 6171 14262
rect 6227 14206 6237 14262
rect 4425 14138 6237 14206
rect 4425 14082 4435 14138
rect 4491 14082 4559 14138
rect 4615 14082 4683 14138
rect 4739 14082 4807 14138
rect 4863 14082 4931 14138
rect 4987 14082 5055 14138
rect 5111 14082 5179 14138
rect 5235 14082 5303 14138
rect 5359 14082 5427 14138
rect 5483 14082 5551 14138
rect 5607 14082 5675 14138
rect 5731 14082 5799 14138
rect 5855 14082 5923 14138
rect 5979 14082 6047 14138
rect 6103 14082 6171 14138
rect 6227 14082 6237 14138
rect 4425 14014 6237 14082
rect 4425 13958 4435 14014
rect 4491 13958 4559 14014
rect 4615 13958 4683 14014
rect 4739 13958 4807 14014
rect 4863 13958 4931 14014
rect 4987 13958 5055 14014
rect 5111 13958 5179 14014
rect 5235 13958 5303 14014
rect 5359 13958 5427 14014
rect 5483 13958 5551 14014
rect 5607 13958 5675 14014
rect 5731 13958 5799 14014
rect 5855 13958 5923 14014
rect 5979 13958 6047 14014
rect 6103 13958 6171 14014
rect 6227 13958 6237 14014
rect 4425 13890 6237 13958
rect 4425 13834 4435 13890
rect 4491 13834 4559 13890
rect 4615 13834 4683 13890
rect 4739 13834 4807 13890
rect 4863 13834 4931 13890
rect 4987 13834 5055 13890
rect 5111 13834 5179 13890
rect 5235 13834 5303 13890
rect 5359 13834 5427 13890
rect 5483 13834 5551 13890
rect 5607 13834 5675 13890
rect 5731 13834 5799 13890
rect 5855 13834 5923 13890
rect 5979 13834 6047 13890
rect 6103 13834 6171 13890
rect 6227 13834 6237 13890
rect 4425 13766 6237 13834
rect 4425 13710 4435 13766
rect 4491 13710 4559 13766
rect 4615 13710 4683 13766
rect 4739 13710 4807 13766
rect 4863 13710 4931 13766
rect 4987 13710 5055 13766
rect 5111 13710 5179 13766
rect 5235 13710 5303 13766
rect 5359 13710 5427 13766
rect 5483 13710 5551 13766
rect 5607 13710 5675 13766
rect 5731 13710 5799 13766
rect 5855 13710 5923 13766
rect 5979 13710 6047 13766
rect 6103 13710 6171 13766
rect 6227 13710 6237 13766
rect 4425 13642 6237 13710
rect 4425 13586 4435 13642
rect 4491 13586 4559 13642
rect 4615 13586 4683 13642
rect 4739 13586 4807 13642
rect 4863 13586 4931 13642
rect 4987 13586 5055 13642
rect 5111 13586 5179 13642
rect 5235 13586 5303 13642
rect 5359 13586 5427 13642
rect 5483 13586 5551 13642
rect 5607 13586 5675 13642
rect 5731 13586 5799 13642
rect 5855 13586 5923 13642
rect 5979 13586 6047 13642
rect 6103 13586 6171 13642
rect 6227 13586 6237 13642
rect 4425 13518 6237 13586
rect 4425 13462 4435 13518
rect 4491 13462 4559 13518
rect 4615 13462 4683 13518
rect 4739 13462 4807 13518
rect 4863 13462 4931 13518
rect 4987 13462 5055 13518
rect 5111 13462 5179 13518
rect 5235 13462 5303 13518
rect 5359 13462 5427 13518
rect 5483 13462 5551 13518
rect 5607 13462 5675 13518
rect 5731 13462 5799 13518
rect 5855 13462 5923 13518
rect 5979 13462 6047 13518
rect 6103 13462 6171 13518
rect 6227 13462 6237 13518
rect 4425 13394 6237 13462
rect 4425 13338 4435 13394
rect 4491 13338 4559 13394
rect 4615 13338 4683 13394
rect 4739 13338 4807 13394
rect 4863 13338 4931 13394
rect 4987 13338 5055 13394
rect 5111 13338 5179 13394
rect 5235 13338 5303 13394
rect 5359 13338 5427 13394
rect 5483 13338 5551 13394
rect 5607 13338 5675 13394
rect 5731 13338 5799 13394
rect 5855 13338 5923 13394
rect 5979 13338 6047 13394
rect 6103 13338 6171 13394
rect 6227 13338 6237 13394
rect 4425 13270 6237 13338
rect 4425 13214 4435 13270
rect 4491 13214 4559 13270
rect 4615 13214 4683 13270
rect 4739 13214 4807 13270
rect 4863 13214 4931 13270
rect 4987 13214 5055 13270
rect 5111 13214 5179 13270
rect 5235 13214 5303 13270
rect 5359 13214 5427 13270
rect 5483 13214 5551 13270
rect 5607 13214 5675 13270
rect 5731 13214 5799 13270
rect 5855 13214 5923 13270
rect 5979 13214 6047 13270
rect 6103 13214 6171 13270
rect 6227 13214 6237 13270
rect 4425 13146 6237 13214
rect 4425 13090 4435 13146
rect 4491 13090 4559 13146
rect 4615 13090 4683 13146
rect 4739 13090 4807 13146
rect 4863 13090 4931 13146
rect 4987 13090 5055 13146
rect 5111 13090 5179 13146
rect 5235 13090 5303 13146
rect 5359 13090 5427 13146
rect 5483 13090 5551 13146
rect 5607 13090 5675 13146
rect 5731 13090 5799 13146
rect 5855 13090 5923 13146
rect 5979 13090 6047 13146
rect 6103 13090 6171 13146
rect 6227 13090 6237 13146
rect 4425 13022 6237 13090
rect 4425 12966 4435 13022
rect 4491 12966 4559 13022
rect 4615 12966 4683 13022
rect 4739 12966 4807 13022
rect 4863 12966 4931 13022
rect 4987 12966 5055 13022
rect 5111 12966 5179 13022
rect 5235 12966 5303 13022
rect 5359 12966 5427 13022
rect 5483 12966 5551 13022
rect 5607 12966 5675 13022
rect 5731 12966 5799 13022
rect 5855 12966 5923 13022
rect 5979 12966 6047 13022
rect 6103 12966 6171 13022
rect 6227 12966 6237 13022
rect 4425 12898 6237 12966
rect 4425 12842 4435 12898
rect 4491 12842 4559 12898
rect 4615 12842 4683 12898
rect 4739 12842 4807 12898
rect 4863 12842 4931 12898
rect 4987 12842 5055 12898
rect 5111 12842 5179 12898
rect 5235 12842 5303 12898
rect 5359 12842 5427 12898
rect 5483 12842 5551 12898
rect 5607 12842 5675 12898
rect 5731 12842 5799 12898
rect 5855 12842 5923 12898
rect 5979 12842 6047 12898
rect 6103 12842 6171 12898
rect 6227 12842 6237 12898
rect 4425 12832 6237 12842
rect 7552 15750 8620 15760
rect 7552 15694 7562 15750
rect 7618 15694 7686 15750
rect 7742 15694 7810 15750
rect 7866 15694 7934 15750
rect 7990 15694 8058 15750
rect 8114 15694 8182 15750
rect 8238 15694 8306 15750
rect 8362 15694 8430 15750
rect 8486 15694 8554 15750
rect 8610 15694 8620 15750
rect 7552 15626 8620 15694
rect 7552 15570 7562 15626
rect 7618 15570 7686 15626
rect 7742 15570 7810 15626
rect 7866 15570 7934 15626
rect 7990 15570 8058 15626
rect 8114 15570 8182 15626
rect 8238 15570 8306 15626
rect 8362 15570 8430 15626
rect 8486 15570 8554 15626
rect 8610 15570 8620 15626
rect 7552 15502 8620 15570
rect 7552 15446 7562 15502
rect 7618 15446 7686 15502
rect 7742 15446 7810 15502
rect 7866 15446 7934 15502
rect 7990 15446 8058 15502
rect 8114 15446 8182 15502
rect 8238 15446 8306 15502
rect 8362 15446 8430 15502
rect 8486 15446 8554 15502
rect 8610 15446 8620 15502
rect 7552 15378 8620 15446
rect 7552 15322 7562 15378
rect 7618 15322 7686 15378
rect 7742 15322 7810 15378
rect 7866 15322 7934 15378
rect 7990 15322 8058 15378
rect 8114 15322 8182 15378
rect 8238 15322 8306 15378
rect 8362 15322 8430 15378
rect 8486 15322 8554 15378
rect 8610 15322 8620 15378
rect 7552 15254 8620 15322
rect 7552 15198 7562 15254
rect 7618 15198 7686 15254
rect 7742 15198 7810 15254
rect 7866 15198 7934 15254
rect 7990 15198 8058 15254
rect 8114 15198 8182 15254
rect 8238 15198 8306 15254
rect 8362 15198 8430 15254
rect 8486 15198 8554 15254
rect 8610 15198 8620 15254
rect 7552 15130 8620 15198
rect 7552 15074 7562 15130
rect 7618 15074 7686 15130
rect 7742 15074 7810 15130
rect 7866 15074 7934 15130
rect 7990 15074 8058 15130
rect 8114 15074 8182 15130
rect 8238 15074 8306 15130
rect 8362 15074 8430 15130
rect 8486 15074 8554 15130
rect 8610 15074 8620 15130
rect 7552 15006 8620 15074
rect 7552 14950 7562 15006
rect 7618 14950 7686 15006
rect 7742 14950 7810 15006
rect 7866 14950 7934 15006
rect 7990 14950 8058 15006
rect 8114 14950 8182 15006
rect 8238 14950 8306 15006
rect 8362 14950 8430 15006
rect 8486 14950 8554 15006
rect 8610 14950 8620 15006
rect 7552 14882 8620 14950
rect 7552 14826 7562 14882
rect 7618 14826 7686 14882
rect 7742 14826 7810 14882
rect 7866 14826 7934 14882
rect 7990 14826 8058 14882
rect 8114 14826 8182 14882
rect 8238 14826 8306 14882
rect 8362 14826 8430 14882
rect 8486 14826 8554 14882
rect 8610 14826 8620 14882
rect 7552 14758 8620 14826
rect 7552 14702 7562 14758
rect 7618 14702 7686 14758
rect 7742 14702 7810 14758
rect 7866 14702 7934 14758
rect 7990 14702 8058 14758
rect 8114 14702 8182 14758
rect 8238 14702 8306 14758
rect 8362 14702 8430 14758
rect 8486 14702 8554 14758
rect 8610 14702 8620 14758
rect 7552 14634 8620 14702
rect 7552 14578 7562 14634
rect 7618 14578 7686 14634
rect 7742 14578 7810 14634
rect 7866 14578 7934 14634
rect 7990 14578 8058 14634
rect 8114 14578 8182 14634
rect 8238 14578 8306 14634
rect 8362 14578 8430 14634
rect 8486 14578 8554 14634
rect 8610 14578 8620 14634
rect 7552 14510 8620 14578
rect 7552 14454 7562 14510
rect 7618 14454 7686 14510
rect 7742 14454 7810 14510
rect 7866 14454 7934 14510
rect 7990 14454 8058 14510
rect 8114 14454 8182 14510
rect 8238 14454 8306 14510
rect 8362 14454 8430 14510
rect 8486 14454 8554 14510
rect 8610 14454 8620 14510
rect 7552 14386 8620 14454
rect 7552 14330 7562 14386
rect 7618 14330 7686 14386
rect 7742 14330 7810 14386
rect 7866 14330 7934 14386
rect 7990 14330 8058 14386
rect 8114 14330 8182 14386
rect 8238 14330 8306 14386
rect 8362 14330 8430 14386
rect 8486 14330 8554 14386
rect 8610 14330 8620 14386
rect 7552 14262 8620 14330
rect 7552 14206 7562 14262
rect 7618 14206 7686 14262
rect 7742 14206 7810 14262
rect 7866 14206 7934 14262
rect 7990 14206 8058 14262
rect 8114 14206 8182 14262
rect 8238 14206 8306 14262
rect 8362 14206 8430 14262
rect 8486 14206 8554 14262
rect 8610 14206 8620 14262
rect 7552 14138 8620 14206
rect 7552 14082 7562 14138
rect 7618 14082 7686 14138
rect 7742 14082 7810 14138
rect 7866 14082 7934 14138
rect 7990 14082 8058 14138
rect 8114 14082 8182 14138
rect 8238 14082 8306 14138
rect 8362 14082 8430 14138
rect 8486 14082 8554 14138
rect 8610 14082 8620 14138
rect 7552 14014 8620 14082
rect 7552 13958 7562 14014
rect 7618 13958 7686 14014
rect 7742 13958 7810 14014
rect 7866 13958 7934 14014
rect 7990 13958 8058 14014
rect 8114 13958 8182 14014
rect 8238 13958 8306 14014
rect 8362 13958 8430 14014
rect 8486 13958 8554 14014
rect 8610 13958 8620 14014
rect 7552 13890 8620 13958
rect 7552 13834 7562 13890
rect 7618 13834 7686 13890
rect 7742 13834 7810 13890
rect 7866 13834 7934 13890
rect 7990 13834 8058 13890
rect 8114 13834 8182 13890
rect 8238 13834 8306 13890
rect 8362 13834 8430 13890
rect 8486 13834 8554 13890
rect 8610 13834 8620 13890
rect 7552 13766 8620 13834
rect 7552 13710 7562 13766
rect 7618 13710 7686 13766
rect 7742 13710 7810 13766
rect 7866 13710 7934 13766
rect 7990 13710 8058 13766
rect 8114 13710 8182 13766
rect 8238 13710 8306 13766
rect 8362 13710 8430 13766
rect 8486 13710 8554 13766
rect 8610 13710 8620 13766
rect 7552 13642 8620 13710
rect 7552 13586 7562 13642
rect 7618 13586 7686 13642
rect 7742 13586 7810 13642
rect 7866 13586 7934 13642
rect 7990 13586 8058 13642
rect 8114 13586 8182 13642
rect 8238 13586 8306 13642
rect 8362 13586 8430 13642
rect 8486 13586 8554 13642
rect 8610 13586 8620 13642
rect 7552 13518 8620 13586
rect 7552 13462 7562 13518
rect 7618 13462 7686 13518
rect 7742 13462 7810 13518
rect 7866 13462 7934 13518
rect 7990 13462 8058 13518
rect 8114 13462 8182 13518
rect 8238 13462 8306 13518
rect 8362 13462 8430 13518
rect 8486 13462 8554 13518
rect 8610 13462 8620 13518
rect 7552 13394 8620 13462
rect 7552 13338 7562 13394
rect 7618 13338 7686 13394
rect 7742 13338 7810 13394
rect 7866 13338 7934 13394
rect 7990 13338 8058 13394
rect 8114 13338 8182 13394
rect 8238 13338 8306 13394
rect 8362 13338 8430 13394
rect 8486 13338 8554 13394
rect 8610 13338 8620 13394
rect 7552 13270 8620 13338
rect 7552 13214 7562 13270
rect 7618 13214 7686 13270
rect 7742 13214 7810 13270
rect 7866 13214 7934 13270
rect 7990 13214 8058 13270
rect 8114 13214 8182 13270
rect 8238 13214 8306 13270
rect 8362 13214 8430 13270
rect 8486 13214 8554 13270
rect 8610 13214 8620 13270
rect 7552 13146 8620 13214
rect 7552 13090 7562 13146
rect 7618 13090 7686 13146
rect 7742 13090 7810 13146
rect 7866 13090 7934 13146
rect 7990 13090 8058 13146
rect 8114 13090 8182 13146
rect 8238 13090 8306 13146
rect 8362 13090 8430 13146
rect 8486 13090 8554 13146
rect 8610 13090 8620 13146
rect 7552 13022 8620 13090
rect 7552 12966 7562 13022
rect 7618 12966 7686 13022
rect 7742 12966 7810 13022
rect 7866 12966 7934 13022
rect 7990 12966 8058 13022
rect 8114 12966 8182 13022
rect 8238 12966 8306 13022
rect 8362 12966 8430 13022
rect 8486 12966 8554 13022
rect 8610 12966 8620 13022
rect 7552 12898 8620 12966
rect 7552 12842 7562 12898
rect 7618 12842 7686 12898
rect 7742 12842 7810 12898
rect 7866 12842 7934 12898
rect 7990 12842 8058 12898
rect 8114 12842 8182 12898
rect 8238 12842 8306 12898
rect 8362 12842 8430 12898
rect 8486 12842 8554 12898
rect 8610 12842 8620 12898
rect 7552 12832 8620 12842
rect 10669 15750 12481 15760
rect 10669 15694 10679 15750
rect 10735 15694 10803 15750
rect 10859 15694 10927 15750
rect 10983 15694 11051 15750
rect 11107 15694 11175 15750
rect 11231 15694 11299 15750
rect 11355 15694 11423 15750
rect 11479 15694 11547 15750
rect 11603 15694 11671 15750
rect 11727 15694 11795 15750
rect 11851 15694 11919 15750
rect 11975 15694 12043 15750
rect 12099 15694 12167 15750
rect 12223 15694 12291 15750
rect 12347 15694 12415 15750
rect 12471 15694 12481 15750
rect 10669 15626 12481 15694
rect 10669 15570 10679 15626
rect 10735 15570 10803 15626
rect 10859 15570 10927 15626
rect 10983 15570 11051 15626
rect 11107 15570 11175 15626
rect 11231 15570 11299 15626
rect 11355 15570 11423 15626
rect 11479 15570 11547 15626
rect 11603 15570 11671 15626
rect 11727 15570 11795 15626
rect 11851 15570 11919 15626
rect 11975 15570 12043 15626
rect 12099 15570 12167 15626
rect 12223 15570 12291 15626
rect 12347 15570 12415 15626
rect 12471 15570 12481 15626
rect 10669 15502 12481 15570
rect 10669 15446 10679 15502
rect 10735 15446 10803 15502
rect 10859 15446 10927 15502
rect 10983 15446 11051 15502
rect 11107 15446 11175 15502
rect 11231 15446 11299 15502
rect 11355 15446 11423 15502
rect 11479 15446 11547 15502
rect 11603 15446 11671 15502
rect 11727 15446 11795 15502
rect 11851 15446 11919 15502
rect 11975 15446 12043 15502
rect 12099 15446 12167 15502
rect 12223 15446 12291 15502
rect 12347 15446 12415 15502
rect 12471 15446 12481 15502
rect 10669 15378 12481 15446
rect 10669 15322 10679 15378
rect 10735 15322 10803 15378
rect 10859 15322 10927 15378
rect 10983 15322 11051 15378
rect 11107 15322 11175 15378
rect 11231 15322 11299 15378
rect 11355 15322 11423 15378
rect 11479 15322 11547 15378
rect 11603 15322 11671 15378
rect 11727 15322 11795 15378
rect 11851 15322 11919 15378
rect 11975 15322 12043 15378
rect 12099 15322 12167 15378
rect 12223 15322 12291 15378
rect 12347 15322 12415 15378
rect 12471 15322 12481 15378
rect 10669 15254 12481 15322
rect 10669 15198 10679 15254
rect 10735 15198 10803 15254
rect 10859 15198 10927 15254
rect 10983 15198 11051 15254
rect 11107 15198 11175 15254
rect 11231 15198 11299 15254
rect 11355 15198 11423 15254
rect 11479 15198 11547 15254
rect 11603 15198 11671 15254
rect 11727 15198 11795 15254
rect 11851 15198 11919 15254
rect 11975 15198 12043 15254
rect 12099 15198 12167 15254
rect 12223 15198 12291 15254
rect 12347 15198 12415 15254
rect 12471 15198 12481 15254
rect 10669 15130 12481 15198
rect 10669 15074 10679 15130
rect 10735 15074 10803 15130
rect 10859 15074 10927 15130
rect 10983 15074 11051 15130
rect 11107 15074 11175 15130
rect 11231 15074 11299 15130
rect 11355 15074 11423 15130
rect 11479 15074 11547 15130
rect 11603 15074 11671 15130
rect 11727 15074 11795 15130
rect 11851 15074 11919 15130
rect 11975 15074 12043 15130
rect 12099 15074 12167 15130
rect 12223 15074 12291 15130
rect 12347 15074 12415 15130
rect 12471 15074 12481 15130
rect 10669 15006 12481 15074
rect 10669 14950 10679 15006
rect 10735 14950 10803 15006
rect 10859 14950 10927 15006
rect 10983 14950 11051 15006
rect 11107 14950 11175 15006
rect 11231 14950 11299 15006
rect 11355 14950 11423 15006
rect 11479 14950 11547 15006
rect 11603 14950 11671 15006
rect 11727 14950 11795 15006
rect 11851 14950 11919 15006
rect 11975 14950 12043 15006
rect 12099 14950 12167 15006
rect 12223 14950 12291 15006
rect 12347 14950 12415 15006
rect 12471 14950 12481 15006
rect 10669 14882 12481 14950
rect 10669 14826 10679 14882
rect 10735 14826 10803 14882
rect 10859 14826 10927 14882
rect 10983 14826 11051 14882
rect 11107 14826 11175 14882
rect 11231 14826 11299 14882
rect 11355 14826 11423 14882
rect 11479 14826 11547 14882
rect 11603 14826 11671 14882
rect 11727 14826 11795 14882
rect 11851 14826 11919 14882
rect 11975 14826 12043 14882
rect 12099 14826 12167 14882
rect 12223 14826 12291 14882
rect 12347 14826 12415 14882
rect 12471 14826 12481 14882
rect 10669 14758 12481 14826
rect 10669 14702 10679 14758
rect 10735 14702 10803 14758
rect 10859 14702 10927 14758
rect 10983 14702 11051 14758
rect 11107 14702 11175 14758
rect 11231 14702 11299 14758
rect 11355 14702 11423 14758
rect 11479 14702 11547 14758
rect 11603 14702 11671 14758
rect 11727 14702 11795 14758
rect 11851 14702 11919 14758
rect 11975 14702 12043 14758
rect 12099 14702 12167 14758
rect 12223 14702 12291 14758
rect 12347 14702 12415 14758
rect 12471 14702 12481 14758
rect 10669 14634 12481 14702
rect 10669 14578 10679 14634
rect 10735 14578 10803 14634
rect 10859 14578 10927 14634
rect 10983 14578 11051 14634
rect 11107 14578 11175 14634
rect 11231 14578 11299 14634
rect 11355 14578 11423 14634
rect 11479 14578 11547 14634
rect 11603 14578 11671 14634
rect 11727 14578 11795 14634
rect 11851 14578 11919 14634
rect 11975 14578 12043 14634
rect 12099 14578 12167 14634
rect 12223 14578 12291 14634
rect 12347 14578 12415 14634
rect 12471 14578 12481 14634
rect 10669 14510 12481 14578
rect 10669 14454 10679 14510
rect 10735 14454 10803 14510
rect 10859 14454 10927 14510
rect 10983 14454 11051 14510
rect 11107 14454 11175 14510
rect 11231 14454 11299 14510
rect 11355 14454 11423 14510
rect 11479 14454 11547 14510
rect 11603 14454 11671 14510
rect 11727 14454 11795 14510
rect 11851 14454 11919 14510
rect 11975 14454 12043 14510
rect 12099 14454 12167 14510
rect 12223 14454 12291 14510
rect 12347 14454 12415 14510
rect 12471 14454 12481 14510
rect 10669 14386 12481 14454
rect 10669 14330 10679 14386
rect 10735 14330 10803 14386
rect 10859 14330 10927 14386
rect 10983 14330 11051 14386
rect 11107 14330 11175 14386
rect 11231 14330 11299 14386
rect 11355 14330 11423 14386
rect 11479 14330 11547 14386
rect 11603 14330 11671 14386
rect 11727 14330 11795 14386
rect 11851 14330 11919 14386
rect 11975 14330 12043 14386
rect 12099 14330 12167 14386
rect 12223 14330 12291 14386
rect 12347 14330 12415 14386
rect 12471 14330 12481 14386
rect 10669 14262 12481 14330
rect 10669 14206 10679 14262
rect 10735 14206 10803 14262
rect 10859 14206 10927 14262
rect 10983 14206 11051 14262
rect 11107 14206 11175 14262
rect 11231 14206 11299 14262
rect 11355 14206 11423 14262
rect 11479 14206 11547 14262
rect 11603 14206 11671 14262
rect 11727 14206 11795 14262
rect 11851 14206 11919 14262
rect 11975 14206 12043 14262
rect 12099 14206 12167 14262
rect 12223 14206 12291 14262
rect 12347 14206 12415 14262
rect 12471 14206 12481 14262
rect 10669 14138 12481 14206
rect 10669 14082 10679 14138
rect 10735 14082 10803 14138
rect 10859 14082 10927 14138
rect 10983 14082 11051 14138
rect 11107 14082 11175 14138
rect 11231 14082 11299 14138
rect 11355 14082 11423 14138
rect 11479 14082 11547 14138
rect 11603 14082 11671 14138
rect 11727 14082 11795 14138
rect 11851 14082 11919 14138
rect 11975 14082 12043 14138
rect 12099 14082 12167 14138
rect 12223 14082 12291 14138
rect 12347 14082 12415 14138
rect 12471 14082 12481 14138
rect 10669 14014 12481 14082
rect 10669 13958 10679 14014
rect 10735 13958 10803 14014
rect 10859 13958 10927 14014
rect 10983 13958 11051 14014
rect 11107 13958 11175 14014
rect 11231 13958 11299 14014
rect 11355 13958 11423 14014
rect 11479 13958 11547 14014
rect 11603 13958 11671 14014
rect 11727 13958 11795 14014
rect 11851 13958 11919 14014
rect 11975 13958 12043 14014
rect 12099 13958 12167 14014
rect 12223 13958 12291 14014
rect 12347 13958 12415 14014
rect 12471 13958 12481 14014
rect 10669 13890 12481 13958
rect 10669 13834 10679 13890
rect 10735 13834 10803 13890
rect 10859 13834 10927 13890
rect 10983 13834 11051 13890
rect 11107 13834 11175 13890
rect 11231 13834 11299 13890
rect 11355 13834 11423 13890
rect 11479 13834 11547 13890
rect 11603 13834 11671 13890
rect 11727 13834 11795 13890
rect 11851 13834 11919 13890
rect 11975 13834 12043 13890
rect 12099 13834 12167 13890
rect 12223 13834 12291 13890
rect 12347 13834 12415 13890
rect 12471 13834 12481 13890
rect 10669 13766 12481 13834
rect 10669 13710 10679 13766
rect 10735 13710 10803 13766
rect 10859 13710 10927 13766
rect 10983 13710 11051 13766
rect 11107 13710 11175 13766
rect 11231 13710 11299 13766
rect 11355 13710 11423 13766
rect 11479 13710 11547 13766
rect 11603 13710 11671 13766
rect 11727 13710 11795 13766
rect 11851 13710 11919 13766
rect 11975 13710 12043 13766
rect 12099 13710 12167 13766
rect 12223 13710 12291 13766
rect 12347 13710 12415 13766
rect 12471 13710 12481 13766
rect 10669 13642 12481 13710
rect 10669 13586 10679 13642
rect 10735 13586 10803 13642
rect 10859 13586 10927 13642
rect 10983 13586 11051 13642
rect 11107 13586 11175 13642
rect 11231 13586 11299 13642
rect 11355 13586 11423 13642
rect 11479 13586 11547 13642
rect 11603 13586 11671 13642
rect 11727 13586 11795 13642
rect 11851 13586 11919 13642
rect 11975 13586 12043 13642
rect 12099 13586 12167 13642
rect 12223 13586 12291 13642
rect 12347 13586 12415 13642
rect 12471 13586 12481 13642
rect 10669 13518 12481 13586
rect 10669 13462 10679 13518
rect 10735 13462 10803 13518
rect 10859 13462 10927 13518
rect 10983 13462 11051 13518
rect 11107 13462 11175 13518
rect 11231 13462 11299 13518
rect 11355 13462 11423 13518
rect 11479 13462 11547 13518
rect 11603 13462 11671 13518
rect 11727 13462 11795 13518
rect 11851 13462 11919 13518
rect 11975 13462 12043 13518
rect 12099 13462 12167 13518
rect 12223 13462 12291 13518
rect 12347 13462 12415 13518
rect 12471 13462 12481 13518
rect 10669 13394 12481 13462
rect 10669 13338 10679 13394
rect 10735 13338 10803 13394
rect 10859 13338 10927 13394
rect 10983 13338 11051 13394
rect 11107 13338 11175 13394
rect 11231 13338 11299 13394
rect 11355 13338 11423 13394
rect 11479 13338 11547 13394
rect 11603 13338 11671 13394
rect 11727 13338 11795 13394
rect 11851 13338 11919 13394
rect 11975 13338 12043 13394
rect 12099 13338 12167 13394
rect 12223 13338 12291 13394
rect 12347 13338 12415 13394
rect 12471 13338 12481 13394
rect 10669 13270 12481 13338
rect 10669 13214 10679 13270
rect 10735 13214 10803 13270
rect 10859 13214 10927 13270
rect 10983 13214 11051 13270
rect 11107 13214 11175 13270
rect 11231 13214 11299 13270
rect 11355 13214 11423 13270
rect 11479 13214 11547 13270
rect 11603 13214 11671 13270
rect 11727 13214 11795 13270
rect 11851 13214 11919 13270
rect 11975 13214 12043 13270
rect 12099 13214 12167 13270
rect 12223 13214 12291 13270
rect 12347 13214 12415 13270
rect 12471 13214 12481 13270
rect 10669 13146 12481 13214
rect 10669 13090 10679 13146
rect 10735 13090 10803 13146
rect 10859 13090 10927 13146
rect 10983 13090 11051 13146
rect 11107 13090 11175 13146
rect 11231 13090 11299 13146
rect 11355 13090 11423 13146
rect 11479 13090 11547 13146
rect 11603 13090 11671 13146
rect 11727 13090 11795 13146
rect 11851 13090 11919 13146
rect 11975 13090 12043 13146
rect 12099 13090 12167 13146
rect 12223 13090 12291 13146
rect 12347 13090 12415 13146
rect 12471 13090 12481 13146
rect 10669 13022 12481 13090
rect 10669 12966 10679 13022
rect 10735 12966 10803 13022
rect 10859 12966 10927 13022
rect 10983 12966 11051 13022
rect 11107 12966 11175 13022
rect 11231 12966 11299 13022
rect 11355 12966 11423 13022
rect 11479 12966 11547 13022
rect 11603 12966 11671 13022
rect 11727 12966 11795 13022
rect 11851 12966 11919 13022
rect 11975 12966 12043 13022
rect 12099 12966 12167 13022
rect 12223 12966 12291 13022
rect 12347 12966 12415 13022
rect 12471 12966 12481 13022
rect 10669 12898 12481 12966
rect 10669 12842 10679 12898
rect 10735 12842 10803 12898
rect 10859 12842 10927 12898
rect 10983 12842 11051 12898
rect 11107 12842 11175 12898
rect 11231 12842 11299 12898
rect 11355 12842 11423 12898
rect 11479 12842 11547 12898
rect 11603 12842 11671 12898
rect 11727 12842 11795 12898
rect 11851 12842 11919 12898
rect 11975 12842 12043 12898
rect 12099 12842 12167 12898
rect 12223 12842 12291 12898
rect 12347 12842 12415 12898
rect 12471 12842 12481 12898
rect 10669 12832 12481 12842
rect 2497 12544 4309 12554
rect 2497 12488 2507 12544
rect 2563 12488 2631 12544
rect 2687 12488 2755 12544
rect 2811 12488 2879 12544
rect 2935 12488 3003 12544
rect 3059 12488 3127 12544
rect 3183 12488 3251 12544
rect 3307 12488 3375 12544
rect 3431 12488 3499 12544
rect 3555 12488 3623 12544
rect 3679 12488 3747 12544
rect 3803 12488 3871 12544
rect 3927 12488 3995 12544
rect 4051 12488 4119 12544
rect 4175 12488 4243 12544
rect 4299 12488 4309 12544
rect 2497 12420 4309 12488
rect 2497 12364 2507 12420
rect 2563 12364 2631 12420
rect 2687 12364 2755 12420
rect 2811 12364 2879 12420
rect 2935 12364 3003 12420
rect 3059 12364 3127 12420
rect 3183 12364 3251 12420
rect 3307 12364 3375 12420
rect 3431 12364 3499 12420
rect 3555 12364 3623 12420
rect 3679 12364 3747 12420
rect 3803 12364 3871 12420
rect 3927 12364 3995 12420
rect 4051 12364 4119 12420
rect 4175 12364 4243 12420
rect 4299 12364 4309 12420
rect 2497 12296 4309 12364
rect 2497 12240 2507 12296
rect 2563 12240 2631 12296
rect 2687 12240 2755 12296
rect 2811 12240 2879 12296
rect 2935 12240 3003 12296
rect 3059 12240 3127 12296
rect 3183 12240 3251 12296
rect 3307 12240 3375 12296
rect 3431 12240 3499 12296
rect 3555 12240 3623 12296
rect 3679 12240 3747 12296
rect 3803 12240 3871 12296
rect 3927 12240 3995 12296
rect 4051 12240 4119 12296
rect 4175 12240 4243 12296
rect 4299 12240 4309 12296
rect 2497 12172 4309 12240
rect 2497 12116 2507 12172
rect 2563 12116 2631 12172
rect 2687 12116 2755 12172
rect 2811 12116 2879 12172
rect 2935 12116 3003 12172
rect 3059 12116 3127 12172
rect 3183 12116 3251 12172
rect 3307 12116 3375 12172
rect 3431 12116 3499 12172
rect 3555 12116 3623 12172
rect 3679 12116 3747 12172
rect 3803 12116 3871 12172
rect 3927 12116 3995 12172
rect 4051 12116 4119 12172
rect 4175 12116 4243 12172
rect 4299 12116 4309 12172
rect 2497 12048 4309 12116
rect 2497 11992 2507 12048
rect 2563 11992 2631 12048
rect 2687 11992 2755 12048
rect 2811 11992 2879 12048
rect 2935 11992 3003 12048
rect 3059 11992 3127 12048
rect 3183 11992 3251 12048
rect 3307 11992 3375 12048
rect 3431 11992 3499 12048
rect 3555 11992 3623 12048
rect 3679 11992 3747 12048
rect 3803 11992 3871 12048
rect 3927 11992 3995 12048
rect 4051 11992 4119 12048
rect 4175 11992 4243 12048
rect 4299 11992 4309 12048
rect 2497 11924 4309 11992
rect 2497 11868 2507 11924
rect 2563 11868 2631 11924
rect 2687 11868 2755 11924
rect 2811 11868 2879 11924
rect 2935 11868 3003 11924
rect 3059 11868 3127 11924
rect 3183 11868 3251 11924
rect 3307 11868 3375 11924
rect 3431 11868 3499 11924
rect 3555 11868 3623 11924
rect 3679 11868 3747 11924
rect 3803 11868 3871 11924
rect 3927 11868 3995 11924
rect 4051 11868 4119 11924
rect 4175 11868 4243 11924
rect 4299 11868 4309 11924
rect 2497 11800 4309 11868
rect 2497 11744 2507 11800
rect 2563 11744 2631 11800
rect 2687 11744 2755 11800
rect 2811 11744 2879 11800
rect 2935 11744 3003 11800
rect 3059 11744 3127 11800
rect 3183 11744 3251 11800
rect 3307 11744 3375 11800
rect 3431 11744 3499 11800
rect 3555 11744 3623 11800
rect 3679 11744 3747 11800
rect 3803 11744 3871 11800
rect 3927 11744 3995 11800
rect 4051 11744 4119 11800
rect 4175 11744 4243 11800
rect 4299 11744 4309 11800
rect 2497 11676 4309 11744
rect 2497 11620 2507 11676
rect 2563 11620 2631 11676
rect 2687 11620 2755 11676
rect 2811 11620 2879 11676
rect 2935 11620 3003 11676
rect 3059 11620 3127 11676
rect 3183 11620 3251 11676
rect 3307 11620 3375 11676
rect 3431 11620 3499 11676
rect 3555 11620 3623 11676
rect 3679 11620 3747 11676
rect 3803 11620 3871 11676
rect 3927 11620 3995 11676
rect 4051 11620 4119 11676
rect 4175 11620 4243 11676
rect 4299 11620 4309 11676
rect 2497 11552 4309 11620
rect 2497 11496 2507 11552
rect 2563 11496 2631 11552
rect 2687 11496 2755 11552
rect 2811 11496 2879 11552
rect 2935 11496 3003 11552
rect 3059 11496 3127 11552
rect 3183 11496 3251 11552
rect 3307 11496 3375 11552
rect 3431 11496 3499 11552
rect 3555 11496 3623 11552
rect 3679 11496 3747 11552
rect 3803 11496 3871 11552
rect 3927 11496 3995 11552
rect 4051 11496 4119 11552
rect 4175 11496 4243 11552
rect 4299 11496 4309 11552
rect 2497 11428 4309 11496
rect 2497 11372 2507 11428
rect 2563 11372 2631 11428
rect 2687 11372 2755 11428
rect 2811 11372 2879 11428
rect 2935 11372 3003 11428
rect 3059 11372 3127 11428
rect 3183 11372 3251 11428
rect 3307 11372 3375 11428
rect 3431 11372 3499 11428
rect 3555 11372 3623 11428
rect 3679 11372 3747 11428
rect 3803 11372 3871 11428
rect 3927 11372 3995 11428
rect 4051 11372 4119 11428
rect 4175 11372 4243 11428
rect 4299 11372 4309 11428
rect 2497 11304 4309 11372
rect 2497 11248 2507 11304
rect 2563 11248 2631 11304
rect 2687 11248 2755 11304
rect 2811 11248 2879 11304
rect 2935 11248 3003 11304
rect 3059 11248 3127 11304
rect 3183 11248 3251 11304
rect 3307 11248 3375 11304
rect 3431 11248 3499 11304
rect 3555 11248 3623 11304
rect 3679 11248 3747 11304
rect 3803 11248 3871 11304
rect 3927 11248 3995 11304
rect 4051 11248 4119 11304
rect 4175 11248 4243 11304
rect 4299 11248 4309 11304
rect 2497 11238 4309 11248
rect 6358 12544 7426 12554
rect 6358 12488 6368 12544
rect 6424 12488 6492 12544
rect 6548 12488 6616 12544
rect 6672 12488 6740 12544
rect 6796 12488 6864 12544
rect 6920 12488 6988 12544
rect 7044 12488 7112 12544
rect 7168 12488 7236 12544
rect 7292 12488 7360 12544
rect 7416 12488 7426 12544
rect 6358 12420 7426 12488
rect 6358 12364 6368 12420
rect 6424 12364 6492 12420
rect 6548 12364 6616 12420
rect 6672 12364 6740 12420
rect 6796 12364 6864 12420
rect 6920 12364 6988 12420
rect 7044 12364 7112 12420
rect 7168 12364 7236 12420
rect 7292 12364 7360 12420
rect 7416 12364 7426 12420
rect 6358 12296 7426 12364
rect 6358 12240 6368 12296
rect 6424 12240 6492 12296
rect 6548 12240 6616 12296
rect 6672 12240 6740 12296
rect 6796 12240 6864 12296
rect 6920 12240 6988 12296
rect 7044 12240 7112 12296
rect 7168 12240 7236 12296
rect 7292 12240 7360 12296
rect 7416 12240 7426 12296
rect 6358 12172 7426 12240
rect 6358 12116 6368 12172
rect 6424 12116 6492 12172
rect 6548 12116 6616 12172
rect 6672 12116 6740 12172
rect 6796 12116 6864 12172
rect 6920 12116 6988 12172
rect 7044 12116 7112 12172
rect 7168 12116 7236 12172
rect 7292 12116 7360 12172
rect 7416 12116 7426 12172
rect 6358 12048 7426 12116
rect 6358 11992 6368 12048
rect 6424 11992 6492 12048
rect 6548 11992 6616 12048
rect 6672 11992 6740 12048
rect 6796 11992 6864 12048
rect 6920 11992 6988 12048
rect 7044 11992 7112 12048
rect 7168 11992 7236 12048
rect 7292 11992 7360 12048
rect 7416 11992 7426 12048
rect 6358 11924 7426 11992
rect 6358 11868 6368 11924
rect 6424 11868 6492 11924
rect 6548 11868 6616 11924
rect 6672 11868 6740 11924
rect 6796 11868 6864 11924
rect 6920 11868 6988 11924
rect 7044 11868 7112 11924
rect 7168 11868 7236 11924
rect 7292 11868 7360 11924
rect 7416 11868 7426 11924
rect 6358 11800 7426 11868
rect 6358 11744 6368 11800
rect 6424 11744 6492 11800
rect 6548 11744 6616 11800
rect 6672 11744 6740 11800
rect 6796 11744 6864 11800
rect 6920 11744 6988 11800
rect 7044 11744 7112 11800
rect 7168 11744 7236 11800
rect 7292 11744 7360 11800
rect 7416 11744 7426 11800
rect 6358 11676 7426 11744
rect 6358 11620 6368 11676
rect 6424 11620 6492 11676
rect 6548 11620 6616 11676
rect 6672 11620 6740 11676
rect 6796 11620 6864 11676
rect 6920 11620 6988 11676
rect 7044 11620 7112 11676
rect 7168 11620 7236 11676
rect 7292 11620 7360 11676
rect 7416 11620 7426 11676
rect 6358 11552 7426 11620
rect 6358 11496 6368 11552
rect 6424 11496 6492 11552
rect 6548 11496 6616 11552
rect 6672 11496 6740 11552
rect 6796 11496 6864 11552
rect 6920 11496 6988 11552
rect 7044 11496 7112 11552
rect 7168 11496 7236 11552
rect 7292 11496 7360 11552
rect 7416 11496 7426 11552
rect 6358 11428 7426 11496
rect 6358 11372 6368 11428
rect 6424 11372 6492 11428
rect 6548 11372 6616 11428
rect 6672 11372 6740 11428
rect 6796 11372 6864 11428
rect 6920 11372 6988 11428
rect 7044 11372 7112 11428
rect 7168 11372 7236 11428
rect 7292 11372 7360 11428
rect 7416 11372 7426 11428
rect 6358 11304 7426 11372
rect 6358 11248 6368 11304
rect 6424 11248 6492 11304
rect 6548 11248 6616 11304
rect 6672 11248 6740 11304
rect 6796 11248 6864 11304
rect 6920 11248 6988 11304
rect 7044 11248 7112 11304
rect 7168 11248 7236 11304
rect 7292 11248 7360 11304
rect 7416 11248 7426 11304
rect 6358 11238 7426 11248
rect 8741 12544 10553 12554
rect 8741 12488 8751 12544
rect 8807 12488 8875 12544
rect 8931 12488 8999 12544
rect 9055 12488 9123 12544
rect 9179 12488 9247 12544
rect 9303 12488 9371 12544
rect 9427 12488 9495 12544
rect 9551 12488 9619 12544
rect 9675 12488 9743 12544
rect 9799 12488 9867 12544
rect 9923 12488 9991 12544
rect 10047 12488 10115 12544
rect 10171 12488 10239 12544
rect 10295 12488 10363 12544
rect 10419 12488 10487 12544
rect 10543 12488 10553 12544
rect 8741 12420 10553 12488
rect 8741 12364 8751 12420
rect 8807 12364 8875 12420
rect 8931 12364 8999 12420
rect 9055 12364 9123 12420
rect 9179 12364 9247 12420
rect 9303 12364 9371 12420
rect 9427 12364 9495 12420
rect 9551 12364 9619 12420
rect 9675 12364 9743 12420
rect 9799 12364 9867 12420
rect 9923 12364 9991 12420
rect 10047 12364 10115 12420
rect 10171 12364 10239 12420
rect 10295 12364 10363 12420
rect 10419 12364 10487 12420
rect 10543 12364 10553 12420
rect 8741 12296 10553 12364
rect 8741 12240 8751 12296
rect 8807 12240 8875 12296
rect 8931 12240 8999 12296
rect 9055 12240 9123 12296
rect 9179 12240 9247 12296
rect 9303 12240 9371 12296
rect 9427 12240 9495 12296
rect 9551 12240 9619 12296
rect 9675 12240 9743 12296
rect 9799 12240 9867 12296
rect 9923 12240 9991 12296
rect 10047 12240 10115 12296
rect 10171 12240 10239 12296
rect 10295 12240 10363 12296
rect 10419 12240 10487 12296
rect 10543 12240 10553 12296
rect 8741 12172 10553 12240
rect 8741 12116 8751 12172
rect 8807 12116 8875 12172
rect 8931 12116 8999 12172
rect 9055 12116 9123 12172
rect 9179 12116 9247 12172
rect 9303 12116 9371 12172
rect 9427 12116 9495 12172
rect 9551 12116 9619 12172
rect 9675 12116 9743 12172
rect 9799 12116 9867 12172
rect 9923 12116 9991 12172
rect 10047 12116 10115 12172
rect 10171 12116 10239 12172
rect 10295 12116 10363 12172
rect 10419 12116 10487 12172
rect 10543 12116 10553 12172
rect 8741 12048 10553 12116
rect 8741 11992 8751 12048
rect 8807 11992 8875 12048
rect 8931 11992 8999 12048
rect 9055 11992 9123 12048
rect 9179 11992 9247 12048
rect 9303 11992 9371 12048
rect 9427 11992 9495 12048
rect 9551 11992 9619 12048
rect 9675 11992 9743 12048
rect 9799 11992 9867 12048
rect 9923 11992 9991 12048
rect 10047 11992 10115 12048
rect 10171 11992 10239 12048
rect 10295 11992 10363 12048
rect 10419 11992 10487 12048
rect 10543 11992 10553 12048
rect 8741 11924 10553 11992
rect 8741 11868 8751 11924
rect 8807 11868 8875 11924
rect 8931 11868 8999 11924
rect 9055 11868 9123 11924
rect 9179 11868 9247 11924
rect 9303 11868 9371 11924
rect 9427 11868 9495 11924
rect 9551 11868 9619 11924
rect 9675 11868 9743 11924
rect 9799 11868 9867 11924
rect 9923 11868 9991 11924
rect 10047 11868 10115 11924
rect 10171 11868 10239 11924
rect 10295 11868 10363 11924
rect 10419 11868 10487 11924
rect 10543 11868 10553 11924
rect 8741 11800 10553 11868
rect 8741 11744 8751 11800
rect 8807 11744 8875 11800
rect 8931 11744 8999 11800
rect 9055 11744 9123 11800
rect 9179 11744 9247 11800
rect 9303 11744 9371 11800
rect 9427 11744 9495 11800
rect 9551 11744 9619 11800
rect 9675 11744 9743 11800
rect 9799 11744 9867 11800
rect 9923 11744 9991 11800
rect 10047 11744 10115 11800
rect 10171 11744 10239 11800
rect 10295 11744 10363 11800
rect 10419 11744 10487 11800
rect 10543 11744 10553 11800
rect 8741 11676 10553 11744
rect 8741 11620 8751 11676
rect 8807 11620 8875 11676
rect 8931 11620 8999 11676
rect 9055 11620 9123 11676
rect 9179 11620 9247 11676
rect 9303 11620 9371 11676
rect 9427 11620 9495 11676
rect 9551 11620 9619 11676
rect 9675 11620 9743 11676
rect 9799 11620 9867 11676
rect 9923 11620 9991 11676
rect 10047 11620 10115 11676
rect 10171 11620 10239 11676
rect 10295 11620 10363 11676
rect 10419 11620 10487 11676
rect 10543 11620 10553 11676
rect 8741 11552 10553 11620
rect 8741 11496 8751 11552
rect 8807 11496 8875 11552
rect 8931 11496 8999 11552
rect 9055 11496 9123 11552
rect 9179 11496 9247 11552
rect 9303 11496 9371 11552
rect 9427 11496 9495 11552
rect 9551 11496 9619 11552
rect 9675 11496 9743 11552
rect 9799 11496 9867 11552
rect 9923 11496 9991 11552
rect 10047 11496 10115 11552
rect 10171 11496 10239 11552
rect 10295 11496 10363 11552
rect 10419 11496 10487 11552
rect 10543 11496 10553 11552
rect 8741 11428 10553 11496
rect 8741 11372 8751 11428
rect 8807 11372 8875 11428
rect 8931 11372 8999 11428
rect 9055 11372 9123 11428
rect 9179 11372 9247 11428
rect 9303 11372 9371 11428
rect 9427 11372 9495 11428
rect 9551 11372 9619 11428
rect 9675 11372 9743 11428
rect 9799 11372 9867 11428
rect 9923 11372 9991 11428
rect 10047 11372 10115 11428
rect 10171 11372 10239 11428
rect 10295 11372 10363 11428
rect 10419 11372 10487 11428
rect 10543 11372 10553 11428
rect 8741 11304 10553 11372
rect 8741 11248 8751 11304
rect 8807 11248 8875 11304
rect 8931 11248 8999 11304
rect 9055 11248 9123 11304
rect 9179 11248 9247 11304
rect 9303 11248 9371 11304
rect 9427 11248 9495 11304
rect 9551 11248 9619 11304
rect 9675 11248 9743 11304
rect 9799 11248 9867 11304
rect 9923 11248 9991 11304
rect 10047 11248 10115 11304
rect 10171 11248 10239 11304
rect 10295 11248 10363 11304
rect 10419 11248 10487 11304
rect 10543 11248 10553 11304
rect 8741 11238 10553 11248
rect 12842 12544 13910 12554
rect 12842 12488 12852 12544
rect 12908 12488 12976 12544
rect 13032 12488 13100 12544
rect 13156 12488 13224 12544
rect 13280 12488 13348 12544
rect 13404 12488 13472 12544
rect 13528 12488 13596 12544
rect 13652 12488 13720 12544
rect 13776 12488 13844 12544
rect 13900 12488 13910 12544
rect 12842 12420 13910 12488
rect 12842 12364 12852 12420
rect 12908 12364 12976 12420
rect 13032 12364 13100 12420
rect 13156 12364 13224 12420
rect 13280 12364 13348 12420
rect 13404 12364 13472 12420
rect 13528 12364 13596 12420
rect 13652 12364 13720 12420
rect 13776 12364 13844 12420
rect 13900 12364 13910 12420
rect 12842 12296 13910 12364
rect 12842 12240 12852 12296
rect 12908 12240 12976 12296
rect 13032 12240 13100 12296
rect 13156 12240 13224 12296
rect 13280 12240 13348 12296
rect 13404 12240 13472 12296
rect 13528 12240 13596 12296
rect 13652 12240 13720 12296
rect 13776 12240 13844 12296
rect 13900 12240 13910 12296
rect 12842 12172 13910 12240
rect 12842 12116 12852 12172
rect 12908 12116 12976 12172
rect 13032 12116 13100 12172
rect 13156 12116 13224 12172
rect 13280 12116 13348 12172
rect 13404 12116 13472 12172
rect 13528 12116 13596 12172
rect 13652 12116 13720 12172
rect 13776 12116 13844 12172
rect 13900 12116 13910 12172
rect 12842 12048 13910 12116
rect 12842 11992 12852 12048
rect 12908 11992 12976 12048
rect 13032 11992 13100 12048
rect 13156 11992 13224 12048
rect 13280 11992 13348 12048
rect 13404 11992 13472 12048
rect 13528 11992 13596 12048
rect 13652 11992 13720 12048
rect 13776 11992 13844 12048
rect 13900 11992 13910 12048
rect 12842 11924 13910 11992
rect 12842 11868 12852 11924
rect 12908 11868 12976 11924
rect 13032 11868 13100 11924
rect 13156 11868 13224 11924
rect 13280 11868 13348 11924
rect 13404 11868 13472 11924
rect 13528 11868 13596 11924
rect 13652 11868 13720 11924
rect 13776 11868 13844 11924
rect 13900 11868 13910 11924
rect 12842 11800 13910 11868
rect 12842 11744 12852 11800
rect 12908 11744 12976 11800
rect 13032 11744 13100 11800
rect 13156 11744 13224 11800
rect 13280 11744 13348 11800
rect 13404 11744 13472 11800
rect 13528 11744 13596 11800
rect 13652 11744 13720 11800
rect 13776 11744 13844 11800
rect 13900 11744 13910 11800
rect 12842 11676 13910 11744
rect 12842 11620 12852 11676
rect 12908 11620 12976 11676
rect 13032 11620 13100 11676
rect 13156 11620 13224 11676
rect 13280 11620 13348 11676
rect 13404 11620 13472 11676
rect 13528 11620 13596 11676
rect 13652 11620 13720 11676
rect 13776 11620 13844 11676
rect 13900 11620 13910 11676
rect 12842 11552 13910 11620
rect 12842 11496 12852 11552
rect 12908 11496 12976 11552
rect 13032 11496 13100 11552
rect 13156 11496 13224 11552
rect 13280 11496 13348 11552
rect 13404 11496 13472 11552
rect 13528 11496 13596 11552
rect 13652 11496 13720 11552
rect 13776 11496 13844 11552
rect 13900 11496 13910 11552
rect 12842 11428 13910 11496
rect 12842 11372 12852 11428
rect 12908 11372 12976 11428
rect 13032 11372 13100 11428
rect 13156 11372 13224 11428
rect 13280 11372 13348 11428
rect 13404 11372 13472 11428
rect 13528 11372 13596 11428
rect 13652 11372 13720 11428
rect 13776 11372 13844 11428
rect 13900 11372 13910 11428
rect 12842 11304 13910 11372
rect 12842 11248 12852 11304
rect 12908 11248 12976 11304
rect 13032 11248 13100 11304
rect 13156 11248 13224 11304
rect 13280 11248 13348 11304
rect 13404 11248 13472 11304
rect 13528 11248 13596 11304
rect 13652 11248 13720 11304
rect 13776 11248 13844 11304
rect 13900 11248 13910 11304
rect 12842 11238 13910 11248
rect 1068 10944 2136 10954
rect 1068 10888 1078 10944
rect 1134 10888 1202 10944
rect 1258 10888 1326 10944
rect 1382 10888 1450 10944
rect 1506 10888 1574 10944
rect 1630 10888 1698 10944
rect 1754 10888 1822 10944
rect 1878 10888 1946 10944
rect 2002 10888 2070 10944
rect 2126 10888 2136 10944
rect 1068 10820 2136 10888
rect 1068 10764 1078 10820
rect 1134 10764 1202 10820
rect 1258 10764 1326 10820
rect 1382 10764 1450 10820
rect 1506 10764 1574 10820
rect 1630 10764 1698 10820
rect 1754 10764 1822 10820
rect 1878 10764 1946 10820
rect 2002 10764 2070 10820
rect 2126 10764 2136 10820
rect 1068 10696 2136 10764
rect 1068 10640 1078 10696
rect 1134 10640 1202 10696
rect 1258 10640 1326 10696
rect 1382 10640 1450 10696
rect 1506 10640 1574 10696
rect 1630 10640 1698 10696
rect 1754 10640 1822 10696
rect 1878 10640 1946 10696
rect 2002 10640 2070 10696
rect 2126 10640 2136 10696
rect 1068 10572 2136 10640
rect 1068 10516 1078 10572
rect 1134 10516 1202 10572
rect 1258 10516 1326 10572
rect 1382 10516 1450 10572
rect 1506 10516 1574 10572
rect 1630 10516 1698 10572
rect 1754 10516 1822 10572
rect 1878 10516 1946 10572
rect 2002 10516 2070 10572
rect 2126 10516 2136 10572
rect 1068 10448 2136 10516
rect 1068 10392 1078 10448
rect 1134 10392 1202 10448
rect 1258 10392 1326 10448
rect 1382 10392 1450 10448
rect 1506 10392 1574 10448
rect 1630 10392 1698 10448
rect 1754 10392 1822 10448
rect 1878 10392 1946 10448
rect 2002 10392 2070 10448
rect 2126 10392 2136 10448
rect 1068 10324 2136 10392
rect 1068 10268 1078 10324
rect 1134 10268 1202 10324
rect 1258 10268 1326 10324
rect 1382 10268 1450 10324
rect 1506 10268 1574 10324
rect 1630 10268 1698 10324
rect 1754 10268 1822 10324
rect 1878 10268 1946 10324
rect 2002 10268 2070 10324
rect 2126 10268 2136 10324
rect 1068 10200 2136 10268
rect 1068 10144 1078 10200
rect 1134 10144 1202 10200
rect 1258 10144 1326 10200
rect 1382 10144 1450 10200
rect 1506 10144 1574 10200
rect 1630 10144 1698 10200
rect 1754 10144 1822 10200
rect 1878 10144 1946 10200
rect 2002 10144 2070 10200
rect 2126 10144 2136 10200
rect 1068 10076 2136 10144
rect 1068 10020 1078 10076
rect 1134 10020 1202 10076
rect 1258 10020 1326 10076
rect 1382 10020 1450 10076
rect 1506 10020 1574 10076
rect 1630 10020 1698 10076
rect 1754 10020 1822 10076
rect 1878 10020 1946 10076
rect 2002 10020 2070 10076
rect 2126 10020 2136 10076
rect 1068 9952 2136 10020
rect 1068 9896 1078 9952
rect 1134 9896 1202 9952
rect 1258 9896 1326 9952
rect 1382 9896 1450 9952
rect 1506 9896 1574 9952
rect 1630 9896 1698 9952
rect 1754 9896 1822 9952
rect 1878 9896 1946 9952
rect 2002 9896 2070 9952
rect 2126 9896 2136 9952
rect 1068 9828 2136 9896
rect 1068 9772 1078 9828
rect 1134 9772 1202 9828
rect 1258 9772 1326 9828
rect 1382 9772 1450 9828
rect 1506 9772 1574 9828
rect 1630 9772 1698 9828
rect 1754 9772 1822 9828
rect 1878 9772 1946 9828
rect 2002 9772 2070 9828
rect 2126 9772 2136 9828
rect 1068 9704 2136 9772
rect 1068 9648 1078 9704
rect 1134 9648 1202 9704
rect 1258 9648 1326 9704
rect 1382 9648 1450 9704
rect 1506 9648 1574 9704
rect 1630 9648 1698 9704
rect 1754 9648 1822 9704
rect 1878 9648 1946 9704
rect 2002 9648 2070 9704
rect 2126 9648 2136 9704
rect 1068 9638 2136 9648
rect 4425 10944 6237 10954
rect 4425 10888 4435 10944
rect 4491 10888 4559 10944
rect 4615 10888 4683 10944
rect 4739 10888 4807 10944
rect 4863 10888 4931 10944
rect 4987 10888 5055 10944
rect 5111 10888 5179 10944
rect 5235 10888 5303 10944
rect 5359 10888 5427 10944
rect 5483 10888 5551 10944
rect 5607 10888 5675 10944
rect 5731 10888 5799 10944
rect 5855 10888 5923 10944
rect 5979 10888 6047 10944
rect 6103 10888 6171 10944
rect 6227 10888 6237 10944
rect 4425 10820 6237 10888
rect 4425 10764 4435 10820
rect 4491 10764 4559 10820
rect 4615 10764 4683 10820
rect 4739 10764 4807 10820
rect 4863 10764 4931 10820
rect 4987 10764 5055 10820
rect 5111 10764 5179 10820
rect 5235 10764 5303 10820
rect 5359 10764 5427 10820
rect 5483 10764 5551 10820
rect 5607 10764 5675 10820
rect 5731 10764 5799 10820
rect 5855 10764 5923 10820
rect 5979 10764 6047 10820
rect 6103 10764 6171 10820
rect 6227 10764 6237 10820
rect 4425 10696 6237 10764
rect 4425 10640 4435 10696
rect 4491 10640 4559 10696
rect 4615 10640 4683 10696
rect 4739 10640 4807 10696
rect 4863 10640 4931 10696
rect 4987 10640 5055 10696
rect 5111 10640 5179 10696
rect 5235 10640 5303 10696
rect 5359 10640 5427 10696
rect 5483 10640 5551 10696
rect 5607 10640 5675 10696
rect 5731 10640 5799 10696
rect 5855 10640 5923 10696
rect 5979 10640 6047 10696
rect 6103 10640 6171 10696
rect 6227 10640 6237 10696
rect 4425 10572 6237 10640
rect 4425 10516 4435 10572
rect 4491 10516 4559 10572
rect 4615 10516 4683 10572
rect 4739 10516 4807 10572
rect 4863 10516 4931 10572
rect 4987 10516 5055 10572
rect 5111 10516 5179 10572
rect 5235 10516 5303 10572
rect 5359 10516 5427 10572
rect 5483 10516 5551 10572
rect 5607 10516 5675 10572
rect 5731 10516 5799 10572
rect 5855 10516 5923 10572
rect 5979 10516 6047 10572
rect 6103 10516 6171 10572
rect 6227 10516 6237 10572
rect 4425 10448 6237 10516
rect 4425 10392 4435 10448
rect 4491 10392 4559 10448
rect 4615 10392 4683 10448
rect 4739 10392 4807 10448
rect 4863 10392 4931 10448
rect 4987 10392 5055 10448
rect 5111 10392 5179 10448
rect 5235 10392 5303 10448
rect 5359 10392 5427 10448
rect 5483 10392 5551 10448
rect 5607 10392 5675 10448
rect 5731 10392 5799 10448
rect 5855 10392 5923 10448
rect 5979 10392 6047 10448
rect 6103 10392 6171 10448
rect 6227 10392 6237 10448
rect 4425 10324 6237 10392
rect 4425 10268 4435 10324
rect 4491 10268 4559 10324
rect 4615 10268 4683 10324
rect 4739 10268 4807 10324
rect 4863 10268 4931 10324
rect 4987 10268 5055 10324
rect 5111 10268 5179 10324
rect 5235 10268 5303 10324
rect 5359 10268 5427 10324
rect 5483 10268 5551 10324
rect 5607 10268 5675 10324
rect 5731 10268 5799 10324
rect 5855 10268 5923 10324
rect 5979 10268 6047 10324
rect 6103 10268 6171 10324
rect 6227 10268 6237 10324
rect 4425 10200 6237 10268
rect 4425 10144 4435 10200
rect 4491 10144 4559 10200
rect 4615 10144 4683 10200
rect 4739 10144 4807 10200
rect 4863 10144 4931 10200
rect 4987 10144 5055 10200
rect 5111 10144 5179 10200
rect 5235 10144 5303 10200
rect 5359 10144 5427 10200
rect 5483 10144 5551 10200
rect 5607 10144 5675 10200
rect 5731 10144 5799 10200
rect 5855 10144 5923 10200
rect 5979 10144 6047 10200
rect 6103 10144 6171 10200
rect 6227 10144 6237 10200
rect 4425 10076 6237 10144
rect 4425 10020 4435 10076
rect 4491 10020 4559 10076
rect 4615 10020 4683 10076
rect 4739 10020 4807 10076
rect 4863 10020 4931 10076
rect 4987 10020 5055 10076
rect 5111 10020 5179 10076
rect 5235 10020 5303 10076
rect 5359 10020 5427 10076
rect 5483 10020 5551 10076
rect 5607 10020 5675 10076
rect 5731 10020 5799 10076
rect 5855 10020 5923 10076
rect 5979 10020 6047 10076
rect 6103 10020 6171 10076
rect 6227 10020 6237 10076
rect 4425 9952 6237 10020
rect 4425 9896 4435 9952
rect 4491 9896 4559 9952
rect 4615 9896 4683 9952
rect 4739 9896 4807 9952
rect 4863 9896 4931 9952
rect 4987 9896 5055 9952
rect 5111 9896 5179 9952
rect 5235 9896 5303 9952
rect 5359 9896 5427 9952
rect 5483 9896 5551 9952
rect 5607 9896 5675 9952
rect 5731 9896 5799 9952
rect 5855 9896 5923 9952
rect 5979 9896 6047 9952
rect 6103 9896 6171 9952
rect 6227 9896 6237 9952
rect 4425 9828 6237 9896
rect 4425 9772 4435 9828
rect 4491 9772 4559 9828
rect 4615 9772 4683 9828
rect 4739 9772 4807 9828
rect 4863 9772 4931 9828
rect 4987 9772 5055 9828
rect 5111 9772 5179 9828
rect 5235 9772 5303 9828
rect 5359 9772 5427 9828
rect 5483 9772 5551 9828
rect 5607 9772 5675 9828
rect 5731 9772 5799 9828
rect 5855 9772 5923 9828
rect 5979 9772 6047 9828
rect 6103 9772 6171 9828
rect 6227 9772 6237 9828
rect 4425 9704 6237 9772
rect 4425 9648 4435 9704
rect 4491 9648 4559 9704
rect 4615 9648 4683 9704
rect 4739 9648 4807 9704
rect 4863 9648 4931 9704
rect 4987 9648 5055 9704
rect 5111 9648 5179 9704
rect 5235 9648 5303 9704
rect 5359 9648 5427 9704
rect 5483 9648 5551 9704
rect 5607 9648 5675 9704
rect 5731 9648 5799 9704
rect 5855 9648 5923 9704
rect 5979 9648 6047 9704
rect 6103 9648 6171 9704
rect 6227 9648 6237 9704
rect 4425 9638 6237 9648
rect 7552 10944 8620 10954
rect 7552 10888 7562 10944
rect 7618 10888 7686 10944
rect 7742 10888 7810 10944
rect 7866 10888 7934 10944
rect 7990 10888 8058 10944
rect 8114 10888 8182 10944
rect 8238 10888 8306 10944
rect 8362 10888 8430 10944
rect 8486 10888 8554 10944
rect 8610 10888 8620 10944
rect 7552 10820 8620 10888
rect 7552 10764 7562 10820
rect 7618 10764 7686 10820
rect 7742 10764 7810 10820
rect 7866 10764 7934 10820
rect 7990 10764 8058 10820
rect 8114 10764 8182 10820
rect 8238 10764 8306 10820
rect 8362 10764 8430 10820
rect 8486 10764 8554 10820
rect 8610 10764 8620 10820
rect 7552 10696 8620 10764
rect 7552 10640 7562 10696
rect 7618 10640 7686 10696
rect 7742 10640 7810 10696
rect 7866 10640 7934 10696
rect 7990 10640 8058 10696
rect 8114 10640 8182 10696
rect 8238 10640 8306 10696
rect 8362 10640 8430 10696
rect 8486 10640 8554 10696
rect 8610 10640 8620 10696
rect 7552 10572 8620 10640
rect 7552 10516 7562 10572
rect 7618 10516 7686 10572
rect 7742 10516 7810 10572
rect 7866 10516 7934 10572
rect 7990 10516 8058 10572
rect 8114 10516 8182 10572
rect 8238 10516 8306 10572
rect 8362 10516 8430 10572
rect 8486 10516 8554 10572
rect 8610 10516 8620 10572
rect 7552 10448 8620 10516
rect 7552 10392 7562 10448
rect 7618 10392 7686 10448
rect 7742 10392 7810 10448
rect 7866 10392 7934 10448
rect 7990 10392 8058 10448
rect 8114 10392 8182 10448
rect 8238 10392 8306 10448
rect 8362 10392 8430 10448
rect 8486 10392 8554 10448
rect 8610 10392 8620 10448
rect 7552 10324 8620 10392
rect 7552 10268 7562 10324
rect 7618 10268 7686 10324
rect 7742 10268 7810 10324
rect 7866 10268 7934 10324
rect 7990 10268 8058 10324
rect 8114 10268 8182 10324
rect 8238 10268 8306 10324
rect 8362 10268 8430 10324
rect 8486 10268 8554 10324
rect 8610 10268 8620 10324
rect 7552 10200 8620 10268
rect 7552 10144 7562 10200
rect 7618 10144 7686 10200
rect 7742 10144 7810 10200
rect 7866 10144 7934 10200
rect 7990 10144 8058 10200
rect 8114 10144 8182 10200
rect 8238 10144 8306 10200
rect 8362 10144 8430 10200
rect 8486 10144 8554 10200
rect 8610 10144 8620 10200
rect 7552 10076 8620 10144
rect 7552 10020 7562 10076
rect 7618 10020 7686 10076
rect 7742 10020 7810 10076
rect 7866 10020 7934 10076
rect 7990 10020 8058 10076
rect 8114 10020 8182 10076
rect 8238 10020 8306 10076
rect 8362 10020 8430 10076
rect 8486 10020 8554 10076
rect 8610 10020 8620 10076
rect 7552 9952 8620 10020
rect 7552 9896 7562 9952
rect 7618 9896 7686 9952
rect 7742 9896 7810 9952
rect 7866 9896 7934 9952
rect 7990 9896 8058 9952
rect 8114 9896 8182 9952
rect 8238 9896 8306 9952
rect 8362 9896 8430 9952
rect 8486 9896 8554 9952
rect 8610 9896 8620 9952
rect 7552 9828 8620 9896
rect 7552 9772 7562 9828
rect 7618 9772 7686 9828
rect 7742 9772 7810 9828
rect 7866 9772 7934 9828
rect 7990 9772 8058 9828
rect 8114 9772 8182 9828
rect 8238 9772 8306 9828
rect 8362 9772 8430 9828
rect 8486 9772 8554 9828
rect 8610 9772 8620 9828
rect 7552 9704 8620 9772
rect 7552 9648 7562 9704
rect 7618 9648 7686 9704
rect 7742 9648 7810 9704
rect 7866 9648 7934 9704
rect 7990 9648 8058 9704
rect 8114 9648 8182 9704
rect 8238 9648 8306 9704
rect 8362 9648 8430 9704
rect 8486 9648 8554 9704
rect 8610 9648 8620 9704
rect 7552 9638 8620 9648
rect 10669 10944 12481 10954
rect 10669 10888 10679 10944
rect 10735 10888 10803 10944
rect 10859 10888 10927 10944
rect 10983 10888 11051 10944
rect 11107 10888 11175 10944
rect 11231 10888 11299 10944
rect 11355 10888 11423 10944
rect 11479 10888 11547 10944
rect 11603 10888 11671 10944
rect 11727 10888 11795 10944
rect 11851 10888 11919 10944
rect 11975 10888 12043 10944
rect 12099 10888 12167 10944
rect 12223 10888 12291 10944
rect 12347 10888 12415 10944
rect 12471 10888 12481 10944
rect 10669 10820 12481 10888
rect 10669 10764 10679 10820
rect 10735 10764 10803 10820
rect 10859 10764 10927 10820
rect 10983 10764 11051 10820
rect 11107 10764 11175 10820
rect 11231 10764 11299 10820
rect 11355 10764 11423 10820
rect 11479 10764 11547 10820
rect 11603 10764 11671 10820
rect 11727 10764 11795 10820
rect 11851 10764 11919 10820
rect 11975 10764 12043 10820
rect 12099 10764 12167 10820
rect 12223 10764 12291 10820
rect 12347 10764 12415 10820
rect 12471 10764 12481 10820
rect 10669 10696 12481 10764
rect 10669 10640 10679 10696
rect 10735 10640 10803 10696
rect 10859 10640 10927 10696
rect 10983 10640 11051 10696
rect 11107 10640 11175 10696
rect 11231 10640 11299 10696
rect 11355 10640 11423 10696
rect 11479 10640 11547 10696
rect 11603 10640 11671 10696
rect 11727 10640 11795 10696
rect 11851 10640 11919 10696
rect 11975 10640 12043 10696
rect 12099 10640 12167 10696
rect 12223 10640 12291 10696
rect 12347 10640 12415 10696
rect 12471 10640 12481 10696
rect 10669 10572 12481 10640
rect 10669 10516 10679 10572
rect 10735 10516 10803 10572
rect 10859 10516 10927 10572
rect 10983 10516 11051 10572
rect 11107 10516 11175 10572
rect 11231 10516 11299 10572
rect 11355 10516 11423 10572
rect 11479 10516 11547 10572
rect 11603 10516 11671 10572
rect 11727 10516 11795 10572
rect 11851 10516 11919 10572
rect 11975 10516 12043 10572
rect 12099 10516 12167 10572
rect 12223 10516 12291 10572
rect 12347 10516 12415 10572
rect 12471 10516 12481 10572
rect 10669 10448 12481 10516
rect 10669 10392 10679 10448
rect 10735 10392 10803 10448
rect 10859 10392 10927 10448
rect 10983 10392 11051 10448
rect 11107 10392 11175 10448
rect 11231 10392 11299 10448
rect 11355 10392 11423 10448
rect 11479 10392 11547 10448
rect 11603 10392 11671 10448
rect 11727 10392 11795 10448
rect 11851 10392 11919 10448
rect 11975 10392 12043 10448
rect 12099 10392 12167 10448
rect 12223 10392 12291 10448
rect 12347 10392 12415 10448
rect 12471 10392 12481 10448
rect 10669 10324 12481 10392
rect 10669 10268 10679 10324
rect 10735 10268 10803 10324
rect 10859 10268 10927 10324
rect 10983 10268 11051 10324
rect 11107 10268 11175 10324
rect 11231 10268 11299 10324
rect 11355 10268 11423 10324
rect 11479 10268 11547 10324
rect 11603 10268 11671 10324
rect 11727 10268 11795 10324
rect 11851 10268 11919 10324
rect 11975 10268 12043 10324
rect 12099 10268 12167 10324
rect 12223 10268 12291 10324
rect 12347 10268 12415 10324
rect 12471 10268 12481 10324
rect 10669 10200 12481 10268
rect 10669 10144 10679 10200
rect 10735 10144 10803 10200
rect 10859 10144 10927 10200
rect 10983 10144 11051 10200
rect 11107 10144 11175 10200
rect 11231 10144 11299 10200
rect 11355 10144 11423 10200
rect 11479 10144 11547 10200
rect 11603 10144 11671 10200
rect 11727 10144 11795 10200
rect 11851 10144 11919 10200
rect 11975 10144 12043 10200
rect 12099 10144 12167 10200
rect 12223 10144 12291 10200
rect 12347 10144 12415 10200
rect 12471 10144 12481 10200
rect 10669 10076 12481 10144
rect 10669 10020 10679 10076
rect 10735 10020 10803 10076
rect 10859 10020 10927 10076
rect 10983 10020 11051 10076
rect 11107 10020 11175 10076
rect 11231 10020 11299 10076
rect 11355 10020 11423 10076
rect 11479 10020 11547 10076
rect 11603 10020 11671 10076
rect 11727 10020 11795 10076
rect 11851 10020 11919 10076
rect 11975 10020 12043 10076
rect 12099 10020 12167 10076
rect 12223 10020 12291 10076
rect 12347 10020 12415 10076
rect 12471 10020 12481 10076
rect 10669 9952 12481 10020
rect 10669 9896 10679 9952
rect 10735 9896 10803 9952
rect 10859 9896 10927 9952
rect 10983 9896 11051 9952
rect 11107 9896 11175 9952
rect 11231 9896 11299 9952
rect 11355 9896 11423 9952
rect 11479 9896 11547 9952
rect 11603 9896 11671 9952
rect 11727 9896 11795 9952
rect 11851 9896 11919 9952
rect 11975 9896 12043 9952
rect 12099 9896 12167 9952
rect 12223 9896 12291 9952
rect 12347 9896 12415 9952
rect 12471 9896 12481 9952
rect 10669 9828 12481 9896
rect 10669 9772 10679 9828
rect 10735 9772 10803 9828
rect 10859 9772 10927 9828
rect 10983 9772 11051 9828
rect 11107 9772 11175 9828
rect 11231 9772 11299 9828
rect 11355 9772 11423 9828
rect 11479 9772 11547 9828
rect 11603 9772 11671 9828
rect 11727 9772 11795 9828
rect 11851 9772 11919 9828
rect 11975 9772 12043 9828
rect 12099 9772 12167 9828
rect 12223 9772 12291 9828
rect 12347 9772 12415 9828
rect 12471 9772 12481 9828
rect 10669 9704 12481 9772
rect 10669 9648 10679 9704
rect 10735 9648 10803 9704
rect 10859 9648 10927 9704
rect 10983 9648 11051 9704
rect 11107 9648 11175 9704
rect 11231 9648 11299 9704
rect 11355 9648 11423 9704
rect 11479 9648 11547 9704
rect 11603 9648 11671 9704
rect 11727 9648 11795 9704
rect 11851 9648 11919 9704
rect 11975 9648 12043 9704
rect 12099 9648 12167 9704
rect 12223 9648 12291 9704
rect 12347 9648 12415 9704
rect 12471 9648 12481 9704
rect 10669 9638 12481 9648
rect 2497 9350 4309 9360
rect 2497 9294 2507 9350
rect 2563 9294 2631 9350
rect 2687 9294 2755 9350
rect 2811 9294 2879 9350
rect 2935 9294 3003 9350
rect 3059 9294 3127 9350
rect 3183 9294 3251 9350
rect 3307 9294 3375 9350
rect 3431 9294 3499 9350
rect 3555 9294 3623 9350
rect 3679 9294 3747 9350
rect 3803 9294 3871 9350
rect 3927 9294 3995 9350
rect 4051 9294 4119 9350
rect 4175 9294 4243 9350
rect 4299 9294 4309 9350
rect 2497 9226 4309 9294
rect 2497 9170 2507 9226
rect 2563 9170 2631 9226
rect 2687 9170 2755 9226
rect 2811 9170 2879 9226
rect 2935 9170 3003 9226
rect 3059 9170 3127 9226
rect 3183 9170 3251 9226
rect 3307 9170 3375 9226
rect 3431 9170 3499 9226
rect 3555 9170 3623 9226
rect 3679 9170 3747 9226
rect 3803 9170 3871 9226
rect 3927 9170 3995 9226
rect 4051 9170 4119 9226
rect 4175 9170 4243 9226
rect 4299 9170 4309 9226
rect 2497 9102 4309 9170
rect 2497 9046 2507 9102
rect 2563 9046 2631 9102
rect 2687 9046 2755 9102
rect 2811 9046 2879 9102
rect 2935 9046 3003 9102
rect 3059 9046 3127 9102
rect 3183 9046 3251 9102
rect 3307 9046 3375 9102
rect 3431 9046 3499 9102
rect 3555 9046 3623 9102
rect 3679 9046 3747 9102
rect 3803 9046 3871 9102
rect 3927 9046 3995 9102
rect 4051 9046 4119 9102
rect 4175 9046 4243 9102
rect 4299 9046 4309 9102
rect 2497 8978 4309 9046
rect 2497 8922 2507 8978
rect 2563 8922 2631 8978
rect 2687 8922 2755 8978
rect 2811 8922 2879 8978
rect 2935 8922 3003 8978
rect 3059 8922 3127 8978
rect 3183 8922 3251 8978
rect 3307 8922 3375 8978
rect 3431 8922 3499 8978
rect 3555 8922 3623 8978
rect 3679 8922 3747 8978
rect 3803 8922 3871 8978
rect 3927 8922 3995 8978
rect 4051 8922 4119 8978
rect 4175 8922 4243 8978
rect 4299 8922 4309 8978
rect 2497 8854 4309 8922
rect 2497 8798 2507 8854
rect 2563 8798 2631 8854
rect 2687 8798 2755 8854
rect 2811 8798 2879 8854
rect 2935 8798 3003 8854
rect 3059 8798 3127 8854
rect 3183 8798 3251 8854
rect 3307 8798 3375 8854
rect 3431 8798 3499 8854
rect 3555 8798 3623 8854
rect 3679 8798 3747 8854
rect 3803 8798 3871 8854
rect 3927 8798 3995 8854
rect 4051 8798 4119 8854
rect 4175 8798 4243 8854
rect 4299 8798 4309 8854
rect 2497 8730 4309 8798
rect 2497 8674 2507 8730
rect 2563 8674 2631 8730
rect 2687 8674 2755 8730
rect 2811 8674 2879 8730
rect 2935 8674 3003 8730
rect 3059 8674 3127 8730
rect 3183 8674 3251 8730
rect 3307 8674 3375 8730
rect 3431 8674 3499 8730
rect 3555 8674 3623 8730
rect 3679 8674 3747 8730
rect 3803 8674 3871 8730
rect 3927 8674 3995 8730
rect 4051 8674 4119 8730
rect 4175 8674 4243 8730
rect 4299 8674 4309 8730
rect 2497 8606 4309 8674
rect 2497 8550 2507 8606
rect 2563 8550 2631 8606
rect 2687 8550 2755 8606
rect 2811 8550 2879 8606
rect 2935 8550 3003 8606
rect 3059 8550 3127 8606
rect 3183 8550 3251 8606
rect 3307 8550 3375 8606
rect 3431 8550 3499 8606
rect 3555 8550 3623 8606
rect 3679 8550 3747 8606
rect 3803 8550 3871 8606
rect 3927 8550 3995 8606
rect 4051 8550 4119 8606
rect 4175 8550 4243 8606
rect 4299 8550 4309 8606
rect 2497 8482 4309 8550
rect 2497 8426 2507 8482
rect 2563 8426 2631 8482
rect 2687 8426 2755 8482
rect 2811 8426 2879 8482
rect 2935 8426 3003 8482
rect 3059 8426 3127 8482
rect 3183 8426 3251 8482
rect 3307 8426 3375 8482
rect 3431 8426 3499 8482
rect 3555 8426 3623 8482
rect 3679 8426 3747 8482
rect 3803 8426 3871 8482
rect 3927 8426 3995 8482
rect 4051 8426 4119 8482
rect 4175 8426 4243 8482
rect 4299 8426 4309 8482
rect 2497 8358 4309 8426
rect 2497 8302 2507 8358
rect 2563 8302 2631 8358
rect 2687 8302 2755 8358
rect 2811 8302 2879 8358
rect 2935 8302 3003 8358
rect 3059 8302 3127 8358
rect 3183 8302 3251 8358
rect 3307 8302 3375 8358
rect 3431 8302 3499 8358
rect 3555 8302 3623 8358
rect 3679 8302 3747 8358
rect 3803 8302 3871 8358
rect 3927 8302 3995 8358
rect 4051 8302 4119 8358
rect 4175 8302 4243 8358
rect 4299 8302 4309 8358
rect 2497 8234 4309 8302
rect 2497 8178 2507 8234
rect 2563 8178 2631 8234
rect 2687 8178 2755 8234
rect 2811 8178 2879 8234
rect 2935 8178 3003 8234
rect 3059 8178 3127 8234
rect 3183 8178 3251 8234
rect 3307 8178 3375 8234
rect 3431 8178 3499 8234
rect 3555 8178 3623 8234
rect 3679 8178 3747 8234
rect 3803 8178 3871 8234
rect 3927 8178 3995 8234
rect 4051 8178 4119 8234
rect 4175 8178 4243 8234
rect 4299 8178 4309 8234
rect 2497 8110 4309 8178
rect 2497 8054 2507 8110
rect 2563 8054 2631 8110
rect 2687 8054 2755 8110
rect 2811 8054 2879 8110
rect 2935 8054 3003 8110
rect 3059 8054 3127 8110
rect 3183 8054 3251 8110
rect 3307 8054 3375 8110
rect 3431 8054 3499 8110
rect 3555 8054 3623 8110
rect 3679 8054 3747 8110
rect 3803 8054 3871 8110
rect 3927 8054 3995 8110
rect 4051 8054 4119 8110
rect 4175 8054 4243 8110
rect 4299 8054 4309 8110
rect 2497 7986 4309 8054
rect 2497 7930 2507 7986
rect 2563 7930 2631 7986
rect 2687 7930 2755 7986
rect 2811 7930 2879 7986
rect 2935 7930 3003 7986
rect 3059 7930 3127 7986
rect 3183 7930 3251 7986
rect 3307 7930 3375 7986
rect 3431 7930 3499 7986
rect 3555 7930 3623 7986
rect 3679 7930 3747 7986
rect 3803 7930 3871 7986
rect 3927 7930 3995 7986
rect 4051 7930 4119 7986
rect 4175 7930 4243 7986
rect 4299 7930 4309 7986
rect 2497 7862 4309 7930
rect 2497 7806 2507 7862
rect 2563 7806 2631 7862
rect 2687 7806 2755 7862
rect 2811 7806 2879 7862
rect 2935 7806 3003 7862
rect 3059 7806 3127 7862
rect 3183 7806 3251 7862
rect 3307 7806 3375 7862
rect 3431 7806 3499 7862
rect 3555 7806 3623 7862
rect 3679 7806 3747 7862
rect 3803 7806 3871 7862
rect 3927 7806 3995 7862
rect 4051 7806 4119 7862
rect 4175 7806 4243 7862
rect 4299 7806 4309 7862
rect 2497 7738 4309 7806
rect 2497 7682 2507 7738
rect 2563 7682 2631 7738
rect 2687 7682 2755 7738
rect 2811 7682 2879 7738
rect 2935 7682 3003 7738
rect 3059 7682 3127 7738
rect 3183 7682 3251 7738
rect 3307 7682 3375 7738
rect 3431 7682 3499 7738
rect 3555 7682 3623 7738
rect 3679 7682 3747 7738
rect 3803 7682 3871 7738
rect 3927 7682 3995 7738
rect 4051 7682 4119 7738
rect 4175 7682 4243 7738
rect 4299 7682 4309 7738
rect 2497 7614 4309 7682
rect 2497 7558 2507 7614
rect 2563 7558 2631 7614
rect 2687 7558 2755 7614
rect 2811 7558 2879 7614
rect 2935 7558 3003 7614
rect 3059 7558 3127 7614
rect 3183 7558 3251 7614
rect 3307 7558 3375 7614
rect 3431 7558 3499 7614
rect 3555 7558 3623 7614
rect 3679 7558 3747 7614
rect 3803 7558 3871 7614
rect 3927 7558 3995 7614
rect 4051 7558 4119 7614
rect 4175 7558 4243 7614
rect 4299 7558 4309 7614
rect 2497 7490 4309 7558
rect 2497 7434 2507 7490
rect 2563 7434 2631 7490
rect 2687 7434 2755 7490
rect 2811 7434 2879 7490
rect 2935 7434 3003 7490
rect 3059 7434 3127 7490
rect 3183 7434 3251 7490
rect 3307 7434 3375 7490
rect 3431 7434 3499 7490
rect 3555 7434 3623 7490
rect 3679 7434 3747 7490
rect 3803 7434 3871 7490
rect 3927 7434 3995 7490
rect 4051 7434 4119 7490
rect 4175 7434 4243 7490
rect 4299 7434 4309 7490
rect 2497 7366 4309 7434
rect 2497 7310 2507 7366
rect 2563 7310 2631 7366
rect 2687 7310 2755 7366
rect 2811 7310 2879 7366
rect 2935 7310 3003 7366
rect 3059 7310 3127 7366
rect 3183 7310 3251 7366
rect 3307 7310 3375 7366
rect 3431 7310 3499 7366
rect 3555 7310 3623 7366
rect 3679 7310 3747 7366
rect 3803 7310 3871 7366
rect 3927 7310 3995 7366
rect 4051 7310 4119 7366
rect 4175 7310 4243 7366
rect 4299 7310 4309 7366
rect 2497 7242 4309 7310
rect 2497 7186 2507 7242
rect 2563 7186 2631 7242
rect 2687 7186 2755 7242
rect 2811 7186 2879 7242
rect 2935 7186 3003 7242
rect 3059 7186 3127 7242
rect 3183 7186 3251 7242
rect 3307 7186 3375 7242
rect 3431 7186 3499 7242
rect 3555 7186 3623 7242
rect 3679 7186 3747 7242
rect 3803 7186 3871 7242
rect 3927 7186 3995 7242
rect 4051 7186 4119 7242
rect 4175 7186 4243 7242
rect 4299 7186 4309 7242
rect 2497 7118 4309 7186
rect 2497 7062 2507 7118
rect 2563 7062 2631 7118
rect 2687 7062 2755 7118
rect 2811 7062 2879 7118
rect 2935 7062 3003 7118
rect 3059 7062 3127 7118
rect 3183 7062 3251 7118
rect 3307 7062 3375 7118
rect 3431 7062 3499 7118
rect 3555 7062 3623 7118
rect 3679 7062 3747 7118
rect 3803 7062 3871 7118
rect 3927 7062 3995 7118
rect 4051 7062 4119 7118
rect 4175 7062 4243 7118
rect 4299 7062 4309 7118
rect 2497 6994 4309 7062
rect 2497 6938 2507 6994
rect 2563 6938 2631 6994
rect 2687 6938 2755 6994
rect 2811 6938 2879 6994
rect 2935 6938 3003 6994
rect 3059 6938 3127 6994
rect 3183 6938 3251 6994
rect 3307 6938 3375 6994
rect 3431 6938 3499 6994
rect 3555 6938 3623 6994
rect 3679 6938 3747 6994
rect 3803 6938 3871 6994
rect 3927 6938 3995 6994
rect 4051 6938 4119 6994
rect 4175 6938 4243 6994
rect 4299 6938 4309 6994
rect 2497 6870 4309 6938
rect 2497 6814 2507 6870
rect 2563 6814 2631 6870
rect 2687 6814 2755 6870
rect 2811 6814 2879 6870
rect 2935 6814 3003 6870
rect 3059 6814 3127 6870
rect 3183 6814 3251 6870
rect 3307 6814 3375 6870
rect 3431 6814 3499 6870
rect 3555 6814 3623 6870
rect 3679 6814 3747 6870
rect 3803 6814 3871 6870
rect 3927 6814 3995 6870
rect 4051 6814 4119 6870
rect 4175 6814 4243 6870
rect 4299 6814 4309 6870
rect 2497 6746 4309 6814
rect 2497 6690 2507 6746
rect 2563 6690 2631 6746
rect 2687 6690 2755 6746
rect 2811 6690 2879 6746
rect 2935 6690 3003 6746
rect 3059 6690 3127 6746
rect 3183 6690 3251 6746
rect 3307 6690 3375 6746
rect 3431 6690 3499 6746
rect 3555 6690 3623 6746
rect 3679 6690 3747 6746
rect 3803 6690 3871 6746
rect 3927 6690 3995 6746
rect 4051 6690 4119 6746
rect 4175 6690 4243 6746
rect 4299 6690 4309 6746
rect 2497 6622 4309 6690
rect 2497 6566 2507 6622
rect 2563 6566 2631 6622
rect 2687 6566 2755 6622
rect 2811 6566 2879 6622
rect 2935 6566 3003 6622
rect 3059 6566 3127 6622
rect 3183 6566 3251 6622
rect 3307 6566 3375 6622
rect 3431 6566 3499 6622
rect 3555 6566 3623 6622
rect 3679 6566 3747 6622
rect 3803 6566 3871 6622
rect 3927 6566 3995 6622
rect 4051 6566 4119 6622
rect 4175 6566 4243 6622
rect 4299 6566 4309 6622
rect 2497 6498 4309 6566
rect 2497 6442 2507 6498
rect 2563 6442 2631 6498
rect 2687 6442 2755 6498
rect 2811 6442 2879 6498
rect 2935 6442 3003 6498
rect 3059 6442 3127 6498
rect 3183 6442 3251 6498
rect 3307 6442 3375 6498
rect 3431 6442 3499 6498
rect 3555 6442 3623 6498
rect 3679 6442 3747 6498
rect 3803 6442 3871 6498
rect 3927 6442 3995 6498
rect 4051 6442 4119 6498
rect 4175 6442 4243 6498
rect 4299 6442 4309 6498
rect 2497 6432 4309 6442
rect 6358 9350 7426 9360
rect 6358 9294 6368 9350
rect 6424 9294 6492 9350
rect 6548 9294 6616 9350
rect 6672 9294 6740 9350
rect 6796 9294 6864 9350
rect 6920 9294 6988 9350
rect 7044 9294 7112 9350
rect 7168 9294 7236 9350
rect 7292 9294 7360 9350
rect 7416 9294 7426 9350
rect 6358 9226 7426 9294
rect 6358 9170 6368 9226
rect 6424 9170 6492 9226
rect 6548 9170 6616 9226
rect 6672 9170 6740 9226
rect 6796 9170 6864 9226
rect 6920 9170 6988 9226
rect 7044 9170 7112 9226
rect 7168 9170 7236 9226
rect 7292 9170 7360 9226
rect 7416 9170 7426 9226
rect 6358 9102 7426 9170
rect 6358 9046 6368 9102
rect 6424 9046 6492 9102
rect 6548 9046 6616 9102
rect 6672 9046 6740 9102
rect 6796 9046 6864 9102
rect 6920 9046 6988 9102
rect 7044 9046 7112 9102
rect 7168 9046 7236 9102
rect 7292 9046 7360 9102
rect 7416 9046 7426 9102
rect 6358 8978 7426 9046
rect 6358 8922 6368 8978
rect 6424 8922 6492 8978
rect 6548 8922 6616 8978
rect 6672 8922 6740 8978
rect 6796 8922 6864 8978
rect 6920 8922 6988 8978
rect 7044 8922 7112 8978
rect 7168 8922 7236 8978
rect 7292 8922 7360 8978
rect 7416 8922 7426 8978
rect 6358 8854 7426 8922
rect 6358 8798 6368 8854
rect 6424 8798 6492 8854
rect 6548 8798 6616 8854
rect 6672 8798 6740 8854
rect 6796 8798 6864 8854
rect 6920 8798 6988 8854
rect 7044 8798 7112 8854
rect 7168 8798 7236 8854
rect 7292 8798 7360 8854
rect 7416 8798 7426 8854
rect 6358 8730 7426 8798
rect 6358 8674 6368 8730
rect 6424 8674 6492 8730
rect 6548 8674 6616 8730
rect 6672 8674 6740 8730
rect 6796 8674 6864 8730
rect 6920 8674 6988 8730
rect 7044 8674 7112 8730
rect 7168 8674 7236 8730
rect 7292 8674 7360 8730
rect 7416 8674 7426 8730
rect 6358 8606 7426 8674
rect 6358 8550 6368 8606
rect 6424 8550 6492 8606
rect 6548 8550 6616 8606
rect 6672 8550 6740 8606
rect 6796 8550 6864 8606
rect 6920 8550 6988 8606
rect 7044 8550 7112 8606
rect 7168 8550 7236 8606
rect 7292 8550 7360 8606
rect 7416 8550 7426 8606
rect 6358 8482 7426 8550
rect 6358 8426 6368 8482
rect 6424 8426 6492 8482
rect 6548 8426 6616 8482
rect 6672 8426 6740 8482
rect 6796 8426 6864 8482
rect 6920 8426 6988 8482
rect 7044 8426 7112 8482
rect 7168 8426 7236 8482
rect 7292 8426 7360 8482
rect 7416 8426 7426 8482
rect 6358 8358 7426 8426
rect 6358 8302 6368 8358
rect 6424 8302 6492 8358
rect 6548 8302 6616 8358
rect 6672 8302 6740 8358
rect 6796 8302 6864 8358
rect 6920 8302 6988 8358
rect 7044 8302 7112 8358
rect 7168 8302 7236 8358
rect 7292 8302 7360 8358
rect 7416 8302 7426 8358
rect 6358 8234 7426 8302
rect 6358 8178 6368 8234
rect 6424 8178 6492 8234
rect 6548 8178 6616 8234
rect 6672 8178 6740 8234
rect 6796 8178 6864 8234
rect 6920 8178 6988 8234
rect 7044 8178 7112 8234
rect 7168 8178 7236 8234
rect 7292 8178 7360 8234
rect 7416 8178 7426 8234
rect 6358 8110 7426 8178
rect 6358 8054 6368 8110
rect 6424 8054 6492 8110
rect 6548 8054 6616 8110
rect 6672 8054 6740 8110
rect 6796 8054 6864 8110
rect 6920 8054 6988 8110
rect 7044 8054 7112 8110
rect 7168 8054 7236 8110
rect 7292 8054 7360 8110
rect 7416 8054 7426 8110
rect 6358 7986 7426 8054
rect 6358 7930 6368 7986
rect 6424 7930 6492 7986
rect 6548 7930 6616 7986
rect 6672 7930 6740 7986
rect 6796 7930 6864 7986
rect 6920 7930 6988 7986
rect 7044 7930 7112 7986
rect 7168 7930 7236 7986
rect 7292 7930 7360 7986
rect 7416 7930 7426 7986
rect 6358 7862 7426 7930
rect 6358 7806 6368 7862
rect 6424 7806 6492 7862
rect 6548 7806 6616 7862
rect 6672 7806 6740 7862
rect 6796 7806 6864 7862
rect 6920 7806 6988 7862
rect 7044 7806 7112 7862
rect 7168 7806 7236 7862
rect 7292 7806 7360 7862
rect 7416 7806 7426 7862
rect 6358 7738 7426 7806
rect 6358 7682 6368 7738
rect 6424 7682 6492 7738
rect 6548 7682 6616 7738
rect 6672 7682 6740 7738
rect 6796 7682 6864 7738
rect 6920 7682 6988 7738
rect 7044 7682 7112 7738
rect 7168 7682 7236 7738
rect 7292 7682 7360 7738
rect 7416 7682 7426 7738
rect 6358 7614 7426 7682
rect 6358 7558 6368 7614
rect 6424 7558 6492 7614
rect 6548 7558 6616 7614
rect 6672 7558 6740 7614
rect 6796 7558 6864 7614
rect 6920 7558 6988 7614
rect 7044 7558 7112 7614
rect 7168 7558 7236 7614
rect 7292 7558 7360 7614
rect 7416 7558 7426 7614
rect 6358 7490 7426 7558
rect 6358 7434 6368 7490
rect 6424 7434 6492 7490
rect 6548 7434 6616 7490
rect 6672 7434 6740 7490
rect 6796 7434 6864 7490
rect 6920 7434 6988 7490
rect 7044 7434 7112 7490
rect 7168 7434 7236 7490
rect 7292 7434 7360 7490
rect 7416 7434 7426 7490
rect 6358 7366 7426 7434
rect 6358 7310 6368 7366
rect 6424 7310 6492 7366
rect 6548 7310 6616 7366
rect 6672 7310 6740 7366
rect 6796 7310 6864 7366
rect 6920 7310 6988 7366
rect 7044 7310 7112 7366
rect 7168 7310 7236 7366
rect 7292 7310 7360 7366
rect 7416 7310 7426 7366
rect 6358 7242 7426 7310
rect 6358 7186 6368 7242
rect 6424 7186 6492 7242
rect 6548 7186 6616 7242
rect 6672 7186 6740 7242
rect 6796 7186 6864 7242
rect 6920 7186 6988 7242
rect 7044 7186 7112 7242
rect 7168 7186 7236 7242
rect 7292 7186 7360 7242
rect 7416 7186 7426 7242
rect 6358 7118 7426 7186
rect 6358 7062 6368 7118
rect 6424 7062 6492 7118
rect 6548 7062 6616 7118
rect 6672 7062 6740 7118
rect 6796 7062 6864 7118
rect 6920 7062 6988 7118
rect 7044 7062 7112 7118
rect 7168 7062 7236 7118
rect 7292 7062 7360 7118
rect 7416 7062 7426 7118
rect 6358 6994 7426 7062
rect 6358 6938 6368 6994
rect 6424 6938 6492 6994
rect 6548 6938 6616 6994
rect 6672 6938 6740 6994
rect 6796 6938 6864 6994
rect 6920 6938 6988 6994
rect 7044 6938 7112 6994
rect 7168 6938 7236 6994
rect 7292 6938 7360 6994
rect 7416 6938 7426 6994
rect 6358 6870 7426 6938
rect 6358 6814 6368 6870
rect 6424 6814 6492 6870
rect 6548 6814 6616 6870
rect 6672 6814 6740 6870
rect 6796 6814 6864 6870
rect 6920 6814 6988 6870
rect 7044 6814 7112 6870
rect 7168 6814 7236 6870
rect 7292 6814 7360 6870
rect 7416 6814 7426 6870
rect 6358 6746 7426 6814
rect 6358 6690 6368 6746
rect 6424 6690 6492 6746
rect 6548 6690 6616 6746
rect 6672 6690 6740 6746
rect 6796 6690 6864 6746
rect 6920 6690 6988 6746
rect 7044 6690 7112 6746
rect 7168 6690 7236 6746
rect 7292 6690 7360 6746
rect 7416 6690 7426 6746
rect 6358 6622 7426 6690
rect 6358 6566 6368 6622
rect 6424 6566 6492 6622
rect 6548 6566 6616 6622
rect 6672 6566 6740 6622
rect 6796 6566 6864 6622
rect 6920 6566 6988 6622
rect 7044 6566 7112 6622
rect 7168 6566 7236 6622
rect 7292 6566 7360 6622
rect 7416 6566 7426 6622
rect 6358 6498 7426 6566
rect 6358 6442 6368 6498
rect 6424 6442 6492 6498
rect 6548 6442 6616 6498
rect 6672 6442 6740 6498
rect 6796 6442 6864 6498
rect 6920 6442 6988 6498
rect 7044 6442 7112 6498
rect 7168 6442 7236 6498
rect 7292 6442 7360 6498
rect 7416 6442 7426 6498
rect 6358 6432 7426 6442
rect 8741 9350 10553 9360
rect 8741 9294 8751 9350
rect 8807 9294 8875 9350
rect 8931 9294 8999 9350
rect 9055 9294 9123 9350
rect 9179 9294 9247 9350
rect 9303 9294 9371 9350
rect 9427 9294 9495 9350
rect 9551 9294 9619 9350
rect 9675 9294 9743 9350
rect 9799 9294 9867 9350
rect 9923 9294 9991 9350
rect 10047 9294 10115 9350
rect 10171 9294 10239 9350
rect 10295 9294 10363 9350
rect 10419 9294 10487 9350
rect 10543 9294 10553 9350
rect 8741 9226 10553 9294
rect 8741 9170 8751 9226
rect 8807 9170 8875 9226
rect 8931 9170 8999 9226
rect 9055 9170 9123 9226
rect 9179 9170 9247 9226
rect 9303 9170 9371 9226
rect 9427 9170 9495 9226
rect 9551 9170 9619 9226
rect 9675 9170 9743 9226
rect 9799 9170 9867 9226
rect 9923 9170 9991 9226
rect 10047 9170 10115 9226
rect 10171 9170 10239 9226
rect 10295 9170 10363 9226
rect 10419 9170 10487 9226
rect 10543 9170 10553 9226
rect 8741 9102 10553 9170
rect 8741 9046 8751 9102
rect 8807 9046 8875 9102
rect 8931 9046 8999 9102
rect 9055 9046 9123 9102
rect 9179 9046 9247 9102
rect 9303 9046 9371 9102
rect 9427 9046 9495 9102
rect 9551 9046 9619 9102
rect 9675 9046 9743 9102
rect 9799 9046 9867 9102
rect 9923 9046 9991 9102
rect 10047 9046 10115 9102
rect 10171 9046 10239 9102
rect 10295 9046 10363 9102
rect 10419 9046 10487 9102
rect 10543 9046 10553 9102
rect 8741 8978 10553 9046
rect 8741 8922 8751 8978
rect 8807 8922 8875 8978
rect 8931 8922 8999 8978
rect 9055 8922 9123 8978
rect 9179 8922 9247 8978
rect 9303 8922 9371 8978
rect 9427 8922 9495 8978
rect 9551 8922 9619 8978
rect 9675 8922 9743 8978
rect 9799 8922 9867 8978
rect 9923 8922 9991 8978
rect 10047 8922 10115 8978
rect 10171 8922 10239 8978
rect 10295 8922 10363 8978
rect 10419 8922 10487 8978
rect 10543 8922 10553 8978
rect 8741 8854 10553 8922
rect 8741 8798 8751 8854
rect 8807 8798 8875 8854
rect 8931 8798 8999 8854
rect 9055 8798 9123 8854
rect 9179 8798 9247 8854
rect 9303 8798 9371 8854
rect 9427 8798 9495 8854
rect 9551 8798 9619 8854
rect 9675 8798 9743 8854
rect 9799 8798 9867 8854
rect 9923 8798 9991 8854
rect 10047 8798 10115 8854
rect 10171 8798 10239 8854
rect 10295 8798 10363 8854
rect 10419 8798 10487 8854
rect 10543 8798 10553 8854
rect 8741 8730 10553 8798
rect 8741 8674 8751 8730
rect 8807 8674 8875 8730
rect 8931 8674 8999 8730
rect 9055 8674 9123 8730
rect 9179 8674 9247 8730
rect 9303 8674 9371 8730
rect 9427 8674 9495 8730
rect 9551 8674 9619 8730
rect 9675 8674 9743 8730
rect 9799 8674 9867 8730
rect 9923 8674 9991 8730
rect 10047 8674 10115 8730
rect 10171 8674 10239 8730
rect 10295 8674 10363 8730
rect 10419 8674 10487 8730
rect 10543 8674 10553 8730
rect 8741 8606 10553 8674
rect 8741 8550 8751 8606
rect 8807 8550 8875 8606
rect 8931 8550 8999 8606
rect 9055 8550 9123 8606
rect 9179 8550 9247 8606
rect 9303 8550 9371 8606
rect 9427 8550 9495 8606
rect 9551 8550 9619 8606
rect 9675 8550 9743 8606
rect 9799 8550 9867 8606
rect 9923 8550 9991 8606
rect 10047 8550 10115 8606
rect 10171 8550 10239 8606
rect 10295 8550 10363 8606
rect 10419 8550 10487 8606
rect 10543 8550 10553 8606
rect 8741 8482 10553 8550
rect 8741 8426 8751 8482
rect 8807 8426 8875 8482
rect 8931 8426 8999 8482
rect 9055 8426 9123 8482
rect 9179 8426 9247 8482
rect 9303 8426 9371 8482
rect 9427 8426 9495 8482
rect 9551 8426 9619 8482
rect 9675 8426 9743 8482
rect 9799 8426 9867 8482
rect 9923 8426 9991 8482
rect 10047 8426 10115 8482
rect 10171 8426 10239 8482
rect 10295 8426 10363 8482
rect 10419 8426 10487 8482
rect 10543 8426 10553 8482
rect 8741 8358 10553 8426
rect 8741 8302 8751 8358
rect 8807 8302 8875 8358
rect 8931 8302 8999 8358
rect 9055 8302 9123 8358
rect 9179 8302 9247 8358
rect 9303 8302 9371 8358
rect 9427 8302 9495 8358
rect 9551 8302 9619 8358
rect 9675 8302 9743 8358
rect 9799 8302 9867 8358
rect 9923 8302 9991 8358
rect 10047 8302 10115 8358
rect 10171 8302 10239 8358
rect 10295 8302 10363 8358
rect 10419 8302 10487 8358
rect 10543 8302 10553 8358
rect 8741 8234 10553 8302
rect 8741 8178 8751 8234
rect 8807 8178 8875 8234
rect 8931 8178 8999 8234
rect 9055 8178 9123 8234
rect 9179 8178 9247 8234
rect 9303 8178 9371 8234
rect 9427 8178 9495 8234
rect 9551 8178 9619 8234
rect 9675 8178 9743 8234
rect 9799 8178 9867 8234
rect 9923 8178 9991 8234
rect 10047 8178 10115 8234
rect 10171 8178 10239 8234
rect 10295 8178 10363 8234
rect 10419 8178 10487 8234
rect 10543 8178 10553 8234
rect 8741 8110 10553 8178
rect 8741 8054 8751 8110
rect 8807 8054 8875 8110
rect 8931 8054 8999 8110
rect 9055 8054 9123 8110
rect 9179 8054 9247 8110
rect 9303 8054 9371 8110
rect 9427 8054 9495 8110
rect 9551 8054 9619 8110
rect 9675 8054 9743 8110
rect 9799 8054 9867 8110
rect 9923 8054 9991 8110
rect 10047 8054 10115 8110
rect 10171 8054 10239 8110
rect 10295 8054 10363 8110
rect 10419 8054 10487 8110
rect 10543 8054 10553 8110
rect 8741 7986 10553 8054
rect 8741 7930 8751 7986
rect 8807 7930 8875 7986
rect 8931 7930 8999 7986
rect 9055 7930 9123 7986
rect 9179 7930 9247 7986
rect 9303 7930 9371 7986
rect 9427 7930 9495 7986
rect 9551 7930 9619 7986
rect 9675 7930 9743 7986
rect 9799 7930 9867 7986
rect 9923 7930 9991 7986
rect 10047 7930 10115 7986
rect 10171 7930 10239 7986
rect 10295 7930 10363 7986
rect 10419 7930 10487 7986
rect 10543 7930 10553 7986
rect 8741 7862 10553 7930
rect 8741 7806 8751 7862
rect 8807 7806 8875 7862
rect 8931 7806 8999 7862
rect 9055 7806 9123 7862
rect 9179 7806 9247 7862
rect 9303 7806 9371 7862
rect 9427 7806 9495 7862
rect 9551 7806 9619 7862
rect 9675 7806 9743 7862
rect 9799 7806 9867 7862
rect 9923 7806 9991 7862
rect 10047 7806 10115 7862
rect 10171 7806 10239 7862
rect 10295 7806 10363 7862
rect 10419 7806 10487 7862
rect 10543 7806 10553 7862
rect 8741 7738 10553 7806
rect 8741 7682 8751 7738
rect 8807 7682 8875 7738
rect 8931 7682 8999 7738
rect 9055 7682 9123 7738
rect 9179 7682 9247 7738
rect 9303 7682 9371 7738
rect 9427 7682 9495 7738
rect 9551 7682 9619 7738
rect 9675 7682 9743 7738
rect 9799 7682 9867 7738
rect 9923 7682 9991 7738
rect 10047 7682 10115 7738
rect 10171 7682 10239 7738
rect 10295 7682 10363 7738
rect 10419 7682 10487 7738
rect 10543 7682 10553 7738
rect 8741 7614 10553 7682
rect 8741 7558 8751 7614
rect 8807 7558 8875 7614
rect 8931 7558 8999 7614
rect 9055 7558 9123 7614
rect 9179 7558 9247 7614
rect 9303 7558 9371 7614
rect 9427 7558 9495 7614
rect 9551 7558 9619 7614
rect 9675 7558 9743 7614
rect 9799 7558 9867 7614
rect 9923 7558 9991 7614
rect 10047 7558 10115 7614
rect 10171 7558 10239 7614
rect 10295 7558 10363 7614
rect 10419 7558 10487 7614
rect 10543 7558 10553 7614
rect 8741 7490 10553 7558
rect 8741 7434 8751 7490
rect 8807 7434 8875 7490
rect 8931 7434 8999 7490
rect 9055 7434 9123 7490
rect 9179 7434 9247 7490
rect 9303 7434 9371 7490
rect 9427 7434 9495 7490
rect 9551 7434 9619 7490
rect 9675 7434 9743 7490
rect 9799 7434 9867 7490
rect 9923 7434 9991 7490
rect 10047 7434 10115 7490
rect 10171 7434 10239 7490
rect 10295 7434 10363 7490
rect 10419 7434 10487 7490
rect 10543 7434 10553 7490
rect 8741 7366 10553 7434
rect 8741 7310 8751 7366
rect 8807 7310 8875 7366
rect 8931 7310 8999 7366
rect 9055 7310 9123 7366
rect 9179 7310 9247 7366
rect 9303 7310 9371 7366
rect 9427 7310 9495 7366
rect 9551 7310 9619 7366
rect 9675 7310 9743 7366
rect 9799 7310 9867 7366
rect 9923 7310 9991 7366
rect 10047 7310 10115 7366
rect 10171 7310 10239 7366
rect 10295 7310 10363 7366
rect 10419 7310 10487 7366
rect 10543 7310 10553 7366
rect 8741 7242 10553 7310
rect 8741 7186 8751 7242
rect 8807 7186 8875 7242
rect 8931 7186 8999 7242
rect 9055 7186 9123 7242
rect 9179 7186 9247 7242
rect 9303 7186 9371 7242
rect 9427 7186 9495 7242
rect 9551 7186 9619 7242
rect 9675 7186 9743 7242
rect 9799 7186 9867 7242
rect 9923 7186 9991 7242
rect 10047 7186 10115 7242
rect 10171 7186 10239 7242
rect 10295 7186 10363 7242
rect 10419 7186 10487 7242
rect 10543 7186 10553 7242
rect 8741 7118 10553 7186
rect 8741 7062 8751 7118
rect 8807 7062 8875 7118
rect 8931 7062 8999 7118
rect 9055 7062 9123 7118
rect 9179 7062 9247 7118
rect 9303 7062 9371 7118
rect 9427 7062 9495 7118
rect 9551 7062 9619 7118
rect 9675 7062 9743 7118
rect 9799 7062 9867 7118
rect 9923 7062 9991 7118
rect 10047 7062 10115 7118
rect 10171 7062 10239 7118
rect 10295 7062 10363 7118
rect 10419 7062 10487 7118
rect 10543 7062 10553 7118
rect 8741 6994 10553 7062
rect 8741 6938 8751 6994
rect 8807 6938 8875 6994
rect 8931 6938 8999 6994
rect 9055 6938 9123 6994
rect 9179 6938 9247 6994
rect 9303 6938 9371 6994
rect 9427 6938 9495 6994
rect 9551 6938 9619 6994
rect 9675 6938 9743 6994
rect 9799 6938 9867 6994
rect 9923 6938 9991 6994
rect 10047 6938 10115 6994
rect 10171 6938 10239 6994
rect 10295 6938 10363 6994
rect 10419 6938 10487 6994
rect 10543 6938 10553 6994
rect 8741 6870 10553 6938
rect 8741 6814 8751 6870
rect 8807 6814 8875 6870
rect 8931 6814 8999 6870
rect 9055 6814 9123 6870
rect 9179 6814 9247 6870
rect 9303 6814 9371 6870
rect 9427 6814 9495 6870
rect 9551 6814 9619 6870
rect 9675 6814 9743 6870
rect 9799 6814 9867 6870
rect 9923 6814 9991 6870
rect 10047 6814 10115 6870
rect 10171 6814 10239 6870
rect 10295 6814 10363 6870
rect 10419 6814 10487 6870
rect 10543 6814 10553 6870
rect 8741 6746 10553 6814
rect 8741 6690 8751 6746
rect 8807 6690 8875 6746
rect 8931 6690 8999 6746
rect 9055 6690 9123 6746
rect 9179 6690 9247 6746
rect 9303 6690 9371 6746
rect 9427 6690 9495 6746
rect 9551 6690 9619 6746
rect 9675 6690 9743 6746
rect 9799 6690 9867 6746
rect 9923 6690 9991 6746
rect 10047 6690 10115 6746
rect 10171 6690 10239 6746
rect 10295 6690 10363 6746
rect 10419 6690 10487 6746
rect 10543 6690 10553 6746
rect 8741 6622 10553 6690
rect 8741 6566 8751 6622
rect 8807 6566 8875 6622
rect 8931 6566 8999 6622
rect 9055 6566 9123 6622
rect 9179 6566 9247 6622
rect 9303 6566 9371 6622
rect 9427 6566 9495 6622
rect 9551 6566 9619 6622
rect 9675 6566 9743 6622
rect 9799 6566 9867 6622
rect 9923 6566 9991 6622
rect 10047 6566 10115 6622
rect 10171 6566 10239 6622
rect 10295 6566 10363 6622
rect 10419 6566 10487 6622
rect 10543 6566 10553 6622
rect 8741 6498 10553 6566
rect 8741 6442 8751 6498
rect 8807 6442 8875 6498
rect 8931 6442 8999 6498
rect 9055 6442 9123 6498
rect 9179 6442 9247 6498
rect 9303 6442 9371 6498
rect 9427 6442 9495 6498
rect 9551 6442 9619 6498
rect 9675 6442 9743 6498
rect 9799 6442 9867 6498
rect 9923 6442 9991 6498
rect 10047 6442 10115 6498
rect 10171 6442 10239 6498
rect 10295 6442 10363 6498
rect 10419 6442 10487 6498
rect 10543 6442 10553 6498
rect 8741 6432 10553 6442
rect 12842 9350 13910 9360
rect 12842 9294 12852 9350
rect 12908 9294 12976 9350
rect 13032 9294 13100 9350
rect 13156 9294 13224 9350
rect 13280 9294 13348 9350
rect 13404 9294 13472 9350
rect 13528 9294 13596 9350
rect 13652 9294 13720 9350
rect 13776 9294 13844 9350
rect 13900 9294 13910 9350
rect 12842 9226 13910 9294
rect 12842 9170 12852 9226
rect 12908 9170 12976 9226
rect 13032 9170 13100 9226
rect 13156 9170 13224 9226
rect 13280 9170 13348 9226
rect 13404 9170 13472 9226
rect 13528 9170 13596 9226
rect 13652 9170 13720 9226
rect 13776 9170 13844 9226
rect 13900 9170 13910 9226
rect 12842 9102 13910 9170
rect 12842 9046 12852 9102
rect 12908 9046 12976 9102
rect 13032 9046 13100 9102
rect 13156 9046 13224 9102
rect 13280 9046 13348 9102
rect 13404 9046 13472 9102
rect 13528 9046 13596 9102
rect 13652 9046 13720 9102
rect 13776 9046 13844 9102
rect 13900 9046 13910 9102
rect 12842 8978 13910 9046
rect 12842 8922 12852 8978
rect 12908 8922 12976 8978
rect 13032 8922 13100 8978
rect 13156 8922 13224 8978
rect 13280 8922 13348 8978
rect 13404 8922 13472 8978
rect 13528 8922 13596 8978
rect 13652 8922 13720 8978
rect 13776 8922 13844 8978
rect 13900 8922 13910 8978
rect 12842 8854 13910 8922
rect 12842 8798 12852 8854
rect 12908 8798 12976 8854
rect 13032 8798 13100 8854
rect 13156 8798 13224 8854
rect 13280 8798 13348 8854
rect 13404 8798 13472 8854
rect 13528 8798 13596 8854
rect 13652 8798 13720 8854
rect 13776 8798 13844 8854
rect 13900 8798 13910 8854
rect 12842 8730 13910 8798
rect 12842 8674 12852 8730
rect 12908 8674 12976 8730
rect 13032 8674 13100 8730
rect 13156 8674 13224 8730
rect 13280 8674 13348 8730
rect 13404 8674 13472 8730
rect 13528 8674 13596 8730
rect 13652 8674 13720 8730
rect 13776 8674 13844 8730
rect 13900 8674 13910 8730
rect 12842 8606 13910 8674
rect 12842 8550 12852 8606
rect 12908 8550 12976 8606
rect 13032 8550 13100 8606
rect 13156 8550 13224 8606
rect 13280 8550 13348 8606
rect 13404 8550 13472 8606
rect 13528 8550 13596 8606
rect 13652 8550 13720 8606
rect 13776 8550 13844 8606
rect 13900 8550 13910 8606
rect 12842 8482 13910 8550
rect 12842 8426 12852 8482
rect 12908 8426 12976 8482
rect 13032 8426 13100 8482
rect 13156 8426 13224 8482
rect 13280 8426 13348 8482
rect 13404 8426 13472 8482
rect 13528 8426 13596 8482
rect 13652 8426 13720 8482
rect 13776 8426 13844 8482
rect 13900 8426 13910 8482
rect 12842 8358 13910 8426
rect 12842 8302 12852 8358
rect 12908 8302 12976 8358
rect 13032 8302 13100 8358
rect 13156 8302 13224 8358
rect 13280 8302 13348 8358
rect 13404 8302 13472 8358
rect 13528 8302 13596 8358
rect 13652 8302 13720 8358
rect 13776 8302 13844 8358
rect 13900 8302 13910 8358
rect 12842 8234 13910 8302
rect 12842 8178 12852 8234
rect 12908 8178 12976 8234
rect 13032 8178 13100 8234
rect 13156 8178 13224 8234
rect 13280 8178 13348 8234
rect 13404 8178 13472 8234
rect 13528 8178 13596 8234
rect 13652 8178 13720 8234
rect 13776 8178 13844 8234
rect 13900 8178 13910 8234
rect 12842 8110 13910 8178
rect 12842 8054 12852 8110
rect 12908 8054 12976 8110
rect 13032 8054 13100 8110
rect 13156 8054 13224 8110
rect 13280 8054 13348 8110
rect 13404 8054 13472 8110
rect 13528 8054 13596 8110
rect 13652 8054 13720 8110
rect 13776 8054 13844 8110
rect 13900 8054 13910 8110
rect 12842 7986 13910 8054
rect 12842 7930 12852 7986
rect 12908 7930 12976 7986
rect 13032 7930 13100 7986
rect 13156 7930 13224 7986
rect 13280 7930 13348 7986
rect 13404 7930 13472 7986
rect 13528 7930 13596 7986
rect 13652 7930 13720 7986
rect 13776 7930 13844 7986
rect 13900 7930 13910 7986
rect 12842 7862 13910 7930
rect 12842 7806 12852 7862
rect 12908 7806 12976 7862
rect 13032 7806 13100 7862
rect 13156 7806 13224 7862
rect 13280 7806 13348 7862
rect 13404 7806 13472 7862
rect 13528 7806 13596 7862
rect 13652 7806 13720 7862
rect 13776 7806 13844 7862
rect 13900 7806 13910 7862
rect 12842 7738 13910 7806
rect 12842 7682 12852 7738
rect 12908 7682 12976 7738
rect 13032 7682 13100 7738
rect 13156 7682 13224 7738
rect 13280 7682 13348 7738
rect 13404 7682 13472 7738
rect 13528 7682 13596 7738
rect 13652 7682 13720 7738
rect 13776 7682 13844 7738
rect 13900 7682 13910 7738
rect 12842 7614 13910 7682
rect 12842 7558 12852 7614
rect 12908 7558 12976 7614
rect 13032 7558 13100 7614
rect 13156 7558 13224 7614
rect 13280 7558 13348 7614
rect 13404 7558 13472 7614
rect 13528 7558 13596 7614
rect 13652 7558 13720 7614
rect 13776 7558 13844 7614
rect 13900 7558 13910 7614
rect 12842 7490 13910 7558
rect 12842 7434 12852 7490
rect 12908 7434 12976 7490
rect 13032 7434 13100 7490
rect 13156 7434 13224 7490
rect 13280 7434 13348 7490
rect 13404 7434 13472 7490
rect 13528 7434 13596 7490
rect 13652 7434 13720 7490
rect 13776 7434 13844 7490
rect 13900 7434 13910 7490
rect 12842 7366 13910 7434
rect 12842 7310 12852 7366
rect 12908 7310 12976 7366
rect 13032 7310 13100 7366
rect 13156 7310 13224 7366
rect 13280 7310 13348 7366
rect 13404 7310 13472 7366
rect 13528 7310 13596 7366
rect 13652 7310 13720 7366
rect 13776 7310 13844 7366
rect 13900 7310 13910 7366
rect 12842 7242 13910 7310
rect 12842 7186 12852 7242
rect 12908 7186 12976 7242
rect 13032 7186 13100 7242
rect 13156 7186 13224 7242
rect 13280 7186 13348 7242
rect 13404 7186 13472 7242
rect 13528 7186 13596 7242
rect 13652 7186 13720 7242
rect 13776 7186 13844 7242
rect 13900 7186 13910 7242
rect 12842 7118 13910 7186
rect 12842 7062 12852 7118
rect 12908 7062 12976 7118
rect 13032 7062 13100 7118
rect 13156 7062 13224 7118
rect 13280 7062 13348 7118
rect 13404 7062 13472 7118
rect 13528 7062 13596 7118
rect 13652 7062 13720 7118
rect 13776 7062 13844 7118
rect 13900 7062 13910 7118
rect 12842 6994 13910 7062
rect 12842 6938 12852 6994
rect 12908 6938 12976 6994
rect 13032 6938 13100 6994
rect 13156 6938 13224 6994
rect 13280 6938 13348 6994
rect 13404 6938 13472 6994
rect 13528 6938 13596 6994
rect 13652 6938 13720 6994
rect 13776 6938 13844 6994
rect 13900 6938 13910 6994
rect 12842 6870 13910 6938
rect 12842 6814 12852 6870
rect 12908 6814 12976 6870
rect 13032 6814 13100 6870
rect 13156 6814 13224 6870
rect 13280 6814 13348 6870
rect 13404 6814 13472 6870
rect 13528 6814 13596 6870
rect 13652 6814 13720 6870
rect 13776 6814 13844 6870
rect 13900 6814 13910 6870
rect 12842 6746 13910 6814
rect 12842 6690 12852 6746
rect 12908 6690 12976 6746
rect 13032 6690 13100 6746
rect 13156 6690 13224 6746
rect 13280 6690 13348 6746
rect 13404 6690 13472 6746
rect 13528 6690 13596 6746
rect 13652 6690 13720 6746
rect 13776 6690 13844 6746
rect 13900 6690 13910 6746
rect 12842 6622 13910 6690
rect 12842 6566 12852 6622
rect 12908 6566 12976 6622
rect 13032 6566 13100 6622
rect 13156 6566 13224 6622
rect 13280 6566 13348 6622
rect 13404 6566 13472 6622
rect 13528 6566 13596 6622
rect 13652 6566 13720 6622
rect 13776 6566 13844 6622
rect 13900 6566 13910 6622
rect 12842 6498 13910 6566
rect 12842 6442 12852 6498
rect 12908 6442 12976 6498
rect 13032 6442 13100 6498
rect 13156 6442 13224 6498
rect 13280 6442 13348 6498
rect 13404 6442 13472 6498
rect 13528 6442 13596 6498
rect 13652 6442 13720 6498
rect 13776 6442 13844 6498
rect 13900 6442 13910 6498
rect 12842 6432 13910 6442
rect 2497 6150 4309 6160
rect 2497 6094 2507 6150
rect 2563 6094 2631 6150
rect 2687 6094 2755 6150
rect 2811 6094 2879 6150
rect 2935 6094 3003 6150
rect 3059 6094 3127 6150
rect 3183 6094 3251 6150
rect 3307 6094 3375 6150
rect 3431 6094 3499 6150
rect 3555 6094 3623 6150
rect 3679 6094 3747 6150
rect 3803 6094 3871 6150
rect 3927 6094 3995 6150
rect 4051 6094 4119 6150
rect 4175 6094 4243 6150
rect 4299 6094 4309 6150
rect 2497 6026 4309 6094
rect 2497 5970 2507 6026
rect 2563 5970 2631 6026
rect 2687 5970 2755 6026
rect 2811 5970 2879 6026
rect 2935 5970 3003 6026
rect 3059 5970 3127 6026
rect 3183 5970 3251 6026
rect 3307 5970 3375 6026
rect 3431 5970 3499 6026
rect 3555 5970 3623 6026
rect 3679 5970 3747 6026
rect 3803 5970 3871 6026
rect 3927 5970 3995 6026
rect 4051 5970 4119 6026
rect 4175 5970 4243 6026
rect 4299 5970 4309 6026
rect 2497 5902 4309 5970
rect 2497 5846 2507 5902
rect 2563 5846 2631 5902
rect 2687 5846 2755 5902
rect 2811 5846 2879 5902
rect 2935 5846 3003 5902
rect 3059 5846 3127 5902
rect 3183 5846 3251 5902
rect 3307 5846 3375 5902
rect 3431 5846 3499 5902
rect 3555 5846 3623 5902
rect 3679 5846 3747 5902
rect 3803 5846 3871 5902
rect 3927 5846 3995 5902
rect 4051 5846 4119 5902
rect 4175 5846 4243 5902
rect 4299 5846 4309 5902
rect 2497 5778 4309 5846
rect 2497 5722 2507 5778
rect 2563 5722 2631 5778
rect 2687 5722 2755 5778
rect 2811 5722 2879 5778
rect 2935 5722 3003 5778
rect 3059 5722 3127 5778
rect 3183 5722 3251 5778
rect 3307 5722 3375 5778
rect 3431 5722 3499 5778
rect 3555 5722 3623 5778
rect 3679 5722 3747 5778
rect 3803 5722 3871 5778
rect 3927 5722 3995 5778
rect 4051 5722 4119 5778
rect 4175 5722 4243 5778
rect 4299 5722 4309 5778
rect 2497 5654 4309 5722
rect 2497 5598 2507 5654
rect 2563 5598 2631 5654
rect 2687 5598 2755 5654
rect 2811 5598 2879 5654
rect 2935 5598 3003 5654
rect 3059 5598 3127 5654
rect 3183 5598 3251 5654
rect 3307 5598 3375 5654
rect 3431 5598 3499 5654
rect 3555 5598 3623 5654
rect 3679 5598 3747 5654
rect 3803 5598 3871 5654
rect 3927 5598 3995 5654
rect 4051 5598 4119 5654
rect 4175 5598 4243 5654
rect 4299 5598 4309 5654
rect 2497 5530 4309 5598
rect 2497 5474 2507 5530
rect 2563 5474 2631 5530
rect 2687 5474 2755 5530
rect 2811 5474 2879 5530
rect 2935 5474 3003 5530
rect 3059 5474 3127 5530
rect 3183 5474 3251 5530
rect 3307 5474 3375 5530
rect 3431 5474 3499 5530
rect 3555 5474 3623 5530
rect 3679 5474 3747 5530
rect 3803 5474 3871 5530
rect 3927 5474 3995 5530
rect 4051 5474 4119 5530
rect 4175 5474 4243 5530
rect 4299 5474 4309 5530
rect 2497 5406 4309 5474
rect 2497 5350 2507 5406
rect 2563 5350 2631 5406
rect 2687 5350 2755 5406
rect 2811 5350 2879 5406
rect 2935 5350 3003 5406
rect 3059 5350 3127 5406
rect 3183 5350 3251 5406
rect 3307 5350 3375 5406
rect 3431 5350 3499 5406
rect 3555 5350 3623 5406
rect 3679 5350 3747 5406
rect 3803 5350 3871 5406
rect 3927 5350 3995 5406
rect 4051 5350 4119 5406
rect 4175 5350 4243 5406
rect 4299 5350 4309 5406
rect 2497 5282 4309 5350
rect 2497 5226 2507 5282
rect 2563 5226 2631 5282
rect 2687 5226 2755 5282
rect 2811 5226 2879 5282
rect 2935 5226 3003 5282
rect 3059 5226 3127 5282
rect 3183 5226 3251 5282
rect 3307 5226 3375 5282
rect 3431 5226 3499 5282
rect 3555 5226 3623 5282
rect 3679 5226 3747 5282
rect 3803 5226 3871 5282
rect 3927 5226 3995 5282
rect 4051 5226 4119 5282
rect 4175 5226 4243 5282
rect 4299 5226 4309 5282
rect 2497 5158 4309 5226
rect 2497 5102 2507 5158
rect 2563 5102 2631 5158
rect 2687 5102 2755 5158
rect 2811 5102 2879 5158
rect 2935 5102 3003 5158
rect 3059 5102 3127 5158
rect 3183 5102 3251 5158
rect 3307 5102 3375 5158
rect 3431 5102 3499 5158
rect 3555 5102 3623 5158
rect 3679 5102 3747 5158
rect 3803 5102 3871 5158
rect 3927 5102 3995 5158
rect 4051 5102 4119 5158
rect 4175 5102 4243 5158
rect 4299 5102 4309 5158
rect 2497 5034 4309 5102
rect 2497 4978 2507 5034
rect 2563 4978 2631 5034
rect 2687 4978 2755 5034
rect 2811 4978 2879 5034
rect 2935 4978 3003 5034
rect 3059 4978 3127 5034
rect 3183 4978 3251 5034
rect 3307 4978 3375 5034
rect 3431 4978 3499 5034
rect 3555 4978 3623 5034
rect 3679 4978 3747 5034
rect 3803 4978 3871 5034
rect 3927 4978 3995 5034
rect 4051 4978 4119 5034
rect 4175 4978 4243 5034
rect 4299 4978 4309 5034
rect 2497 4910 4309 4978
rect 2497 4854 2507 4910
rect 2563 4854 2631 4910
rect 2687 4854 2755 4910
rect 2811 4854 2879 4910
rect 2935 4854 3003 4910
rect 3059 4854 3127 4910
rect 3183 4854 3251 4910
rect 3307 4854 3375 4910
rect 3431 4854 3499 4910
rect 3555 4854 3623 4910
rect 3679 4854 3747 4910
rect 3803 4854 3871 4910
rect 3927 4854 3995 4910
rect 4051 4854 4119 4910
rect 4175 4854 4243 4910
rect 4299 4854 4309 4910
rect 2497 4786 4309 4854
rect 2497 4730 2507 4786
rect 2563 4730 2631 4786
rect 2687 4730 2755 4786
rect 2811 4730 2879 4786
rect 2935 4730 3003 4786
rect 3059 4730 3127 4786
rect 3183 4730 3251 4786
rect 3307 4730 3375 4786
rect 3431 4730 3499 4786
rect 3555 4730 3623 4786
rect 3679 4730 3747 4786
rect 3803 4730 3871 4786
rect 3927 4730 3995 4786
rect 4051 4730 4119 4786
rect 4175 4730 4243 4786
rect 4299 4730 4309 4786
rect 2497 4662 4309 4730
rect 2497 4606 2507 4662
rect 2563 4606 2631 4662
rect 2687 4606 2755 4662
rect 2811 4606 2879 4662
rect 2935 4606 3003 4662
rect 3059 4606 3127 4662
rect 3183 4606 3251 4662
rect 3307 4606 3375 4662
rect 3431 4606 3499 4662
rect 3555 4606 3623 4662
rect 3679 4606 3747 4662
rect 3803 4606 3871 4662
rect 3927 4606 3995 4662
rect 4051 4606 4119 4662
rect 4175 4606 4243 4662
rect 4299 4606 4309 4662
rect 2497 4538 4309 4606
rect 2497 4482 2507 4538
rect 2563 4482 2631 4538
rect 2687 4482 2755 4538
rect 2811 4482 2879 4538
rect 2935 4482 3003 4538
rect 3059 4482 3127 4538
rect 3183 4482 3251 4538
rect 3307 4482 3375 4538
rect 3431 4482 3499 4538
rect 3555 4482 3623 4538
rect 3679 4482 3747 4538
rect 3803 4482 3871 4538
rect 3927 4482 3995 4538
rect 4051 4482 4119 4538
rect 4175 4482 4243 4538
rect 4299 4482 4309 4538
rect 2497 4414 4309 4482
rect 2497 4358 2507 4414
rect 2563 4358 2631 4414
rect 2687 4358 2755 4414
rect 2811 4358 2879 4414
rect 2935 4358 3003 4414
rect 3059 4358 3127 4414
rect 3183 4358 3251 4414
rect 3307 4358 3375 4414
rect 3431 4358 3499 4414
rect 3555 4358 3623 4414
rect 3679 4358 3747 4414
rect 3803 4358 3871 4414
rect 3927 4358 3995 4414
rect 4051 4358 4119 4414
rect 4175 4358 4243 4414
rect 4299 4358 4309 4414
rect 2497 4290 4309 4358
rect 2497 4234 2507 4290
rect 2563 4234 2631 4290
rect 2687 4234 2755 4290
rect 2811 4234 2879 4290
rect 2935 4234 3003 4290
rect 3059 4234 3127 4290
rect 3183 4234 3251 4290
rect 3307 4234 3375 4290
rect 3431 4234 3499 4290
rect 3555 4234 3623 4290
rect 3679 4234 3747 4290
rect 3803 4234 3871 4290
rect 3927 4234 3995 4290
rect 4051 4234 4119 4290
rect 4175 4234 4243 4290
rect 4299 4234 4309 4290
rect 2497 4166 4309 4234
rect 2497 4110 2507 4166
rect 2563 4110 2631 4166
rect 2687 4110 2755 4166
rect 2811 4110 2879 4166
rect 2935 4110 3003 4166
rect 3059 4110 3127 4166
rect 3183 4110 3251 4166
rect 3307 4110 3375 4166
rect 3431 4110 3499 4166
rect 3555 4110 3623 4166
rect 3679 4110 3747 4166
rect 3803 4110 3871 4166
rect 3927 4110 3995 4166
rect 4051 4110 4119 4166
rect 4175 4110 4243 4166
rect 4299 4110 4309 4166
rect 2497 4042 4309 4110
rect 2497 3986 2507 4042
rect 2563 3986 2631 4042
rect 2687 3986 2755 4042
rect 2811 3986 2879 4042
rect 2935 3986 3003 4042
rect 3059 3986 3127 4042
rect 3183 3986 3251 4042
rect 3307 3986 3375 4042
rect 3431 3986 3499 4042
rect 3555 3986 3623 4042
rect 3679 3986 3747 4042
rect 3803 3986 3871 4042
rect 3927 3986 3995 4042
rect 4051 3986 4119 4042
rect 4175 3986 4243 4042
rect 4299 3986 4309 4042
rect 2497 3918 4309 3986
rect 2497 3862 2507 3918
rect 2563 3862 2631 3918
rect 2687 3862 2755 3918
rect 2811 3862 2879 3918
rect 2935 3862 3003 3918
rect 3059 3862 3127 3918
rect 3183 3862 3251 3918
rect 3307 3862 3375 3918
rect 3431 3862 3499 3918
rect 3555 3862 3623 3918
rect 3679 3862 3747 3918
rect 3803 3862 3871 3918
rect 3927 3862 3995 3918
rect 4051 3862 4119 3918
rect 4175 3862 4243 3918
rect 4299 3862 4309 3918
rect 2497 3794 4309 3862
rect 2497 3738 2507 3794
rect 2563 3738 2631 3794
rect 2687 3738 2755 3794
rect 2811 3738 2879 3794
rect 2935 3738 3003 3794
rect 3059 3738 3127 3794
rect 3183 3738 3251 3794
rect 3307 3738 3375 3794
rect 3431 3738 3499 3794
rect 3555 3738 3623 3794
rect 3679 3738 3747 3794
rect 3803 3738 3871 3794
rect 3927 3738 3995 3794
rect 4051 3738 4119 3794
rect 4175 3738 4243 3794
rect 4299 3738 4309 3794
rect 2497 3670 4309 3738
rect 2497 3614 2507 3670
rect 2563 3614 2631 3670
rect 2687 3614 2755 3670
rect 2811 3614 2879 3670
rect 2935 3614 3003 3670
rect 3059 3614 3127 3670
rect 3183 3614 3251 3670
rect 3307 3614 3375 3670
rect 3431 3614 3499 3670
rect 3555 3614 3623 3670
rect 3679 3614 3747 3670
rect 3803 3614 3871 3670
rect 3927 3614 3995 3670
rect 4051 3614 4119 3670
rect 4175 3614 4243 3670
rect 4299 3614 4309 3670
rect 2497 3546 4309 3614
rect 2497 3490 2507 3546
rect 2563 3490 2631 3546
rect 2687 3490 2755 3546
rect 2811 3490 2879 3546
rect 2935 3490 3003 3546
rect 3059 3490 3127 3546
rect 3183 3490 3251 3546
rect 3307 3490 3375 3546
rect 3431 3490 3499 3546
rect 3555 3490 3623 3546
rect 3679 3490 3747 3546
rect 3803 3490 3871 3546
rect 3927 3490 3995 3546
rect 4051 3490 4119 3546
rect 4175 3490 4243 3546
rect 4299 3490 4309 3546
rect 2497 3422 4309 3490
rect 2497 3366 2507 3422
rect 2563 3366 2631 3422
rect 2687 3366 2755 3422
rect 2811 3366 2879 3422
rect 2935 3366 3003 3422
rect 3059 3366 3127 3422
rect 3183 3366 3251 3422
rect 3307 3366 3375 3422
rect 3431 3366 3499 3422
rect 3555 3366 3623 3422
rect 3679 3366 3747 3422
rect 3803 3366 3871 3422
rect 3927 3366 3995 3422
rect 4051 3366 4119 3422
rect 4175 3366 4243 3422
rect 4299 3366 4309 3422
rect 2497 3298 4309 3366
rect 2497 3242 2507 3298
rect 2563 3242 2631 3298
rect 2687 3242 2755 3298
rect 2811 3242 2879 3298
rect 2935 3242 3003 3298
rect 3059 3242 3127 3298
rect 3183 3242 3251 3298
rect 3307 3242 3375 3298
rect 3431 3242 3499 3298
rect 3555 3242 3623 3298
rect 3679 3242 3747 3298
rect 3803 3242 3871 3298
rect 3927 3242 3995 3298
rect 4051 3242 4119 3298
rect 4175 3242 4243 3298
rect 4299 3242 4309 3298
rect 2497 3232 4309 3242
rect 6358 6150 7426 6160
rect 6358 6094 6368 6150
rect 6424 6094 6492 6150
rect 6548 6094 6616 6150
rect 6672 6094 6740 6150
rect 6796 6094 6864 6150
rect 6920 6094 6988 6150
rect 7044 6094 7112 6150
rect 7168 6094 7236 6150
rect 7292 6094 7360 6150
rect 7416 6094 7426 6150
rect 6358 6026 7426 6094
rect 6358 5970 6368 6026
rect 6424 5970 6492 6026
rect 6548 5970 6616 6026
rect 6672 5970 6740 6026
rect 6796 5970 6864 6026
rect 6920 5970 6988 6026
rect 7044 5970 7112 6026
rect 7168 5970 7236 6026
rect 7292 5970 7360 6026
rect 7416 5970 7426 6026
rect 6358 5902 7426 5970
rect 6358 5846 6368 5902
rect 6424 5846 6492 5902
rect 6548 5846 6616 5902
rect 6672 5846 6740 5902
rect 6796 5846 6864 5902
rect 6920 5846 6988 5902
rect 7044 5846 7112 5902
rect 7168 5846 7236 5902
rect 7292 5846 7360 5902
rect 7416 5846 7426 5902
rect 6358 5778 7426 5846
rect 6358 5722 6368 5778
rect 6424 5722 6492 5778
rect 6548 5722 6616 5778
rect 6672 5722 6740 5778
rect 6796 5722 6864 5778
rect 6920 5722 6988 5778
rect 7044 5722 7112 5778
rect 7168 5722 7236 5778
rect 7292 5722 7360 5778
rect 7416 5722 7426 5778
rect 6358 5654 7426 5722
rect 6358 5598 6368 5654
rect 6424 5598 6492 5654
rect 6548 5598 6616 5654
rect 6672 5598 6740 5654
rect 6796 5598 6864 5654
rect 6920 5598 6988 5654
rect 7044 5598 7112 5654
rect 7168 5598 7236 5654
rect 7292 5598 7360 5654
rect 7416 5598 7426 5654
rect 6358 5530 7426 5598
rect 6358 5474 6368 5530
rect 6424 5474 6492 5530
rect 6548 5474 6616 5530
rect 6672 5474 6740 5530
rect 6796 5474 6864 5530
rect 6920 5474 6988 5530
rect 7044 5474 7112 5530
rect 7168 5474 7236 5530
rect 7292 5474 7360 5530
rect 7416 5474 7426 5530
rect 6358 5406 7426 5474
rect 6358 5350 6368 5406
rect 6424 5350 6492 5406
rect 6548 5350 6616 5406
rect 6672 5350 6740 5406
rect 6796 5350 6864 5406
rect 6920 5350 6988 5406
rect 7044 5350 7112 5406
rect 7168 5350 7236 5406
rect 7292 5350 7360 5406
rect 7416 5350 7426 5406
rect 6358 5282 7426 5350
rect 6358 5226 6368 5282
rect 6424 5226 6492 5282
rect 6548 5226 6616 5282
rect 6672 5226 6740 5282
rect 6796 5226 6864 5282
rect 6920 5226 6988 5282
rect 7044 5226 7112 5282
rect 7168 5226 7236 5282
rect 7292 5226 7360 5282
rect 7416 5226 7426 5282
rect 6358 5158 7426 5226
rect 6358 5102 6368 5158
rect 6424 5102 6492 5158
rect 6548 5102 6616 5158
rect 6672 5102 6740 5158
rect 6796 5102 6864 5158
rect 6920 5102 6988 5158
rect 7044 5102 7112 5158
rect 7168 5102 7236 5158
rect 7292 5102 7360 5158
rect 7416 5102 7426 5158
rect 6358 5034 7426 5102
rect 6358 4978 6368 5034
rect 6424 4978 6492 5034
rect 6548 4978 6616 5034
rect 6672 4978 6740 5034
rect 6796 4978 6864 5034
rect 6920 4978 6988 5034
rect 7044 4978 7112 5034
rect 7168 4978 7236 5034
rect 7292 4978 7360 5034
rect 7416 4978 7426 5034
rect 6358 4910 7426 4978
rect 6358 4854 6368 4910
rect 6424 4854 6492 4910
rect 6548 4854 6616 4910
rect 6672 4854 6740 4910
rect 6796 4854 6864 4910
rect 6920 4854 6988 4910
rect 7044 4854 7112 4910
rect 7168 4854 7236 4910
rect 7292 4854 7360 4910
rect 7416 4854 7426 4910
rect 6358 4786 7426 4854
rect 6358 4730 6368 4786
rect 6424 4730 6492 4786
rect 6548 4730 6616 4786
rect 6672 4730 6740 4786
rect 6796 4730 6864 4786
rect 6920 4730 6988 4786
rect 7044 4730 7112 4786
rect 7168 4730 7236 4786
rect 7292 4730 7360 4786
rect 7416 4730 7426 4786
rect 6358 4662 7426 4730
rect 6358 4606 6368 4662
rect 6424 4606 6492 4662
rect 6548 4606 6616 4662
rect 6672 4606 6740 4662
rect 6796 4606 6864 4662
rect 6920 4606 6988 4662
rect 7044 4606 7112 4662
rect 7168 4606 7236 4662
rect 7292 4606 7360 4662
rect 7416 4606 7426 4662
rect 6358 4538 7426 4606
rect 6358 4482 6368 4538
rect 6424 4482 6492 4538
rect 6548 4482 6616 4538
rect 6672 4482 6740 4538
rect 6796 4482 6864 4538
rect 6920 4482 6988 4538
rect 7044 4482 7112 4538
rect 7168 4482 7236 4538
rect 7292 4482 7360 4538
rect 7416 4482 7426 4538
rect 6358 4414 7426 4482
rect 6358 4358 6368 4414
rect 6424 4358 6492 4414
rect 6548 4358 6616 4414
rect 6672 4358 6740 4414
rect 6796 4358 6864 4414
rect 6920 4358 6988 4414
rect 7044 4358 7112 4414
rect 7168 4358 7236 4414
rect 7292 4358 7360 4414
rect 7416 4358 7426 4414
rect 6358 4290 7426 4358
rect 6358 4234 6368 4290
rect 6424 4234 6492 4290
rect 6548 4234 6616 4290
rect 6672 4234 6740 4290
rect 6796 4234 6864 4290
rect 6920 4234 6988 4290
rect 7044 4234 7112 4290
rect 7168 4234 7236 4290
rect 7292 4234 7360 4290
rect 7416 4234 7426 4290
rect 6358 4166 7426 4234
rect 6358 4110 6368 4166
rect 6424 4110 6492 4166
rect 6548 4110 6616 4166
rect 6672 4110 6740 4166
rect 6796 4110 6864 4166
rect 6920 4110 6988 4166
rect 7044 4110 7112 4166
rect 7168 4110 7236 4166
rect 7292 4110 7360 4166
rect 7416 4110 7426 4166
rect 6358 4042 7426 4110
rect 6358 3986 6368 4042
rect 6424 3986 6492 4042
rect 6548 3986 6616 4042
rect 6672 3986 6740 4042
rect 6796 3986 6864 4042
rect 6920 3986 6988 4042
rect 7044 3986 7112 4042
rect 7168 3986 7236 4042
rect 7292 3986 7360 4042
rect 7416 3986 7426 4042
rect 6358 3918 7426 3986
rect 6358 3862 6368 3918
rect 6424 3862 6492 3918
rect 6548 3862 6616 3918
rect 6672 3862 6740 3918
rect 6796 3862 6864 3918
rect 6920 3862 6988 3918
rect 7044 3862 7112 3918
rect 7168 3862 7236 3918
rect 7292 3862 7360 3918
rect 7416 3862 7426 3918
rect 6358 3794 7426 3862
rect 6358 3738 6368 3794
rect 6424 3738 6492 3794
rect 6548 3738 6616 3794
rect 6672 3738 6740 3794
rect 6796 3738 6864 3794
rect 6920 3738 6988 3794
rect 7044 3738 7112 3794
rect 7168 3738 7236 3794
rect 7292 3738 7360 3794
rect 7416 3738 7426 3794
rect 6358 3670 7426 3738
rect 6358 3614 6368 3670
rect 6424 3614 6492 3670
rect 6548 3614 6616 3670
rect 6672 3614 6740 3670
rect 6796 3614 6864 3670
rect 6920 3614 6988 3670
rect 7044 3614 7112 3670
rect 7168 3614 7236 3670
rect 7292 3614 7360 3670
rect 7416 3614 7426 3670
rect 6358 3546 7426 3614
rect 6358 3490 6368 3546
rect 6424 3490 6492 3546
rect 6548 3490 6616 3546
rect 6672 3490 6740 3546
rect 6796 3490 6864 3546
rect 6920 3490 6988 3546
rect 7044 3490 7112 3546
rect 7168 3490 7236 3546
rect 7292 3490 7360 3546
rect 7416 3490 7426 3546
rect 6358 3422 7426 3490
rect 6358 3366 6368 3422
rect 6424 3366 6492 3422
rect 6548 3366 6616 3422
rect 6672 3366 6740 3422
rect 6796 3366 6864 3422
rect 6920 3366 6988 3422
rect 7044 3366 7112 3422
rect 7168 3366 7236 3422
rect 7292 3366 7360 3422
rect 7416 3366 7426 3422
rect 6358 3298 7426 3366
rect 6358 3242 6368 3298
rect 6424 3242 6492 3298
rect 6548 3242 6616 3298
rect 6672 3242 6740 3298
rect 6796 3242 6864 3298
rect 6920 3242 6988 3298
rect 7044 3242 7112 3298
rect 7168 3242 7236 3298
rect 7292 3242 7360 3298
rect 7416 3242 7426 3298
rect 6358 3232 7426 3242
rect 8741 6150 10553 6160
rect 8741 6094 8751 6150
rect 8807 6094 8875 6150
rect 8931 6094 8999 6150
rect 9055 6094 9123 6150
rect 9179 6094 9247 6150
rect 9303 6094 9371 6150
rect 9427 6094 9495 6150
rect 9551 6094 9619 6150
rect 9675 6094 9743 6150
rect 9799 6094 9867 6150
rect 9923 6094 9991 6150
rect 10047 6094 10115 6150
rect 10171 6094 10239 6150
rect 10295 6094 10363 6150
rect 10419 6094 10487 6150
rect 10543 6094 10553 6150
rect 8741 6026 10553 6094
rect 8741 5970 8751 6026
rect 8807 5970 8875 6026
rect 8931 5970 8999 6026
rect 9055 5970 9123 6026
rect 9179 5970 9247 6026
rect 9303 5970 9371 6026
rect 9427 5970 9495 6026
rect 9551 5970 9619 6026
rect 9675 5970 9743 6026
rect 9799 5970 9867 6026
rect 9923 5970 9991 6026
rect 10047 5970 10115 6026
rect 10171 5970 10239 6026
rect 10295 5970 10363 6026
rect 10419 5970 10487 6026
rect 10543 5970 10553 6026
rect 8741 5902 10553 5970
rect 8741 5846 8751 5902
rect 8807 5846 8875 5902
rect 8931 5846 8999 5902
rect 9055 5846 9123 5902
rect 9179 5846 9247 5902
rect 9303 5846 9371 5902
rect 9427 5846 9495 5902
rect 9551 5846 9619 5902
rect 9675 5846 9743 5902
rect 9799 5846 9867 5902
rect 9923 5846 9991 5902
rect 10047 5846 10115 5902
rect 10171 5846 10239 5902
rect 10295 5846 10363 5902
rect 10419 5846 10487 5902
rect 10543 5846 10553 5902
rect 8741 5778 10553 5846
rect 8741 5722 8751 5778
rect 8807 5722 8875 5778
rect 8931 5722 8999 5778
rect 9055 5722 9123 5778
rect 9179 5722 9247 5778
rect 9303 5722 9371 5778
rect 9427 5722 9495 5778
rect 9551 5722 9619 5778
rect 9675 5722 9743 5778
rect 9799 5722 9867 5778
rect 9923 5722 9991 5778
rect 10047 5722 10115 5778
rect 10171 5722 10239 5778
rect 10295 5722 10363 5778
rect 10419 5722 10487 5778
rect 10543 5722 10553 5778
rect 8741 5654 10553 5722
rect 8741 5598 8751 5654
rect 8807 5598 8875 5654
rect 8931 5598 8999 5654
rect 9055 5598 9123 5654
rect 9179 5598 9247 5654
rect 9303 5598 9371 5654
rect 9427 5598 9495 5654
rect 9551 5598 9619 5654
rect 9675 5598 9743 5654
rect 9799 5598 9867 5654
rect 9923 5598 9991 5654
rect 10047 5598 10115 5654
rect 10171 5598 10239 5654
rect 10295 5598 10363 5654
rect 10419 5598 10487 5654
rect 10543 5598 10553 5654
rect 8741 5530 10553 5598
rect 8741 5474 8751 5530
rect 8807 5474 8875 5530
rect 8931 5474 8999 5530
rect 9055 5474 9123 5530
rect 9179 5474 9247 5530
rect 9303 5474 9371 5530
rect 9427 5474 9495 5530
rect 9551 5474 9619 5530
rect 9675 5474 9743 5530
rect 9799 5474 9867 5530
rect 9923 5474 9991 5530
rect 10047 5474 10115 5530
rect 10171 5474 10239 5530
rect 10295 5474 10363 5530
rect 10419 5474 10487 5530
rect 10543 5474 10553 5530
rect 8741 5406 10553 5474
rect 8741 5350 8751 5406
rect 8807 5350 8875 5406
rect 8931 5350 8999 5406
rect 9055 5350 9123 5406
rect 9179 5350 9247 5406
rect 9303 5350 9371 5406
rect 9427 5350 9495 5406
rect 9551 5350 9619 5406
rect 9675 5350 9743 5406
rect 9799 5350 9867 5406
rect 9923 5350 9991 5406
rect 10047 5350 10115 5406
rect 10171 5350 10239 5406
rect 10295 5350 10363 5406
rect 10419 5350 10487 5406
rect 10543 5350 10553 5406
rect 8741 5282 10553 5350
rect 8741 5226 8751 5282
rect 8807 5226 8875 5282
rect 8931 5226 8999 5282
rect 9055 5226 9123 5282
rect 9179 5226 9247 5282
rect 9303 5226 9371 5282
rect 9427 5226 9495 5282
rect 9551 5226 9619 5282
rect 9675 5226 9743 5282
rect 9799 5226 9867 5282
rect 9923 5226 9991 5282
rect 10047 5226 10115 5282
rect 10171 5226 10239 5282
rect 10295 5226 10363 5282
rect 10419 5226 10487 5282
rect 10543 5226 10553 5282
rect 8741 5158 10553 5226
rect 8741 5102 8751 5158
rect 8807 5102 8875 5158
rect 8931 5102 8999 5158
rect 9055 5102 9123 5158
rect 9179 5102 9247 5158
rect 9303 5102 9371 5158
rect 9427 5102 9495 5158
rect 9551 5102 9619 5158
rect 9675 5102 9743 5158
rect 9799 5102 9867 5158
rect 9923 5102 9991 5158
rect 10047 5102 10115 5158
rect 10171 5102 10239 5158
rect 10295 5102 10363 5158
rect 10419 5102 10487 5158
rect 10543 5102 10553 5158
rect 8741 5034 10553 5102
rect 8741 4978 8751 5034
rect 8807 4978 8875 5034
rect 8931 4978 8999 5034
rect 9055 4978 9123 5034
rect 9179 4978 9247 5034
rect 9303 4978 9371 5034
rect 9427 4978 9495 5034
rect 9551 4978 9619 5034
rect 9675 4978 9743 5034
rect 9799 4978 9867 5034
rect 9923 4978 9991 5034
rect 10047 4978 10115 5034
rect 10171 4978 10239 5034
rect 10295 4978 10363 5034
rect 10419 4978 10487 5034
rect 10543 4978 10553 5034
rect 8741 4910 10553 4978
rect 8741 4854 8751 4910
rect 8807 4854 8875 4910
rect 8931 4854 8999 4910
rect 9055 4854 9123 4910
rect 9179 4854 9247 4910
rect 9303 4854 9371 4910
rect 9427 4854 9495 4910
rect 9551 4854 9619 4910
rect 9675 4854 9743 4910
rect 9799 4854 9867 4910
rect 9923 4854 9991 4910
rect 10047 4854 10115 4910
rect 10171 4854 10239 4910
rect 10295 4854 10363 4910
rect 10419 4854 10487 4910
rect 10543 4854 10553 4910
rect 8741 4786 10553 4854
rect 8741 4730 8751 4786
rect 8807 4730 8875 4786
rect 8931 4730 8999 4786
rect 9055 4730 9123 4786
rect 9179 4730 9247 4786
rect 9303 4730 9371 4786
rect 9427 4730 9495 4786
rect 9551 4730 9619 4786
rect 9675 4730 9743 4786
rect 9799 4730 9867 4786
rect 9923 4730 9991 4786
rect 10047 4730 10115 4786
rect 10171 4730 10239 4786
rect 10295 4730 10363 4786
rect 10419 4730 10487 4786
rect 10543 4730 10553 4786
rect 8741 4662 10553 4730
rect 8741 4606 8751 4662
rect 8807 4606 8875 4662
rect 8931 4606 8999 4662
rect 9055 4606 9123 4662
rect 9179 4606 9247 4662
rect 9303 4606 9371 4662
rect 9427 4606 9495 4662
rect 9551 4606 9619 4662
rect 9675 4606 9743 4662
rect 9799 4606 9867 4662
rect 9923 4606 9991 4662
rect 10047 4606 10115 4662
rect 10171 4606 10239 4662
rect 10295 4606 10363 4662
rect 10419 4606 10487 4662
rect 10543 4606 10553 4662
rect 8741 4538 10553 4606
rect 8741 4482 8751 4538
rect 8807 4482 8875 4538
rect 8931 4482 8999 4538
rect 9055 4482 9123 4538
rect 9179 4482 9247 4538
rect 9303 4482 9371 4538
rect 9427 4482 9495 4538
rect 9551 4482 9619 4538
rect 9675 4482 9743 4538
rect 9799 4482 9867 4538
rect 9923 4482 9991 4538
rect 10047 4482 10115 4538
rect 10171 4482 10239 4538
rect 10295 4482 10363 4538
rect 10419 4482 10487 4538
rect 10543 4482 10553 4538
rect 8741 4414 10553 4482
rect 8741 4358 8751 4414
rect 8807 4358 8875 4414
rect 8931 4358 8999 4414
rect 9055 4358 9123 4414
rect 9179 4358 9247 4414
rect 9303 4358 9371 4414
rect 9427 4358 9495 4414
rect 9551 4358 9619 4414
rect 9675 4358 9743 4414
rect 9799 4358 9867 4414
rect 9923 4358 9991 4414
rect 10047 4358 10115 4414
rect 10171 4358 10239 4414
rect 10295 4358 10363 4414
rect 10419 4358 10487 4414
rect 10543 4358 10553 4414
rect 8741 4290 10553 4358
rect 8741 4234 8751 4290
rect 8807 4234 8875 4290
rect 8931 4234 8999 4290
rect 9055 4234 9123 4290
rect 9179 4234 9247 4290
rect 9303 4234 9371 4290
rect 9427 4234 9495 4290
rect 9551 4234 9619 4290
rect 9675 4234 9743 4290
rect 9799 4234 9867 4290
rect 9923 4234 9991 4290
rect 10047 4234 10115 4290
rect 10171 4234 10239 4290
rect 10295 4234 10363 4290
rect 10419 4234 10487 4290
rect 10543 4234 10553 4290
rect 8741 4166 10553 4234
rect 8741 4110 8751 4166
rect 8807 4110 8875 4166
rect 8931 4110 8999 4166
rect 9055 4110 9123 4166
rect 9179 4110 9247 4166
rect 9303 4110 9371 4166
rect 9427 4110 9495 4166
rect 9551 4110 9619 4166
rect 9675 4110 9743 4166
rect 9799 4110 9867 4166
rect 9923 4110 9991 4166
rect 10047 4110 10115 4166
rect 10171 4110 10239 4166
rect 10295 4110 10363 4166
rect 10419 4110 10487 4166
rect 10543 4110 10553 4166
rect 8741 4042 10553 4110
rect 8741 3986 8751 4042
rect 8807 3986 8875 4042
rect 8931 3986 8999 4042
rect 9055 3986 9123 4042
rect 9179 3986 9247 4042
rect 9303 3986 9371 4042
rect 9427 3986 9495 4042
rect 9551 3986 9619 4042
rect 9675 3986 9743 4042
rect 9799 3986 9867 4042
rect 9923 3986 9991 4042
rect 10047 3986 10115 4042
rect 10171 3986 10239 4042
rect 10295 3986 10363 4042
rect 10419 3986 10487 4042
rect 10543 3986 10553 4042
rect 8741 3918 10553 3986
rect 8741 3862 8751 3918
rect 8807 3862 8875 3918
rect 8931 3862 8999 3918
rect 9055 3862 9123 3918
rect 9179 3862 9247 3918
rect 9303 3862 9371 3918
rect 9427 3862 9495 3918
rect 9551 3862 9619 3918
rect 9675 3862 9743 3918
rect 9799 3862 9867 3918
rect 9923 3862 9991 3918
rect 10047 3862 10115 3918
rect 10171 3862 10239 3918
rect 10295 3862 10363 3918
rect 10419 3862 10487 3918
rect 10543 3862 10553 3918
rect 8741 3794 10553 3862
rect 8741 3738 8751 3794
rect 8807 3738 8875 3794
rect 8931 3738 8999 3794
rect 9055 3738 9123 3794
rect 9179 3738 9247 3794
rect 9303 3738 9371 3794
rect 9427 3738 9495 3794
rect 9551 3738 9619 3794
rect 9675 3738 9743 3794
rect 9799 3738 9867 3794
rect 9923 3738 9991 3794
rect 10047 3738 10115 3794
rect 10171 3738 10239 3794
rect 10295 3738 10363 3794
rect 10419 3738 10487 3794
rect 10543 3738 10553 3794
rect 8741 3670 10553 3738
rect 8741 3614 8751 3670
rect 8807 3614 8875 3670
rect 8931 3614 8999 3670
rect 9055 3614 9123 3670
rect 9179 3614 9247 3670
rect 9303 3614 9371 3670
rect 9427 3614 9495 3670
rect 9551 3614 9619 3670
rect 9675 3614 9743 3670
rect 9799 3614 9867 3670
rect 9923 3614 9991 3670
rect 10047 3614 10115 3670
rect 10171 3614 10239 3670
rect 10295 3614 10363 3670
rect 10419 3614 10487 3670
rect 10543 3614 10553 3670
rect 8741 3546 10553 3614
rect 8741 3490 8751 3546
rect 8807 3490 8875 3546
rect 8931 3490 8999 3546
rect 9055 3490 9123 3546
rect 9179 3490 9247 3546
rect 9303 3490 9371 3546
rect 9427 3490 9495 3546
rect 9551 3490 9619 3546
rect 9675 3490 9743 3546
rect 9799 3490 9867 3546
rect 9923 3490 9991 3546
rect 10047 3490 10115 3546
rect 10171 3490 10239 3546
rect 10295 3490 10363 3546
rect 10419 3490 10487 3546
rect 10543 3490 10553 3546
rect 8741 3422 10553 3490
rect 8741 3366 8751 3422
rect 8807 3366 8875 3422
rect 8931 3366 8999 3422
rect 9055 3366 9123 3422
rect 9179 3366 9247 3422
rect 9303 3366 9371 3422
rect 9427 3366 9495 3422
rect 9551 3366 9619 3422
rect 9675 3366 9743 3422
rect 9799 3366 9867 3422
rect 9923 3366 9991 3422
rect 10047 3366 10115 3422
rect 10171 3366 10239 3422
rect 10295 3366 10363 3422
rect 10419 3366 10487 3422
rect 10543 3366 10553 3422
rect 8741 3298 10553 3366
rect 8741 3242 8751 3298
rect 8807 3242 8875 3298
rect 8931 3242 8999 3298
rect 9055 3242 9123 3298
rect 9179 3242 9247 3298
rect 9303 3242 9371 3298
rect 9427 3242 9495 3298
rect 9551 3242 9619 3298
rect 9675 3242 9743 3298
rect 9799 3242 9867 3298
rect 9923 3242 9991 3298
rect 10047 3242 10115 3298
rect 10171 3242 10239 3298
rect 10295 3242 10363 3298
rect 10419 3242 10487 3298
rect 10543 3242 10553 3298
rect 8741 3232 10553 3242
rect 12842 6150 13910 6160
rect 12842 6094 12852 6150
rect 12908 6094 12976 6150
rect 13032 6094 13100 6150
rect 13156 6094 13224 6150
rect 13280 6094 13348 6150
rect 13404 6094 13472 6150
rect 13528 6094 13596 6150
rect 13652 6094 13720 6150
rect 13776 6094 13844 6150
rect 13900 6094 13910 6150
rect 12842 6026 13910 6094
rect 12842 5970 12852 6026
rect 12908 5970 12976 6026
rect 13032 5970 13100 6026
rect 13156 5970 13224 6026
rect 13280 5970 13348 6026
rect 13404 5970 13472 6026
rect 13528 5970 13596 6026
rect 13652 5970 13720 6026
rect 13776 5970 13844 6026
rect 13900 5970 13910 6026
rect 12842 5902 13910 5970
rect 12842 5846 12852 5902
rect 12908 5846 12976 5902
rect 13032 5846 13100 5902
rect 13156 5846 13224 5902
rect 13280 5846 13348 5902
rect 13404 5846 13472 5902
rect 13528 5846 13596 5902
rect 13652 5846 13720 5902
rect 13776 5846 13844 5902
rect 13900 5846 13910 5902
rect 12842 5778 13910 5846
rect 12842 5722 12852 5778
rect 12908 5722 12976 5778
rect 13032 5722 13100 5778
rect 13156 5722 13224 5778
rect 13280 5722 13348 5778
rect 13404 5722 13472 5778
rect 13528 5722 13596 5778
rect 13652 5722 13720 5778
rect 13776 5722 13844 5778
rect 13900 5722 13910 5778
rect 12842 5654 13910 5722
rect 12842 5598 12852 5654
rect 12908 5598 12976 5654
rect 13032 5598 13100 5654
rect 13156 5598 13224 5654
rect 13280 5598 13348 5654
rect 13404 5598 13472 5654
rect 13528 5598 13596 5654
rect 13652 5598 13720 5654
rect 13776 5598 13844 5654
rect 13900 5598 13910 5654
rect 12842 5530 13910 5598
rect 12842 5474 12852 5530
rect 12908 5474 12976 5530
rect 13032 5474 13100 5530
rect 13156 5474 13224 5530
rect 13280 5474 13348 5530
rect 13404 5474 13472 5530
rect 13528 5474 13596 5530
rect 13652 5474 13720 5530
rect 13776 5474 13844 5530
rect 13900 5474 13910 5530
rect 12842 5406 13910 5474
rect 12842 5350 12852 5406
rect 12908 5350 12976 5406
rect 13032 5350 13100 5406
rect 13156 5350 13224 5406
rect 13280 5350 13348 5406
rect 13404 5350 13472 5406
rect 13528 5350 13596 5406
rect 13652 5350 13720 5406
rect 13776 5350 13844 5406
rect 13900 5350 13910 5406
rect 12842 5282 13910 5350
rect 12842 5226 12852 5282
rect 12908 5226 12976 5282
rect 13032 5226 13100 5282
rect 13156 5226 13224 5282
rect 13280 5226 13348 5282
rect 13404 5226 13472 5282
rect 13528 5226 13596 5282
rect 13652 5226 13720 5282
rect 13776 5226 13844 5282
rect 13900 5226 13910 5282
rect 12842 5158 13910 5226
rect 12842 5102 12852 5158
rect 12908 5102 12976 5158
rect 13032 5102 13100 5158
rect 13156 5102 13224 5158
rect 13280 5102 13348 5158
rect 13404 5102 13472 5158
rect 13528 5102 13596 5158
rect 13652 5102 13720 5158
rect 13776 5102 13844 5158
rect 13900 5102 13910 5158
rect 12842 5034 13910 5102
rect 12842 4978 12852 5034
rect 12908 4978 12976 5034
rect 13032 4978 13100 5034
rect 13156 4978 13224 5034
rect 13280 4978 13348 5034
rect 13404 4978 13472 5034
rect 13528 4978 13596 5034
rect 13652 4978 13720 5034
rect 13776 4978 13844 5034
rect 13900 4978 13910 5034
rect 12842 4910 13910 4978
rect 12842 4854 12852 4910
rect 12908 4854 12976 4910
rect 13032 4854 13100 4910
rect 13156 4854 13224 4910
rect 13280 4854 13348 4910
rect 13404 4854 13472 4910
rect 13528 4854 13596 4910
rect 13652 4854 13720 4910
rect 13776 4854 13844 4910
rect 13900 4854 13910 4910
rect 12842 4786 13910 4854
rect 12842 4730 12852 4786
rect 12908 4730 12976 4786
rect 13032 4730 13100 4786
rect 13156 4730 13224 4786
rect 13280 4730 13348 4786
rect 13404 4730 13472 4786
rect 13528 4730 13596 4786
rect 13652 4730 13720 4786
rect 13776 4730 13844 4786
rect 13900 4730 13910 4786
rect 12842 4662 13910 4730
rect 12842 4606 12852 4662
rect 12908 4606 12976 4662
rect 13032 4606 13100 4662
rect 13156 4606 13224 4662
rect 13280 4606 13348 4662
rect 13404 4606 13472 4662
rect 13528 4606 13596 4662
rect 13652 4606 13720 4662
rect 13776 4606 13844 4662
rect 13900 4606 13910 4662
rect 12842 4538 13910 4606
rect 12842 4482 12852 4538
rect 12908 4482 12976 4538
rect 13032 4482 13100 4538
rect 13156 4482 13224 4538
rect 13280 4482 13348 4538
rect 13404 4482 13472 4538
rect 13528 4482 13596 4538
rect 13652 4482 13720 4538
rect 13776 4482 13844 4538
rect 13900 4482 13910 4538
rect 12842 4414 13910 4482
rect 12842 4358 12852 4414
rect 12908 4358 12976 4414
rect 13032 4358 13100 4414
rect 13156 4358 13224 4414
rect 13280 4358 13348 4414
rect 13404 4358 13472 4414
rect 13528 4358 13596 4414
rect 13652 4358 13720 4414
rect 13776 4358 13844 4414
rect 13900 4358 13910 4414
rect 12842 4290 13910 4358
rect 12842 4234 12852 4290
rect 12908 4234 12976 4290
rect 13032 4234 13100 4290
rect 13156 4234 13224 4290
rect 13280 4234 13348 4290
rect 13404 4234 13472 4290
rect 13528 4234 13596 4290
rect 13652 4234 13720 4290
rect 13776 4234 13844 4290
rect 13900 4234 13910 4290
rect 12842 4166 13910 4234
rect 12842 4110 12852 4166
rect 12908 4110 12976 4166
rect 13032 4110 13100 4166
rect 13156 4110 13224 4166
rect 13280 4110 13348 4166
rect 13404 4110 13472 4166
rect 13528 4110 13596 4166
rect 13652 4110 13720 4166
rect 13776 4110 13844 4166
rect 13900 4110 13910 4166
rect 12842 4042 13910 4110
rect 12842 3986 12852 4042
rect 12908 3986 12976 4042
rect 13032 3986 13100 4042
rect 13156 3986 13224 4042
rect 13280 3986 13348 4042
rect 13404 3986 13472 4042
rect 13528 3986 13596 4042
rect 13652 3986 13720 4042
rect 13776 3986 13844 4042
rect 13900 3986 13910 4042
rect 12842 3918 13910 3986
rect 12842 3862 12852 3918
rect 12908 3862 12976 3918
rect 13032 3862 13100 3918
rect 13156 3862 13224 3918
rect 13280 3862 13348 3918
rect 13404 3862 13472 3918
rect 13528 3862 13596 3918
rect 13652 3862 13720 3918
rect 13776 3862 13844 3918
rect 13900 3862 13910 3918
rect 12842 3794 13910 3862
rect 12842 3738 12852 3794
rect 12908 3738 12976 3794
rect 13032 3738 13100 3794
rect 13156 3738 13224 3794
rect 13280 3738 13348 3794
rect 13404 3738 13472 3794
rect 13528 3738 13596 3794
rect 13652 3738 13720 3794
rect 13776 3738 13844 3794
rect 13900 3738 13910 3794
rect 12842 3670 13910 3738
rect 12842 3614 12852 3670
rect 12908 3614 12976 3670
rect 13032 3614 13100 3670
rect 13156 3614 13224 3670
rect 13280 3614 13348 3670
rect 13404 3614 13472 3670
rect 13528 3614 13596 3670
rect 13652 3614 13720 3670
rect 13776 3614 13844 3670
rect 13900 3614 13910 3670
rect 12842 3546 13910 3614
rect 12842 3490 12852 3546
rect 12908 3490 12976 3546
rect 13032 3490 13100 3546
rect 13156 3490 13224 3546
rect 13280 3490 13348 3546
rect 13404 3490 13472 3546
rect 13528 3490 13596 3546
rect 13652 3490 13720 3546
rect 13776 3490 13844 3546
rect 13900 3490 13910 3546
rect 12842 3422 13910 3490
rect 12842 3366 12852 3422
rect 12908 3366 12976 3422
rect 13032 3366 13100 3422
rect 13156 3366 13224 3422
rect 13280 3366 13348 3422
rect 13404 3366 13472 3422
rect 13528 3366 13596 3422
rect 13652 3366 13720 3422
rect 13776 3366 13844 3422
rect 13900 3366 13910 3422
rect 12842 3298 13910 3366
rect 12842 3242 12852 3298
rect 12908 3242 12976 3298
rect 13032 3242 13100 3298
rect 13156 3242 13224 3298
rect 13280 3242 13348 3298
rect 13404 3242 13472 3298
rect 13528 3242 13596 3298
rect 13652 3242 13720 3298
rect 13776 3242 13844 3298
rect 13900 3242 13910 3298
rect 12842 3232 13910 3242
rect 2497 2950 4309 2960
rect 2497 2894 2507 2950
rect 2563 2894 2631 2950
rect 2687 2894 2755 2950
rect 2811 2894 2879 2950
rect 2935 2894 3003 2950
rect 3059 2894 3127 2950
rect 3183 2894 3251 2950
rect 3307 2894 3375 2950
rect 3431 2894 3499 2950
rect 3555 2894 3623 2950
rect 3679 2894 3747 2950
rect 3803 2894 3871 2950
rect 3927 2894 3995 2950
rect 4051 2894 4119 2950
rect 4175 2894 4243 2950
rect 4299 2894 4309 2950
rect 2497 2826 4309 2894
rect 2497 2770 2507 2826
rect 2563 2770 2631 2826
rect 2687 2770 2755 2826
rect 2811 2770 2879 2826
rect 2935 2770 3003 2826
rect 3059 2770 3127 2826
rect 3183 2770 3251 2826
rect 3307 2770 3375 2826
rect 3431 2770 3499 2826
rect 3555 2770 3623 2826
rect 3679 2770 3747 2826
rect 3803 2770 3871 2826
rect 3927 2770 3995 2826
rect 4051 2770 4119 2826
rect 4175 2770 4243 2826
rect 4299 2770 4309 2826
rect 2497 2702 4309 2770
rect 2497 2646 2507 2702
rect 2563 2646 2631 2702
rect 2687 2646 2755 2702
rect 2811 2646 2879 2702
rect 2935 2646 3003 2702
rect 3059 2646 3127 2702
rect 3183 2646 3251 2702
rect 3307 2646 3375 2702
rect 3431 2646 3499 2702
rect 3555 2646 3623 2702
rect 3679 2646 3747 2702
rect 3803 2646 3871 2702
rect 3927 2646 3995 2702
rect 4051 2646 4119 2702
rect 4175 2646 4243 2702
rect 4299 2646 4309 2702
rect 2497 2578 4309 2646
rect 2497 2522 2507 2578
rect 2563 2522 2631 2578
rect 2687 2522 2755 2578
rect 2811 2522 2879 2578
rect 2935 2522 3003 2578
rect 3059 2522 3127 2578
rect 3183 2522 3251 2578
rect 3307 2522 3375 2578
rect 3431 2522 3499 2578
rect 3555 2522 3623 2578
rect 3679 2522 3747 2578
rect 3803 2522 3871 2578
rect 3927 2522 3995 2578
rect 4051 2522 4119 2578
rect 4175 2522 4243 2578
rect 4299 2522 4309 2578
rect 2497 2454 4309 2522
rect 2497 2398 2507 2454
rect 2563 2398 2631 2454
rect 2687 2398 2755 2454
rect 2811 2398 2879 2454
rect 2935 2398 3003 2454
rect 3059 2398 3127 2454
rect 3183 2398 3251 2454
rect 3307 2398 3375 2454
rect 3431 2398 3499 2454
rect 3555 2398 3623 2454
rect 3679 2398 3747 2454
rect 3803 2398 3871 2454
rect 3927 2398 3995 2454
rect 4051 2398 4119 2454
rect 4175 2398 4243 2454
rect 4299 2398 4309 2454
rect 2497 2330 4309 2398
rect 2497 2274 2507 2330
rect 2563 2274 2631 2330
rect 2687 2274 2755 2330
rect 2811 2274 2879 2330
rect 2935 2274 3003 2330
rect 3059 2274 3127 2330
rect 3183 2274 3251 2330
rect 3307 2274 3375 2330
rect 3431 2274 3499 2330
rect 3555 2274 3623 2330
rect 3679 2274 3747 2330
rect 3803 2274 3871 2330
rect 3927 2274 3995 2330
rect 4051 2274 4119 2330
rect 4175 2274 4243 2330
rect 4299 2274 4309 2330
rect 2497 2206 4309 2274
rect 2497 2150 2507 2206
rect 2563 2150 2631 2206
rect 2687 2150 2755 2206
rect 2811 2150 2879 2206
rect 2935 2150 3003 2206
rect 3059 2150 3127 2206
rect 3183 2150 3251 2206
rect 3307 2150 3375 2206
rect 3431 2150 3499 2206
rect 3555 2150 3623 2206
rect 3679 2150 3747 2206
rect 3803 2150 3871 2206
rect 3927 2150 3995 2206
rect 4051 2150 4119 2206
rect 4175 2150 4243 2206
rect 4299 2150 4309 2206
rect 2497 2082 4309 2150
rect 2497 2026 2507 2082
rect 2563 2026 2631 2082
rect 2687 2026 2755 2082
rect 2811 2026 2879 2082
rect 2935 2026 3003 2082
rect 3059 2026 3127 2082
rect 3183 2026 3251 2082
rect 3307 2026 3375 2082
rect 3431 2026 3499 2082
rect 3555 2026 3623 2082
rect 3679 2026 3747 2082
rect 3803 2026 3871 2082
rect 3927 2026 3995 2082
rect 4051 2026 4119 2082
rect 4175 2026 4243 2082
rect 4299 2026 4309 2082
rect 2497 1958 4309 2026
rect 2497 1902 2507 1958
rect 2563 1902 2631 1958
rect 2687 1902 2755 1958
rect 2811 1902 2879 1958
rect 2935 1902 3003 1958
rect 3059 1902 3127 1958
rect 3183 1902 3251 1958
rect 3307 1902 3375 1958
rect 3431 1902 3499 1958
rect 3555 1902 3623 1958
rect 3679 1902 3747 1958
rect 3803 1902 3871 1958
rect 3927 1902 3995 1958
rect 4051 1902 4119 1958
rect 4175 1902 4243 1958
rect 4299 1902 4309 1958
rect 2497 1834 4309 1902
rect 2497 1778 2507 1834
rect 2563 1778 2631 1834
rect 2687 1778 2755 1834
rect 2811 1778 2879 1834
rect 2935 1778 3003 1834
rect 3059 1778 3127 1834
rect 3183 1778 3251 1834
rect 3307 1778 3375 1834
rect 3431 1778 3499 1834
rect 3555 1778 3623 1834
rect 3679 1778 3747 1834
rect 3803 1778 3871 1834
rect 3927 1778 3995 1834
rect 4051 1778 4119 1834
rect 4175 1778 4243 1834
rect 4299 1778 4309 1834
rect 2497 1710 4309 1778
rect 2497 1654 2507 1710
rect 2563 1654 2631 1710
rect 2687 1654 2755 1710
rect 2811 1654 2879 1710
rect 2935 1654 3003 1710
rect 3059 1654 3127 1710
rect 3183 1654 3251 1710
rect 3307 1654 3375 1710
rect 3431 1654 3499 1710
rect 3555 1654 3623 1710
rect 3679 1654 3747 1710
rect 3803 1654 3871 1710
rect 3927 1654 3995 1710
rect 4051 1654 4119 1710
rect 4175 1654 4243 1710
rect 4299 1654 4309 1710
rect 2497 1586 4309 1654
rect 2497 1530 2507 1586
rect 2563 1530 2631 1586
rect 2687 1530 2755 1586
rect 2811 1530 2879 1586
rect 2935 1530 3003 1586
rect 3059 1530 3127 1586
rect 3183 1530 3251 1586
rect 3307 1530 3375 1586
rect 3431 1530 3499 1586
rect 3555 1530 3623 1586
rect 3679 1530 3747 1586
rect 3803 1530 3871 1586
rect 3927 1530 3995 1586
rect 4051 1530 4119 1586
rect 4175 1530 4243 1586
rect 4299 1530 4309 1586
rect 2497 1462 4309 1530
rect 2497 1406 2507 1462
rect 2563 1406 2631 1462
rect 2687 1406 2755 1462
rect 2811 1406 2879 1462
rect 2935 1406 3003 1462
rect 3059 1406 3127 1462
rect 3183 1406 3251 1462
rect 3307 1406 3375 1462
rect 3431 1406 3499 1462
rect 3555 1406 3623 1462
rect 3679 1406 3747 1462
rect 3803 1406 3871 1462
rect 3927 1406 3995 1462
rect 4051 1406 4119 1462
rect 4175 1406 4243 1462
rect 4299 1406 4309 1462
rect 2497 1338 4309 1406
rect 2497 1282 2507 1338
rect 2563 1282 2631 1338
rect 2687 1282 2755 1338
rect 2811 1282 2879 1338
rect 2935 1282 3003 1338
rect 3059 1282 3127 1338
rect 3183 1282 3251 1338
rect 3307 1282 3375 1338
rect 3431 1282 3499 1338
rect 3555 1282 3623 1338
rect 3679 1282 3747 1338
rect 3803 1282 3871 1338
rect 3927 1282 3995 1338
rect 4051 1282 4119 1338
rect 4175 1282 4243 1338
rect 4299 1282 4309 1338
rect 2497 1214 4309 1282
rect 2497 1158 2507 1214
rect 2563 1158 2631 1214
rect 2687 1158 2755 1214
rect 2811 1158 2879 1214
rect 2935 1158 3003 1214
rect 3059 1158 3127 1214
rect 3183 1158 3251 1214
rect 3307 1158 3375 1214
rect 3431 1158 3499 1214
rect 3555 1158 3623 1214
rect 3679 1158 3747 1214
rect 3803 1158 3871 1214
rect 3927 1158 3995 1214
rect 4051 1158 4119 1214
rect 4175 1158 4243 1214
rect 4299 1158 4309 1214
rect 2497 1090 4309 1158
rect 2497 1034 2507 1090
rect 2563 1034 2631 1090
rect 2687 1034 2755 1090
rect 2811 1034 2879 1090
rect 2935 1034 3003 1090
rect 3059 1034 3127 1090
rect 3183 1034 3251 1090
rect 3307 1034 3375 1090
rect 3431 1034 3499 1090
rect 3555 1034 3623 1090
rect 3679 1034 3747 1090
rect 3803 1034 3871 1090
rect 3927 1034 3995 1090
rect 4051 1034 4119 1090
rect 4175 1034 4243 1090
rect 4299 1034 4309 1090
rect 2497 966 4309 1034
rect 2497 910 2507 966
rect 2563 910 2631 966
rect 2687 910 2755 966
rect 2811 910 2879 966
rect 2935 910 3003 966
rect 3059 910 3127 966
rect 3183 910 3251 966
rect 3307 910 3375 966
rect 3431 910 3499 966
rect 3555 910 3623 966
rect 3679 910 3747 966
rect 3803 910 3871 966
rect 3927 910 3995 966
rect 4051 910 4119 966
rect 4175 910 4243 966
rect 4299 910 4309 966
rect 2497 842 4309 910
rect 2497 786 2507 842
rect 2563 786 2631 842
rect 2687 786 2755 842
rect 2811 786 2879 842
rect 2935 786 3003 842
rect 3059 786 3127 842
rect 3183 786 3251 842
rect 3307 786 3375 842
rect 3431 786 3499 842
rect 3555 786 3623 842
rect 3679 786 3747 842
rect 3803 786 3871 842
rect 3927 786 3995 842
rect 4051 786 4119 842
rect 4175 786 4243 842
rect 4299 786 4309 842
rect 2497 718 4309 786
rect 2497 662 2507 718
rect 2563 662 2631 718
rect 2687 662 2755 718
rect 2811 662 2879 718
rect 2935 662 3003 718
rect 3059 662 3127 718
rect 3183 662 3251 718
rect 3307 662 3375 718
rect 3431 662 3499 718
rect 3555 662 3623 718
rect 3679 662 3747 718
rect 3803 662 3871 718
rect 3927 662 3995 718
rect 4051 662 4119 718
rect 4175 662 4243 718
rect 4299 662 4309 718
rect 2497 594 4309 662
rect 2497 538 2507 594
rect 2563 538 2631 594
rect 2687 538 2755 594
rect 2811 538 2879 594
rect 2935 538 3003 594
rect 3059 538 3127 594
rect 3183 538 3251 594
rect 3307 538 3375 594
rect 3431 538 3499 594
rect 3555 538 3623 594
rect 3679 538 3747 594
rect 3803 538 3871 594
rect 3927 538 3995 594
rect 4051 538 4119 594
rect 4175 538 4243 594
rect 4299 538 4309 594
rect 2497 470 4309 538
rect 2497 414 2507 470
rect 2563 414 2631 470
rect 2687 414 2755 470
rect 2811 414 2879 470
rect 2935 414 3003 470
rect 3059 414 3127 470
rect 3183 414 3251 470
rect 3307 414 3375 470
rect 3431 414 3499 470
rect 3555 414 3623 470
rect 3679 414 3747 470
rect 3803 414 3871 470
rect 3927 414 3995 470
rect 4051 414 4119 470
rect 4175 414 4243 470
rect 4299 414 4309 470
rect 2497 346 4309 414
rect 2497 290 2507 346
rect 2563 290 2631 346
rect 2687 290 2755 346
rect 2811 290 2879 346
rect 2935 290 3003 346
rect 3059 290 3127 346
rect 3183 290 3251 346
rect 3307 290 3375 346
rect 3431 290 3499 346
rect 3555 290 3623 346
rect 3679 290 3747 346
rect 3803 290 3871 346
rect 3927 290 3995 346
rect 4051 290 4119 346
rect 4175 290 4243 346
rect 4299 290 4309 346
rect 2497 222 4309 290
rect 2497 166 2507 222
rect 2563 166 2631 222
rect 2687 166 2755 222
rect 2811 166 2879 222
rect 2935 166 3003 222
rect 3059 166 3127 222
rect 3183 166 3251 222
rect 3307 166 3375 222
rect 3431 166 3499 222
rect 3555 166 3623 222
rect 3679 166 3747 222
rect 3803 166 3871 222
rect 3927 166 3995 222
rect 4051 166 4119 222
rect 4175 166 4243 222
rect 4299 166 4309 222
rect 2497 98 4309 166
rect 2497 42 2507 98
rect 2563 42 2631 98
rect 2687 42 2755 98
rect 2811 42 2879 98
rect 2935 42 3003 98
rect 3059 42 3127 98
rect 3183 42 3251 98
rect 3307 42 3375 98
rect 3431 42 3499 98
rect 3555 42 3623 98
rect 3679 42 3747 98
rect 3803 42 3871 98
rect 3927 42 3995 98
rect 4051 42 4119 98
rect 4175 42 4243 98
rect 4299 42 4309 98
rect 2497 32 4309 42
rect 6358 2950 7426 2960
rect 6358 2894 6368 2950
rect 6424 2894 6492 2950
rect 6548 2894 6616 2950
rect 6672 2894 6740 2950
rect 6796 2894 6864 2950
rect 6920 2894 6988 2950
rect 7044 2894 7112 2950
rect 7168 2894 7236 2950
rect 7292 2894 7360 2950
rect 7416 2894 7426 2950
rect 6358 2826 7426 2894
rect 6358 2770 6368 2826
rect 6424 2770 6492 2826
rect 6548 2770 6616 2826
rect 6672 2770 6740 2826
rect 6796 2770 6864 2826
rect 6920 2770 6988 2826
rect 7044 2770 7112 2826
rect 7168 2770 7236 2826
rect 7292 2770 7360 2826
rect 7416 2770 7426 2826
rect 6358 2702 7426 2770
rect 6358 2646 6368 2702
rect 6424 2646 6492 2702
rect 6548 2646 6616 2702
rect 6672 2646 6740 2702
rect 6796 2646 6864 2702
rect 6920 2646 6988 2702
rect 7044 2646 7112 2702
rect 7168 2646 7236 2702
rect 7292 2646 7360 2702
rect 7416 2646 7426 2702
rect 6358 2578 7426 2646
rect 6358 2522 6368 2578
rect 6424 2522 6492 2578
rect 6548 2522 6616 2578
rect 6672 2522 6740 2578
rect 6796 2522 6864 2578
rect 6920 2522 6988 2578
rect 7044 2522 7112 2578
rect 7168 2522 7236 2578
rect 7292 2522 7360 2578
rect 7416 2522 7426 2578
rect 6358 2454 7426 2522
rect 6358 2398 6368 2454
rect 6424 2398 6492 2454
rect 6548 2398 6616 2454
rect 6672 2398 6740 2454
rect 6796 2398 6864 2454
rect 6920 2398 6988 2454
rect 7044 2398 7112 2454
rect 7168 2398 7236 2454
rect 7292 2398 7360 2454
rect 7416 2398 7426 2454
rect 6358 2330 7426 2398
rect 6358 2274 6368 2330
rect 6424 2274 6492 2330
rect 6548 2274 6616 2330
rect 6672 2274 6740 2330
rect 6796 2274 6864 2330
rect 6920 2274 6988 2330
rect 7044 2274 7112 2330
rect 7168 2274 7236 2330
rect 7292 2274 7360 2330
rect 7416 2274 7426 2330
rect 6358 2206 7426 2274
rect 6358 2150 6368 2206
rect 6424 2150 6492 2206
rect 6548 2150 6616 2206
rect 6672 2150 6740 2206
rect 6796 2150 6864 2206
rect 6920 2150 6988 2206
rect 7044 2150 7112 2206
rect 7168 2150 7236 2206
rect 7292 2150 7360 2206
rect 7416 2150 7426 2206
rect 6358 2082 7426 2150
rect 6358 2026 6368 2082
rect 6424 2026 6492 2082
rect 6548 2026 6616 2082
rect 6672 2026 6740 2082
rect 6796 2026 6864 2082
rect 6920 2026 6988 2082
rect 7044 2026 7112 2082
rect 7168 2026 7236 2082
rect 7292 2026 7360 2082
rect 7416 2026 7426 2082
rect 6358 1958 7426 2026
rect 6358 1902 6368 1958
rect 6424 1902 6492 1958
rect 6548 1902 6616 1958
rect 6672 1902 6740 1958
rect 6796 1902 6864 1958
rect 6920 1902 6988 1958
rect 7044 1902 7112 1958
rect 7168 1902 7236 1958
rect 7292 1902 7360 1958
rect 7416 1902 7426 1958
rect 6358 1834 7426 1902
rect 6358 1778 6368 1834
rect 6424 1778 6492 1834
rect 6548 1778 6616 1834
rect 6672 1778 6740 1834
rect 6796 1778 6864 1834
rect 6920 1778 6988 1834
rect 7044 1778 7112 1834
rect 7168 1778 7236 1834
rect 7292 1778 7360 1834
rect 7416 1778 7426 1834
rect 6358 1710 7426 1778
rect 6358 1654 6368 1710
rect 6424 1654 6492 1710
rect 6548 1654 6616 1710
rect 6672 1654 6740 1710
rect 6796 1654 6864 1710
rect 6920 1654 6988 1710
rect 7044 1654 7112 1710
rect 7168 1654 7236 1710
rect 7292 1654 7360 1710
rect 7416 1654 7426 1710
rect 6358 1586 7426 1654
rect 6358 1530 6368 1586
rect 6424 1530 6492 1586
rect 6548 1530 6616 1586
rect 6672 1530 6740 1586
rect 6796 1530 6864 1586
rect 6920 1530 6988 1586
rect 7044 1530 7112 1586
rect 7168 1530 7236 1586
rect 7292 1530 7360 1586
rect 7416 1530 7426 1586
rect 6358 1462 7426 1530
rect 6358 1406 6368 1462
rect 6424 1406 6492 1462
rect 6548 1406 6616 1462
rect 6672 1406 6740 1462
rect 6796 1406 6864 1462
rect 6920 1406 6988 1462
rect 7044 1406 7112 1462
rect 7168 1406 7236 1462
rect 7292 1406 7360 1462
rect 7416 1406 7426 1462
rect 6358 1338 7426 1406
rect 6358 1282 6368 1338
rect 6424 1282 6492 1338
rect 6548 1282 6616 1338
rect 6672 1282 6740 1338
rect 6796 1282 6864 1338
rect 6920 1282 6988 1338
rect 7044 1282 7112 1338
rect 7168 1282 7236 1338
rect 7292 1282 7360 1338
rect 7416 1282 7426 1338
rect 6358 1214 7426 1282
rect 6358 1158 6368 1214
rect 6424 1158 6492 1214
rect 6548 1158 6616 1214
rect 6672 1158 6740 1214
rect 6796 1158 6864 1214
rect 6920 1158 6988 1214
rect 7044 1158 7112 1214
rect 7168 1158 7236 1214
rect 7292 1158 7360 1214
rect 7416 1158 7426 1214
rect 6358 1090 7426 1158
rect 6358 1034 6368 1090
rect 6424 1034 6492 1090
rect 6548 1034 6616 1090
rect 6672 1034 6740 1090
rect 6796 1034 6864 1090
rect 6920 1034 6988 1090
rect 7044 1034 7112 1090
rect 7168 1034 7236 1090
rect 7292 1034 7360 1090
rect 7416 1034 7426 1090
rect 6358 966 7426 1034
rect 6358 910 6368 966
rect 6424 910 6492 966
rect 6548 910 6616 966
rect 6672 910 6740 966
rect 6796 910 6864 966
rect 6920 910 6988 966
rect 7044 910 7112 966
rect 7168 910 7236 966
rect 7292 910 7360 966
rect 7416 910 7426 966
rect 6358 842 7426 910
rect 6358 786 6368 842
rect 6424 786 6492 842
rect 6548 786 6616 842
rect 6672 786 6740 842
rect 6796 786 6864 842
rect 6920 786 6988 842
rect 7044 786 7112 842
rect 7168 786 7236 842
rect 7292 786 7360 842
rect 7416 786 7426 842
rect 6358 718 7426 786
rect 6358 662 6368 718
rect 6424 662 6492 718
rect 6548 662 6616 718
rect 6672 662 6740 718
rect 6796 662 6864 718
rect 6920 662 6988 718
rect 7044 662 7112 718
rect 7168 662 7236 718
rect 7292 662 7360 718
rect 7416 662 7426 718
rect 6358 594 7426 662
rect 6358 538 6368 594
rect 6424 538 6492 594
rect 6548 538 6616 594
rect 6672 538 6740 594
rect 6796 538 6864 594
rect 6920 538 6988 594
rect 7044 538 7112 594
rect 7168 538 7236 594
rect 7292 538 7360 594
rect 7416 538 7426 594
rect 6358 470 7426 538
rect 6358 414 6368 470
rect 6424 414 6492 470
rect 6548 414 6616 470
rect 6672 414 6740 470
rect 6796 414 6864 470
rect 6920 414 6988 470
rect 7044 414 7112 470
rect 7168 414 7236 470
rect 7292 414 7360 470
rect 7416 414 7426 470
rect 6358 346 7426 414
rect 6358 290 6368 346
rect 6424 290 6492 346
rect 6548 290 6616 346
rect 6672 290 6740 346
rect 6796 290 6864 346
rect 6920 290 6988 346
rect 7044 290 7112 346
rect 7168 290 7236 346
rect 7292 290 7360 346
rect 7416 290 7426 346
rect 6358 222 7426 290
rect 6358 166 6368 222
rect 6424 166 6492 222
rect 6548 166 6616 222
rect 6672 166 6740 222
rect 6796 166 6864 222
rect 6920 166 6988 222
rect 7044 166 7112 222
rect 7168 166 7236 222
rect 7292 166 7360 222
rect 7416 166 7426 222
rect 6358 98 7426 166
rect 6358 42 6368 98
rect 6424 42 6492 98
rect 6548 42 6616 98
rect 6672 42 6740 98
rect 6796 42 6864 98
rect 6920 42 6988 98
rect 7044 42 7112 98
rect 7168 42 7236 98
rect 7292 42 7360 98
rect 7416 42 7426 98
rect 6358 32 7426 42
rect 8741 2950 10553 2960
rect 8741 2894 8751 2950
rect 8807 2894 8875 2950
rect 8931 2894 8999 2950
rect 9055 2894 9123 2950
rect 9179 2894 9247 2950
rect 9303 2894 9371 2950
rect 9427 2894 9495 2950
rect 9551 2894 9619 2950
rect 9675 2894 9743 2950
rect 9799 2894 9867 2950
rect 9923 2894 9991 2950
rect 10047 2894 10115 2950
rect 10171 2894 10239 2950
rect 10295 2894 10363 2950
rect 10419 2894 10487 2950
rect 10543 2894 10553 2950
rect 8741 2826 10553 2894
rect 8741 2770 8751 2826
rect 8807 2770 8875 2826
rect 8931 2770 8999 2826
rect 9055 2770 9123 2826
rect 9179 2770 9247 2826
rect 9303 2770 9371 2826
rect 9427 2770 9495 2826
rect 9551 2770 9619 2826
rect 9675 2770 9743 2826
rect 9799 2770 9867 2826
rect 9923 2770 9991 2826
rect 10047 2770 10115 2826
rect 10171 2770 10239 2826
rect 10295 2770 10363 2826
rect 10419 2770 10487 2826
rect 10543 2770 10553 2826
rect 8741 2702 10553 2770
rect 8741 2646 8751 2702
rect 8807 2646 8875 2702
rect 8931 2646 8999 2702
rect 9055 2646 9123 2702
rect 9179 2646 9247 2702
rect 9303 2646 9371 2702
rect 9427 2646 9495 2702
rect 9551 2646 9619 2702
rect 9675 2646 9743 2702
rect 9799 2646 9867 2702
rect 9923 2646 9991 2702
rect 10047 2646 10115 2702
rect 10171 2646 10239 2702
rect 10295 2646 10363 2702
rect 10419 2646 10487 2702
rect 10543 2646 10553 2702
rect 8741 2578 10553 2646
rect 8741 2522 8751 2578
rect 8807 2522 8875 2578
rect 8931 2522 8999 2578
rect 9055 2522 9123 2578
rect 9179 2522 9247 2578
rect 9303 2522 9371 2578
rect 9427 2522 9495 2578
rect 9551 2522 9619 2578
rect 9675 2522 9743 2578
rect 9799 2522 9867 2578
rect 9923 2522 9991 2578
rect 10047 2522 10115 2578
rect 10171 2522 10239 2578
rect 10295 2522 10363 2578
rect 10419 2522 10487 2578
rect 10543 2522 10553 2578
rect 8741 2454 10553 2522
rect 8741 2398 8751 2454
rect 8807 2398 8875 2454
rect 8931 2398 8999 2454
rect 9055 2398 9123 2454
rect 9179 2398 9247 2454
rect 9303 2398 9371 2454
rect 9427 2398 9495 2454
rect 9551 2398 9619 2454
rect 9675 2398 9743 2454
rect 9799 2398 9867 2454
rect 9923 2398 9991 2454
rect 10047 2398 10115 2454
rect 10171 2398 10239 2454
rect 10295 2398 10363 2454
rect 10419 2398 10487 2454
rect 10543 2398 10553 2454
rect 8741 2330 10553 2398
rect 8741 2274 8751 2330
rect 8807 2274 8875 2330
rect 8931 2274 8999 2330
rect 9055 2274 9123 2330
rect 9179 2274 9247 2330
rect 9303 2274 9371 2330
rect 9427 2274 9495 2330
rect 9551 2274 9619 2330
rect 9675 2274 9743 2330
rect 9799 2274 9867 2330
rect 9923 2274 9991 2330
rect 10047 2274 10115 2330
rect 10171 2274 10239 2330
rect 10295 2274 10363 2330
rect 10419 2274 10487 2330
rect 10543 2274 10553 2330
rect 8741 2206 10553 2274
rect 8741 2150 8751 2206
rect 8807 2150 8875 2206
rect 8931 2150 8999 2206
rect 9055 2150 9123 2206
rect 9179 2150 9247 2206
rect 9303 2150 9371 2206
rect 9427 2150 9495 2206
rect 9551 2150 9619 2206
rect 9675 2150 9743 2206
rect 9799 2150 9867 2206
rect 9923 2150 9991 2206
rect 10047 2150 10115 2206
rect 10171 2150 10239 2206
rect 10295 2150 10363 2206
rect 10419 2150 10487 2206
rect 10543 2150 10553 2206
rect 8741 2082 10553 2150
rect 8741 2026 8751 2082
rect 8807 2026 8875 2082
rect 8931 2026 8999 2082
rect 9055 2026 9123 2082
rect 9179 2026 9247 2082
rect 9303 2026 9371 2082
rect 9427 2026 9495 2082
rect 9551 2026 9619 2082
rect 9675 2026 9743 2082
rect 9799 2026 9867 2082
rect 9923 2026 9991 2082
rect 10047 2026 10115 2082
rect 10171 2026 10239 2082
rect 10295 2026 10363 2082
rect 10419 2026 10487 2082
rect 10543 2026 10553 2082
rect 8741 1958 10553 2026
rect 8741 1902 8751 1958
rect 8807 1902 8875 1958
rect 8931 1902 8999 1958
rect 9055 1902 9123 1958
rect 9179 1902 9247 1958
rect 9303 1902 9371 1958
rect 9427 1902 9495 1958
rect 9551 1902 9619 1958
rect 9675 1902 9743 1958
rect 9799 1902 9867 1958
rect 9923 1902 9991 1958
rect 10047 1902 10115 1958
rect 10171 1902 10239 1958
rect 10295 1902 10363 1958
rect 10419 1902 10487 1958
rect 10543 1902 10553 1958
rect 8741 1834 10553 1902
rect 8741 1778 8751 1834
rect 8807 1778 8875 1834
rect 8931 1778 8999 1834
rect 9055 1778 9123 1834
rect 9179 1778 9247 1834
rect 9303 1778 9371 1834
rect 9427 1778 9495 1834
rect 9551 1778 9619 1834
rect 9675 1778 9743 1834
rect 9799 1778 9867 1834
rect 9923 1778 9991 1834
rect 10047 1778 10115 1834
rect 10171 1778 10239 1834
rect 10295 1778 10363 1834
rect 10419 1778 10487 1834
rect 10543 1778 10553 1834
rect 8741 1710 10553 1778
rect 8741 1654 8751 1710
rect 8807 1654 8875 1710
rect 8931 1654 8999 1710
rect 9055 1654 9123 1710
rect 9179 1654 9247 1710
rect 9303 1654 9371 1710
rect 9427 1654 9495 1710
rect 9551 1654 9619 1710
rect 9675 1654 9743 1710
rect 9799 1654 9867 1710
rect 9923 1654 9991 1710
rect 10047 1654 10115 1710
rect 10171 1654 10239 1710
rect 10295 1654 10363 1710
rect 10419 1654 10487 1710
rect 10543 1654 10553 1710
rect 8741 1586 10553 1654
rect 8741 1530 8751 1586
rect 8807 1530 8875 1586
rect 8931 1530 8999 1586
rect 9055 1530 9123 1586
rect 9179 1530 9247 1586
rect 9303 1530 9371 1586
rect 9427 1530 9495 1586
rect 9551 1530 9619 1586
rect 9675 1530 9743 1586
rect 9799 1530 9867 1586
rect 9923 1530 9991 1586
rect 10047 1530 10115 1586
rect 10171 1530 10239 1586
rect 10295 1530 10363 1586
rect 10419 1530 10487 1586
rect 10543 1530 10553 1586
rect 8741 1462 10553 1530
rect 8741 1406 8751 1462
rect 8807 1406 8875 1462
rect 8931 1406 8999 1462
rect 9055 1406 9123 1462
rect 9179 1406 9247 1462
rect 9303 1406 9371 1462
rect 9427 1406 9495 1462
rect 9551 1406 9619 1462
rect 9675 1406 9743 1462
rect 9799 1406 9867 1462
rect 9923 1406 9991 1462
rect 10047 1406 10115 1462
rect 10171 1406 10239 1462
rect 10295 1406 10363 1462
rect 10419 1406 10487 1462
rect 10543 1406 10553 1462
rect 8741 1338 10553 1406
rect 8741 1282 8751 1338
rect 8807 1282 8875 1338
rect 8931 1282 8999 1338
rect 9055 1282 9123 1338
rect 9179 1282 9247 1338
rect 9303 1282 9371 1338
rect 9427 1282 9495 1338
rect 9551 1282 9619 1338
rect 9675 1282 9743 1338
rect 9799 1282 9867 1338
rect 9923 1282 9991 1338
rect 10047 1282 10115 1338
rect 10171 1282 10239 1338
rect 10295 1282 10363 1338
rect 10419 1282 10487 1338
rect 10543 1282 10553 1338
rect 8741 1214 10553 1282
rect 8741 1158 8751 1214
rect 8807 1158 8875 1214
rect 8931 1158 8999 1214
rect 9055 1158 9123 1214
rect 9179 1158 9247 1214
rect 9303 1158 9371 1214
rect 9427 1158 9495 1214
rect 9551 1158 9619 1214
rect 9675 1158 9743 1214
rect 9799 1158 9867 1214
rect 9923 1158 9991 1214
rect 10047 1158 10115 1214
rect 10171 1158 10239 1214
rect 10295 1158 10363 1214
rect 10419 1158 10487 1214
rect 10543 1158 10553 1214
rect 8741 1090 10553 1158
rect 8741 1034 8751 1090
rect 8807 1034 8875 1090
rect 8931 1034 8999 1090
rect 9055 1034 9123 1090
rect 9179 1034 9247 1090
rect 9303 1034 9371 1090
rect 9427 1034 9495 1090
rect 9551 1034 9619 1090
rect 9675 1034 9743 1090
rect 9799 1034 9867 1090
rect 9923 1034 9991 1090
rect 10047 1034 10115 1090
rect 10171 1034 10239 1090
rect 10295 1034 10363 1090
rect 10419 1034 10487 1090
rect 10543 1034 10553 1090
rect 8741 966 10553 1034
rect 8741 910 8751 966
rect 8807 910 8875 966
rect 8931 910 8999 966
rect 9055 910 9123 966
rect 9179 910 9247 966
rect 9303 910 9371 966
rect 9427 910 9495 966
rect 9551 910 9619 966
rect 9675 910 9743 966
rect 9799 910 9867 966
rect 9923 910 9991 966
rect 10047 910 10115 966
rect 10171 910 10239 966
rect 10295 910 10363 966
rect 10419 910 10487 966
rect 10543 910 10553 966
rect 8741 842 10553 910
rect 8741 786 8751 842
rect 8807 786 8875 842
rect 8931 786 8999 842
rect 9055 786 9123 842
rect 9179 786 9247 842
rect 9303 786 9371 842
rect 9427 786 9495 842
rect 9551 786 9619 842
rect 9675 786 9743 842
rect 9799 786 9867 842
rect 9923 786 9991 842
rect 10047 786 10115 842
rect 10171 786 10239 842
rect 10295 786 10363 842
rect 10419 786 10487 842
rect 10543 786 10553 842
rect 8741 718 10553 786
rect 8741 662 8751 718
rect 8807 662 8875 718
rect 8931 662 8999 718
rect 9055 662 9123 718
rect 9179 662 9247 718
rect 9303 662 9371 718
rect 9427 662 9495 718
rect 9551 662 9619 718
rect 9675 662 9743 718
rect 9799 662 9867 718
rect 9923 662 9991 718
rect 10047 662 10115 718
rect 10171 662 10239 718
rect 10295 662 10363 718
rect 10419 662 10487 718
rect 10543 662 10553 718
rect 8741 594 10553 662
rect 8741 538 8751 594
rect 8807 538 8875 594
rect 8931 538 8999 594
rect 9055 538 9123 594
rect 9179 538 9247 594
rect 9303 538 9371 594
rect 9427 538 9495 594
rect 9551 538 9619 594
rect 9675 538 9743 594
rect 9799 538 9867 594
rect 9923 538 9991 594
rect 10047 538 10115 594
rect 10171 538 10239 594
rect 10295 538 10363 594
rect 10419 538 10487 594
rect 10543 538 10553 594
rect 8741 470 10553 538
rect 8741 414 8751 470
rect 8807 414 8875 470
rect 8931 414 8999 470
rect 9055 414 9123 470
rect 9179 414 9247 470
rect 9303 414 9371 470
rect 9427 414 9495 470
rect 9551 414 9619 470
rect 9675 414 9743 470
rect 9799 414 9867 470
rect 9923 414 9991 470
rect 10047 414 10115 470
rect 10171 414 10239 470
rect 10295 414 10363 470
rect 10419 414 10487 470
rect 10543 414 10553 470
rect 8741 346 10553 414
rect 8741 290 8751 346
rect 8807 290 8875 346
rect 8931 290 8999 346
rect 9055 290 9123 346
rect 9179 290 9247 346
rect 9303 290 9371 346
rect 9427 290 9495 346
rect 9551 290 9619 346
rect 9675 290 9743 346
rect 9799 290 9867 346
rect 9923 290 9991 346
rect 10047 290 10115 346
rect 10171 290 10239 346
rect 10295 290 10363 346
rect 10419 290 10487 346
rect 10543 290 10553 346
rect 8741 222 10553 290
rect 8741 166 8751 222
rect 8807 166 8875 222
rect 8931 166 8999 222
rect 9055 166 9123 222
rect 9179 166 9247 222
rect 9303 166 9371 222
rect 9427 166 9495 222
rect 9551 166 9619 222
rect 9675 166 9743 222
rect 9799 166 9867 222
rect 9923 166 9991 222
rect 10047 166 10115 222
rect 10171 166 10239 222
rect 10295 166 10363 222
rect 10419 166 10487 222
rect 10543 166 10553 222
rect 8741 98 10553 166
rect 8741 42 8751 98
rect 8807 42 8875 98
rect 8931 42 8999 98
rect 9055 42 9123 98
rect 9179 42 9247 98
rect 9303 42 9371 98
rect 9427 42 9495 98
rect 9551 42 9619 98
rect 9675 42 9743 98
rect 9799 42 9867 98
rect 9923 42 9991 98
rect 10047 42 10115 98
rect 10171 42 10239 98
rect 10295 42 10363 98
rect 10419 42 10487 98
rect 10543 42 10553 98
rect 8741 32 10553 42
rect 12842 2950 13910 2960
rect 12842 2894 12852 2950
rect 12908 2894 12976 2950
rect 13032 2894 13100 2950
rect 13156 2894 13224 2950
rect 13280 2894 13348 2950
rect 13404 2894 13472 2950
rect 13528 2894 13596 2950
rect 13652 2894 13720 2950
rect 13776 2894 13844 2950
rect 13900 2894 13910 2950
rect 12842 2826 13910 2894
rect 12842 2770 12852 2826
rect 12908 2770 12976 2826
rect 13032 2770 13100 2826
rect 13156 2770 13224 2826
rect 13280 2770 13348 2826
rect 13404 2770 13472 2826
rect 13528 2770 13596 2826
rect 13652 2770 13720 2826
rect 13776 2770 13844 2826
rect 13900 2770 13910 2826
rect 12842 2702 13910 2770
rect 12842 2646 12852 2702
rect 12908 2646 12976 2702
rect 13032 2646 13100 2702
rect 13156 2646 13224 2702
rect 13280 2646 13348 2702
rect 13404 2646 13472 2702
rect 13528 2646 13596 2702
rect 13652 2646 13720 2702
rect 13776 2646 13844 2702
rect 13900 2646 13910 2702
rect 12842 2578 13910 2646
rect 12842 2522 12852 2578
rect 12908 2522 12976 2578
rect 13032 2522 13100 2578
rect 13156 2522 13224 2578
rect 13280 2522 13348 2578
rect 13404 2522 13472 2578
rect 13528 2522 13596 2578
rect 13652 2522 13720 2578
rect 13776 2522 13844 2578
rect 13900 2522 13910 2578
rect 12842 2454 13910 2522
rect 12842 2398 12852 2454
rect 12908 2398 12976 2454
rect 13032 2398 13100 2454
rect 13156 2398 13224 2454
rect 13280 2398 13348 2454
rect 13404 2398 13472 2454
rect 13528 2398 13596 2454
rect 13652 2398 13720 2454
rect 13776 2398 13844 2454
rect 13900 2398 13910 2454
rect 12842 2330 13910 2398
rect 12842 2274 12852 2330
rect 12908 2274 12976 2330
rect 13032 2274 13100 2330
rect 13156 2274 13224 2330
rect 13280 2274 13348 2330
rect 13404 2274 13472 2330
rect 13528 2274 13596 2330
rect 13652 2274 13720 2330
rect 13776 2274 13844 2330
rect 13900 2274 13910 2330
rect 12842 2206 13910 2274
rect 12842 2150 12852 2206
rect 12908 2150 12976 2206
rect 13032 2150 13100 2206
rect 13156 2150 13224 2206
rect 13280 2150 13348 2206
rect 13404 2150 13472 2206
rect 13528 2150 13596 2206
rect 13652 2150 13720 2206
rect 13776 2150 13844 2206
rect 13900 2150 13910 2206
rect 12842 2082 13910 2150
rect 12842 2026 12852 2082
rect 12908 2026 12976 2082
rect 13032 2026 13100 2082
rect 13156 2026 13224 2082
rect 13280 2026 13348 2082
rect 13404 2026 13472 2082
rect 13528 2026 13596 2082
rect 13652 2026 13720 2082
rect 13776 2026 13844 2082
rect 13900 2026 13910 2082
rect 12842 1958 13910 2026
rect 12842 1902 12852 1958
rect 12908 1902 12976 1958
rect 13032 1902 13100 1958
rect 13156 1902 13224 1958
rect 13280 1902 13348 1958
rect 13404 1902 13472 1958
rect 13528 1902 13596 1958
rect 13652 1902 13720 1958
rect 13776 1902 13844 1958
rect 13900 1902 13910 1958
rect 12842 1834 13910 1902
rect 12842 1778 12852 1834
rect 12908 1778 12976 1834
rect 13032 1778 13100 1834
rect 13156 1778 13224 1834
rect 13280 1778 13348 1834
rect 13404 1778 13472 1834
rect 13528 1778 13596 1834
rect 13652 1778 13720 1834
rect 13776 1778 13844 1834
rect 13900 1778 13910 1834
rect 12842 1710 13910 1778
rect 12842 1654 12852 1710
rect 12908 1654 12976 1710
rect 13032 1654 13100 1710
rect 13156 1654 13224 1710
rect 13280 1654 13348 1710
rect 13404 1654 13472 1710
rect 13528 1654 13596 1710
rect 13652 1654 13720 1710
rect 13776 1654 13844 1710
rect 13900 1654 13910 1710
rect 12842 1586 13910 1654
rect 12842 1530 12852 1586
rect 12908 1530 12976 1586
rect 13032 1530 13100 1586
rect 13156 1530 13224 1586
rect 13280 1530 13348 1586
rect 13404 1530 13472 1586
rect 13528 1530 13596 1586
rect 13652 1530 13720 1586
rect 13776 1530 13844 1586
rect 13900 1530 13910 1586
rect 12842 1462 13910 1530
rect 12842 1406 12852 1462
rect 12908 1406 12976 1462
rect 13032 1406 13100 1462
rect 13156 1406 13224 1462
rect 13280 1406 13348 1462
rect 13404 1406 13472 1462
rect 13528 1406 13596 1462
rect 13652 1406 13720 1462
rect 13776 1406 13844 1462
rect 13900 1406 13910 1462
rect 12842 1338 13910 1406
rect 12842 1282 12852 1338
rect 12908 1282 12976 1338
rect 13032 1282 13100 1338
rect 13156 1282 13224 1338
rect 13280 1282 13348 1338
rect 13404 1282 13472 1338
rect 13528 1282 13596 1338
rect 13652 1282 13720 1338
rect 13776 1282 13844 1338
rect 13900 1282 13910 1338
rect 12842 1214 13910 1282
rect 12842 1158 12852 1214
rect 12908 1158 12976 1214
rect 13032 1158 13100 1214
rect 13156 1158 13224 1214
rect 13280 1158 13348 1214
rect 13404 1158 13472 1214
rect 13528 1158 13596 1214
rect 13652 1158 13720 1214
rect 13776 1158 13844 1214
rect 13900 1158 13910 1214
rect 12842 1090 13910 1158
rect 12842 1034 12852 1090
rect 12908 1034 12976 1090
rect 13032 1034 13100 1090
rect 13156 1034 13224 1090
rect 13280 1034 13348 1090
rect 13404 1034 13472 1090
rect 13528 1034 13596 1090
rect 13652 1034 13720 1090
rect 13776 1034 13844 1090
rect 13900 1034 13910 1090
rect 12842 966 13910 1034
rect 12842 910 12852 966
rect 12908 910 12976 966
rect 13032 910 13100 966
rect 13156 910 13224 966
rect 13280 910 13348 966
rect 13404 910 13472 966
rect 13528 910 13596 966
rect 13652 910 13720 966
rect 13776 910 13844 966
rect 13900 910 13910 966
rect 12842 842 13910 910
rect 12842 786 12852 842
rect 12908 786 12976 842
rect 13032 786 13100 842
rect 13156 786 13224 842
rect 13280 786 13348 842
rect 13404 786 13472 842
rect 13528 786 13596 842
rect 13652 786 13720 842
rect 13776 786 13844 842
rect 13900 786 13910 842
rect 12842 718 13910 786
rect 12842 662 12852 718
rect 12908 662 12976 718
rect 13032 662 13100 718
rect 13156 662 13224 718
rect 13280 662 13348 718
rect 13404 662 13472 718
rect 13528 662 13596 718
rect 13652 662 13720 718
rect 13776 662 13844 718
rect 13900 662 13910 718
rect 12842 594 13910 662
rect 12842 538 12852 594
rect 12908 538 12976 594
rect 13032 538 13100 594
rect 13156 538 13224 594
rect 13280 538 13348 594
rect 13404 538 13472 594
rect 13528 538 13596 594
rect 13652 538 13720 594
rect 13776 538 13844 594
rect 13900 538 13910 594
rect 12842 470 13910 538
rect 12842 414 12852 470
rect 12908 414 12976 470
rect 13032 414 13100 470
rect 13156 414 13224 470
rect 13280 414 13348 470
rect 13404 414 13472 470
rect 13528 414 13596 470
rect 13652 414 13720 470
rect 13776 414 13844 470
rect 13900 414 13910 470
rect 12842 346 13910 414
rect 12842 290 12852 346
rect 12908 290 12976 346
rect 13032 290 13100 346
rect 13156 290 13224 346
rect 13280 290 13348 346
rect 13404 290 13472 346
rect 13528 290 13596 346
rect 13652 290 13720 346
rect 13776 290 13844 346
rect 13900 290 13910 346
rect 12842 222 13910 290
rect 12842 166 12852 222
rect 12908 166 12976 222
rect 13032 166 13100 222
rect 13156 166 13224 222
rect 13280 166 13348 222
rect 13404 166 13472 222
rect 13528 166 13596 222
rect 13652 166 13720 222
rect 13776 166 13844 222
rect 13900 166 13910 222
rect 12842 98 13910 166
rect 12842 42 12852 98
rect 12908 42 12976 98
rect 13032 42 13100 98
rect 13156 42 13224 98
rect 13280 42 13348 98
rect 13404 42 13472 98
rect 13528 42 13596 98
rect 13652 42 13720 98
rect 13776 42 13844 98
rect 13900 42 13910 98
rect 12842 32 13910 42
<< via2 >>
rect 14767 50970 14823 50972
rect 14767 50918 14769 50970
rect 14769 50918 14821 50970
rect 14821 50918 14823 50970
rect 14767 50862 14823 50918
rect 14767 50810 14769 50862
rect 14769 50810 14821 50862
rect 14821 50810 14823 50862
rect 14767 50754 14823 50810
rect 14767 50702 14769 50754
rect 14769 50702 14821 50754
rect 14821 50702 14823 50754
rect 14767 50646 14823 50702
rect 14767 50594 14769 50646
rect 14769 50594 14821 50646
rect 14821 50594 14823 50646
rect 14767 50538 14823 50594
rect 14767 50486 14769 50538
rect 14769 50486 14821 50538
rect 14821 50486 14823 50538
rect 14767 50430 14823 50486
rect 14767 50378 14769 50430
rect 14769 50378 14821 50430
rect 14821 50378 14823 50430
rect 14767 50322 14823 50378
rect 14767 50270 14769 50322
rect 14769 50270 14821 50322
rect 14821 50270 14823 50322
rect 14767 50214 14823 50270
rect 14767 50162 14769 50214
rect 14769 50162 14821 50214
rect 14821 50162 14823 50214
rect 14767 50106 14823 50162
rect 14767 50054 14769 50106
rect 14769 50054 14821 50106
rect 14821 50054 14823 50106
rect 14767 49998 14823 50054
rect 14767 49946 14769 49998
rect 14769 49946 14821 49998
rect 14821 49946 14823 49998
rect 14767 49890 14823 49946
rect 14767 49838 14769 49890
rect 14769 49838 14821 49890
rect 14821 49838 14823 49890
rect 14767 49782 14823 49838
rect 14767 49730 14769 49782
rect 14769 49730 14821 49782
rect 14821 49730 14823 49782
rect 14767 49674 14823 49730
rect 14767 49622 14769 49674
rect 14769 49622 14821 49674
rect 14821 49622 14823 49674
rect 14767 49620 14823 49622
rect 6394 46614 6450 46670
rect 6394 46490 6450 46546
rect 6394 46366 6450 46422
rect 4470 46267 4526 46323
rect 6394 46242 6450 46298
rect 4470 46143 4526 46199
rect 4470 46019 4526 46075
rect 4470 45895 4526 45951
rect 4470 45771 4526 45827
rect 4470 45647 4526 45703
rect 4470 45523 4526 45579
rect 4470 45399 4526 45455
rect 4470 45275 4526 45331
rect 1104 45199 1160 45255
rect 4470 45151 4526 45207
rect 1104 45075 1160 45131
rect 1104 44951 1160 45007
rect 1104 44827 1160 44883
rect 1104 44703 1160 44759
rect 1104 44579 1160 44635
rect 1104 44455 1160 44511
rect 1104 44331 1160 44387
rect 1104 44207 1160 44263
rect 1104 44083 1160 44139
rect 1104 43959 1160 44015
rect 1104 43835 1160 43891
rect 1104 43711 1160 43767
rect 1104 43587 1160 43643
rect 1104 43463 1160 43519
rect 1228 45075 1284 45131
rect 4470 45027 4526 45083
rect 1228 44951 1284 45007
rect 1228 44827 1284 44883
rect 1228 44703 1284 44759
rect 1228 44579 1284 44635
rect 1228 44455 1284 44511
rect 1228 44331 1284 44387
rect 1228 44207 1284 44263
rect 1228 44083 1284 44139
rect 1228 43959 1284 44015
rect 1228 43835 1284 43891
rect 1228 43711 1284 43767
rect 1228 43587 1284 43643
rect 1228 43463 1284 43519
rect 1228 43339 1284 43395
rect 1352 44951 1408 45007
rect 4470 44903 4526 44959
rect 1352 44827 1408 44883
rect 1352 44703 1408 44759
rect 1352 44579 1408 44635
rect 1352 44455 1408 44511
rect 1352 44331 1408 44387
rect 1352 44207 1408 44263
rect 1352 44083 1408 44139
rect 1352 43959 1408 44015
rect 1352 43835 1408 43891
rect 1352 43711 1408 43767
rect 1352 43587 1408 43643
rect 1352 43463 1408 43519
rect 1352 43339 1408 43395
rect 1352 43215 1408 43271
rect 1476 44827 1532 44883
rect 4470 44779 4526 44835
rect 1476 44703 1532 44759
rect 1476 44579 1532 44635
rect 1476 44455 1532 44511
rect 1476 44331 1532 44387
rect 1476 44207 1532 44263
rect 1476 44083 1532 44139
rect 1476 43959 1532 44015
rect 1476 43835 1532 43891
rect 1476 43711 1532 43767
rect 1476 43587 1532 43643
rect 1476 43463 1532 43519
rect 1476 43339 1532 43395
rect 1476 43215 1532 43271
rect 1476 43091 1532 43147
rect 1600 44703 1656 44759
rect 4470 44655 4526 44711
rect 4594 46143 4650 46199
rect 6394 46118 6450 46174
rect 4594 46019 4650 46075
rect 4594 45895 4650 45951
rect 4594 45771 4650 45827
rect 4594 45647 4650 45703
rect 4594 45523 4650 45579
rect 4594 45399 4650 45455
rect 4594 45275 4650 45331
rect 4594 45151 4650 45207
rect 4594 45027 4650 45083
rect 4594 44903 4650 44959
rect 4594 44779 4650 44835
rect 4594 44655 4650 44711
rect 1600 44579 1656 44635
rect 1600 44455 1656 44511
rect 1600 44331 1656 44387
rect 1600 44207 1656 44263
rect 1600 44083 1656 44139
rect 1600 43959 1656 44015
rect 1600 43835 1656 43891
rect 1600 43711 1656 43767
rect 1600 43587 1656 43643
rect 1600 43463 1656 43519
rect 1600 43339 1656 43395
rect 1600 43215 1656 43271
rect 1600 43091 1656 43147
rect 1600 42967 1656 43023
rect 1724 44579 1780 44635
rect 4594 44531 4650 44587
rect 4718 46019 4774 46075
rect 6394 45994 6450 46050
rect 4718 45895 4774 45951
rect 4718 45771 4774 45827
rect 4718 45647 4774 45703
rect 4718 45523 4774 45579
rect 4718 45399 4774 45455
rect 4718 45275 4774 45331
rect 4718 45151 4774 45207
rect 4718 45027 4774 45083
rect 4718 44903 4774 44959
rect 4718 44779 4774 44835
rect 4718 44655 4774 44711
rect 4718 44531 4774 44587
rect 1724 44455 1780 44511
rect 1724 44331 1780 44387
rect 1724 44207 1780 44263
rect 1724 44083 1780 44139
rect 1724 43959 1780 44015
rect 1724 43835 1780 43891
rect 1724 43711 1780 43767
rect 1724 43587 1780 43643
rect 1724 43463 1780 43519
rect 1724 43339 1780 43395
rect 1724 43215 1780 43271
rect 1724 43091 1780 43147
rect 1724 42967 1780 43023
rect 1724 42843 1780 42899
rect 1848 44455 1904 44511
rect 4718 44407 4774 44463
rect 4842 45895 4898 45951
rect 6394 45870 6450 45926
rect 4842 45771 4898 45827
rect 4842 45647 4898 45703
rect 4842 45523 4898 45579
rect 4842 45399 4898 45455
rect 4842 45275 4898 45331
rect 4842 45151 4898 45207
rect 4842 45027 4898 45083
rect 4842 44903 4898 44959
rect 4842 44779 4898 44835
rect 4842 44655 4898 44711
rect 4842 44531 4898 44587
rect 4842 44407 4898 44463
rect 1848 44331 1904 44387
rect 1848 44207 1904 44263
rect 1848 44083 1904 44139
rect 1848 43959 1904 44015
rect 1848 43835 1904 43891
rect 1848 43711 1904 43767
rect 1848 43587 1904 43643
rect 1848 43463 1904 43519
rect 1848 43339 1904 43395
rect 1848 43215 1904 43271
rect 1848 43091 1904 43147
rect 1848 42967 1904 43023
rect 1848 42843 1904 42899
rect 1848 42719 1904 42775
rect 1972 44331 2028 44387
rect 4842 44283 4898 44339
rect 4966 45771 5022 45827
rect 6394 45746 6450 45802
rect 4966 45647 5022 45703
rect 4966 45523 5022 45579
rect 4966 45399 5022 45455
rect 4966 45275 5022 45331
rect 4966 45151 5022 45207
rect 4966 45027 5022 45083
rect 4966 44903 5022 44959
rect 4966 44779 5022 44835
rect 4966 44655 5022 44711
rect 4966 44531 5022 44587
rect 4966 44407 5022 44463
rect 4966 44283 5022 44339
rect 1972 44207 2028 44263
rect 4966 44159 5022 44215
rect 5090 45647 5146 45703
rect 6394 45622 6450 45678
rect 5090 45523 5146 45579
rect 5090 45399 5146 45455
rect 5090 45275 5146 45331
rect 5090 45151 5146 45207
rect 5090 45027 5146 45083
rect 5090 44903 5146 44959
rect 5090 44779 5146 44835
rect 5090 44655 5146 44711
rect 5090 44531 5146 44587
rect 5090 44407 5146 44463
rect 5090 44283 5146 44339
rect 5090 44159 5146 44215
rect 1972 44083 2028 44139
rect 5090 44035 5146 44091
rect 1972 43959 2028 44015
rect 1972 43835 2028 43891
rect 1972 43711 2028 43767
rect 1972 43587 2028 43643
rect 1972 43463 2028 43519
rect 1972 43339 2028 43395
rect 1972 43215 2028 43271
rect 1972 43091 2028 43147
rect 1972 42967 2028 43023
rect 1972 42843 2028 42899
rect 1972 42719 2028 42775
rect 1972 42595 2028 42651
rect 5214 45523 5270 45579
rect 6394 45498 6450 45554
rect 5214 45399 5270 45455
rect 5214 45275 5270 45331
rect 5214 45151 5270 45207
rect 5214 45027 5270 45083
rect 5214 44903 5270 44959
rect 5214 44779 5270 44835
rect 5214 44655 5270 44711
rect 5214 44531 5270 44587
rect 5214 44407 5270 44463
rect 5214 44283 5270 44339
rect 5214 44159 5270 44215
rect 5214 44035 5270 44091
rect 4470 43968 4526 44024
rect 5214 43911 5270 43967
rect 4470 43844 4526 43900
rect 4470 43720 4526 43776
rect 4470 43596 4526 43652
rect 4470 43472 4526 43528
rect 4470 43348 4526 43404
rect 4470 43224 4526 43280
rect 4470 43100 4526 43156
rect 4470 42976 4526 43032
rect 4470 42852 4526 42908
rect 4470 42728 4526 42784
rect 4470 42604 4526 42660
rect 4470 42480 4526 42536
rect 4470 42356 4526 42412
rect 5338 45399 5394 45455
rect 6394 45374 6450 45430
rect 5338 45275 5394 45331
rect 5338 45151 5394 45207
rect 5338 45027 5394 45083
rect 5338 44903 5394 44959
rect 5338 44779 5394 44835
rect 5338 44655 5394 44711
rect 5338 44531 5394 44587
rect 5338 44407 5394 44463
rect 5338 44283 5394 44339
rect 5338 44159 5394 44215
rect 5338 44035 5394 44091
rect 5338 43911 5394 43967
rect 4594 43844 4650 43900
rect 5338 43787 5394 43843
rect 4594 43720 4650 43776
rect 4594 43596 4650 43652
rect 4594 43472 4650 43528
rect 4594 43348 4650 43404
rect 4594 43224 4650 43280
rect 4594 43100 4650 43156
rect 4594 42976 4650 43032
rect 4594 42852 4650 42908
rect 4594 42728 4650 42784
rect 4594 42604 4650 42660
rect 4594 42480 4650 42536
rect 4594 42356 4650 42412
rect 4594 42232 4650 42288
rect 5462 45275 5518 45331
rect 6394 45250 6450 45306
rect 5462 45151 5518 45207
rect 5462 45027 5518 45083
rect 5462 44903 5518 44959
rect 5462 44779 5518 44835
rect 5462 44655 5518 44711
rect 5462 44531 5518 44587
rect 5462 44407 5518 44463
rect 5462 44283 5518 44339
rect 5462 44159 5518 44215
rect 5462 44035 5518 44091
rect 5462 43911 5518 43967
rect 5462 43787 5518 43843
rect 4718 43720 4774 43776
rect 5462 43663 5518 43719
rect 4718 43596 4774 43652
rect 4718 43472 4774 43528
rect 4718 43348 4774 43404
rect 4718 43224 4774 43280
rect 4718 43100 4774 43156
rect 4718 42976 4774 43032
rect 4718 42852 4774 42908
rect 4718 42728 4774 42784
rect 4718 42604 4774 42660
rect 4718 42480 4774 42536
rect 4718 42356 4774 42412
rect 4718 42232 4774 42288
rect 4718 42108 4774 42164
rect 5586 45151 5642 45207
rect 6394 45126 6450 45182
rect 5586 45027 5642 45083
rect 5586 44903 5642 44959
rect 5586 44779 5642 44835
rect 5586 44655 5642 44711
rect 5586 44531 5642 44587
rect 5586 44407 5642 44463
rect 5586 44283 5642 44339
rect 5586 44159 5642 44215
rect 5586 44035 5642 44091
rect 5586 43911 5642 43967
rect 5586 43787 5642 43843
rect 5586 43663 5642 43719
rect 4842 43596 4898 43652
rect 5586 43539 5642 43595
rect 4842 43472 4898 43528
rect 4842 43348 4898 43404
rect 4842 43224 4898 43280
rect 4842 43100 4898 43156
rect 4842 42976 4898 43032
rect 4842 42852 4898 42908
rect 4842 42728 4898 42784
rect 4842 42604 4898 42660
rect 4842 42480 4898 42536
rect 4842 42356 4898 42412
rect 4842 42232 4898 42288
rect 4842 42108 4898 42164
rect 4842 41984 4898 42040
rect 5710 45027 5766 45083
rect 6394 45002 6450 45058
rect 6518 46490 6574 46546
rect 6518 46366 6574 46422
rect 6518 46242 6574 46298
rect 6518 46118 6574 46174
rect 6518 45994 6574 46050
rect 6518 45870 6574 45926
rect 6518 45746 6574 45802
rect 6518 45622 6574 45678
rect 6518 45498 6574 45554
rect 6518 45374 6574 45430
rect 6518 45250 6574 45306
rect 6518 45126 6574 45182
rect 6518 45002 6574 45058
rect 5710 44903 5766 44959
rect 5710 44779 5766 44835
rect 5710 44655 5766 44711
rect 5710 44531 5766 44587
rect 5710 44407 5766 44463
rect 5710 44283 5766 44339
rect 5710 44159 5766 44215
rect 5710 44035 5766 44091
rect 5710 43911 5766 43967
rect 5710 43787 5766 43843
rect 5710 43663 5766 43719
rect 5710 43539 5766 43595
rect 4966 43472 5022 43528
rect 5710 43415 5766 43471
rect 4966 43348 5022 43404
rect 4966 43224 5022 43280
rect 4966 43100 5022 43156
rect 4966 42976 5022 43032
rect 4966 42852 5022 42908
rect 4966 42728 5022 42784
rect 4966 42604 5022 42660
rect 4966 42480 5022 42536
rect 4966 42356 5022 42412
rect 4966 42232 5022 42288
rect 4966 42108 5022 42164
rect 4966 41984 5022 42040
rect 4966 41860 5022 41916
rect 5834 44903 5890 44959
rect 6518 44878 6574 44934
rect 6642 46366 6698 46422
rect 6642 46242 6698 46298
rect 6642 46118 6698 46174
rect 6642 45994 6698 46050
rect 6642 45870 6698 45926
rect 6642 45746 6698 45802
rect 6642 45622 6698 45678
rect 6642 45498 6698 45554
rect 6642 45374 6698 45430
rect 6642 45250 6698 45306
rect 6642 45126 6698 45182
rect 6642 45002 6698 45058
rect 6642 44878 6698 44934
rect 5834 44779 5890 44835
rect 5834 44655 5890 44711
rect 5834 44531 5890 44587
rect 5834 44407 5890 44463
rect 5834 44283 5890 44339
rect 5834 44159 5890 44215
rect 5834 44035 5890 44091
rect 5834 43911 5890 43967
rect 5834 43787 5890 43843
rect 5834 43663 5890 43719
rect 5834 43539 5890 43595
rect 5834 43415 5890 43471
rect 5090 43348 5146 43404
rect 5834 43291 5890 43347
rect 5090 43224 5146 43280
rect 5090 43100 5146 43156
rect 5090 42976 5146 43032
rect 5090 42852 5146 42908
rect 5090 42728 5146 42784
rect 5090 42604 5146 42660
rect 5090 42480 5146 42536
rect 5090 42356 5146 42412
rect 5090 42232 5146 42288
rect 5090 42108 5146 42164
rect 5090 41984 5146 42040
rect 5090 41860 5146 41916
rect 4470 41733 4526 41789
rect 5090 41736 5146 41792
rect 5958 44779 6014 44835
rect 6642 44754 6698 44810
rect 6766 46242 6822 46298
rect 6766 46118 6822 46174
rect 6766 45994 6822 46050
rect 6766 45870 6822 45926
rect 6766 45746 6822 45802
rect 6766 45622 6822 45678
rect 6766 45498 6822 45554
rect 6766 45374 6822 45430
rect 6766 45250 6822 45306
rect 6766 45126 6822 45182
rect 6766 45002 6822 45058
rect 6766 44878 6822 44934
rect 6766 44754 6822 44810
rect 5958 44655 6014 44711
rect 5958 44531 6014 44587
rect 5958 44407 6014 44463
rect 5958 44283 6014 44339
rect 5958 44159 6014 44215
rect 5958 44035 6014 44091
rect 5958 43911 6014 43967
rect 5958 43787 6014 43843
rect 5958 43663 6014 43719
rect 5958 43539 6014 43595
rect 5958 43415 6014 43471
rect 5958 43291 6014 43347
rect 5214 43224 5270 43280
rect 5958 43167 6014 43223
rect 5214 43100 5270 43156
rect 5214 42976 5270 43032
rect 5214 42852 5270 42908
rect 5214 42728 5270 42784
rect 5214 42604 5270 42660
rect 5214 42480 5270 42536
rect 5214 42356 5270 42412
rect 5214 42232 5270 42288
rect 5214 42108 5270 42164
rect 5214 41984 5270 42040
rect 5214 41860 5270 41916
rect 5214 41736 5270 41792
rect 4470 41609 4526 41665
rect 4470 41485 4526 41541
rect 4470 41361 4526 41417
rect 4470 41237 4526 41293
rect 4470 41113 4526 41169
rect 4470 40989 4526 41045
rect 4470 40865 4526 40921
rect 4470 40741 4526 40797
rect 4470 40617 4526 40673
rect 4470 40493 4526 40549
rect 4470 40369 4526 40425
rect 4470 40245 4526 40301
rect 4470 40121 4526 40177
rect 4594 41609 4650 41665
rect 5214 41612 5270 41668
rect 6082 44655 6138 44711
rect 6766 44630 6822 44686
rect 6890 46118 6946 46174
rect 6890 45994 6946 46050
rect 6890 45870 6946 45926
rect 6890 45746 6946 45802
rect 6890 45622 6946 45678
rect 6890 45498 6946 45554
rect 6890 45374 6946 45430
rect 6890 45250 6946 45306
rect 6890 45126 6946 45182
rect 6890 45002 6946 45058
rect 6890 44878 6946 44934
rect 6890 44754 6946 44810
rect 6890 44630 6946 44686
rect 6082 44531 6138 44587
rect 6890 44506 6946 44562
rect 7014 45994 7070 46050
rect 7014 45870 7070 45926
rect 7014 45746 7070 45802
rect 7014 45622 7070 45678
rect 7014 45498 7070 45554
rect 7014 45374 7070 45430
rect 7014 45250 7070 45306
rect 7014 45126 7070 45182
rect 7014 45002 7070 45058
rect 7014 44878 7070 44934
rect 7014 44754 7070 44810
rect 7014 44630 7070 44686
rect 7014 44506 7070 44562
rect 6082 44407 6138 44463
rect 7014 44382 7070 44438
rect 7138 45870 7194 45926
rect 7138 45746 7194 45802
rect 7138 45622 7194 45678
rect 7138 45498 7194 45554
rect 7138 45374 7194 45430
rect 7138 45250 7194 45306
rect 7138 45126 7194 45182
rect 7138 45002 7194 45058
rect 7138 44878 7194 44934
rect 7138 44754 7194 44810
rect 7138 44630 7194 44686
rect 7138 44506 7194 44562
rect 7138 44382 7194 44438
rect 6082 44283 6138 44339
rect 7138 44258 7194 44314
rect 7262 45746 7318 45802
rect 7262 45622 7318 45678
rect 7262 45498 7318 45554
rect 7262 45374 7318 45430
rect 7262 45250 7318 45306
rect 7262 45126 7318 45182
rect 7262 45002 7318 45058
rect 7262 44878 7318 44934
rect 7262 44754 7318 44810
rect 7262 44630 7318 44686
rect 7262 44506 7318 44562
rect 7262 44382 7318 44438
rect 7262 44258 7318 44314
rect 6082 44159 6138 44215
rect 7262 44134 7318 44190
rect 8751 44488 8807 44544
rect 8875 44488 8931 44544
rect 8999 44488 9055 44544
rect 9123 44488 9179 44544
rect 9247 44488 9303 44544
rect 9371 44488 9427 44544
rect 9495 44488 9551 44544
rect 9619 44488 9675 44544
rect 9743 44488 9799 44544
rect 9867 44488 9923 44544
rect 9991 44488 10047 44544
rect 10115 44488 10171 44544
rect 10239 44488 10295 44544
rect 10363 44488 10419 44544
rect 10487 44488 10543 44544
rect 8751 44364 8807 44420
rect 8875 44364 8931 44420
rect 8999 44364 9055 44420
rect 9123 44364 9179 44420
rect 9247 44364 9303 44420
rect 9371 44364 9427 44420
rect 9495 44364 9551 44420
rect 9619 44364 9675 44420
rect 9743 44364 9799 44420
rect 9867 44364 9923 44420
rect 9991 44364 10047 44420
rect 10115 44364 10171 44420
rect 10239 44364 10295 44420
rect 10363 44364 10419 44420
rect 10487 44364 10543 44420
rect 8751 44240 8807 44296
rect 8875 44240 8931 44296
rect 8999 44240 9055 44296
rect 9123 44240 9179 44296
rect 9247 44240 9303 44296
rect 9371 44240 9427 44296
rect 9495 44240 9551 44296
rect 9619 44240 9675 44296
rect 9743 44240 9799 44296
rect 9867 44240 9923 44296
rect 9991 44240 10047 44296
rect 10115 44240 10171 44296
rect 10239 44240 10295 44296
rect 10363 44240 10419 44296
rect 10487 44240 10543 44296
rect 6082 44035 6138 44091
rect 6082 43911 6138 43967
rect 6082 43787 6138 43843
rect 6082 43663 6138 43719
rect 6082 43539 6138 43595
rect 6082 43415 6138 43471
rect 6082 43291 6138 43347
rect 8751 44116 8807 44172
rect 8875 44116 8931 44172
rect 8999 44116 9055 44172
rect 9123 44116 9179 44172
rect 9247 44116 9303 44172
rect 9371 44116 9427 44172
rect 9495 44116 9551 44172
rect 9619 44116 9675 44172
rect 9743 44116 9799 44172
rect 9867 44116 9923 44172
rect 9991 44116 10047 44172
rect 10115 44116 10171 44172
rect 10239 44116 10295 44172
rect 10363 44116 10419 44172
rect 10487 44116 10543 44172
rect 8751 43992 8807 44048
rect 8875 43992 8931 44048
rect 8999 43992 9055 44048
rect 9123 43992 9179 44048
rect 9247 43992 9303 44048
rect 9371 43992 9427 44048
rect 9495 43992 9551 44048
rect 9619 43992 9675 44048
rect 9743 43992 9799 44048
rect 9867 43992 9923 44048
rect 9991 43992 10047 44048
rect 10115 43992 10171 44048
rect 10239 43992 10295 44048
rect 10363 43992 10419 44048
rect 10487 43992 10543 44048
rect 8751 43868 8807 43924
rect 8875 43868 8931 43924
rect 8999 43868 9055 43924
rect 9123 43868 9179 43924
rect 9247 43868 9303 43924
rect 9371 43868 9427 43924
rect 9495 43868 9551 43924
rect 9619 43868 9675 43924
rect 9743 43868 9799 43924
rect 9867 43868 9923 43924
rect 9991 43868 10047 43924
rect 10115 43868 10171 43924
rect 10239 43868 10295 43924
rect 10363 43868 10419 43924
rect 10487 43868 10543 43924
rect 8751 43744 8807 43800
rect 8875 43744 8931 43800
rect 8999 43744 9055 43800
rect 9123 43744 9179 43800
rect 9247 43744 9303 43800
rect 9371 43744 9427 43800
rect 9495 43744 9551 43800
rect 9619 43744 9675 43800
rect 9743 43744 9799 43800
rect 9867 43744 9923 43800
rect 9991 43744 10047 43800
rect 10115 43744 10171 43800
rect 10239 43744 10295 43800
rect 10363 43744 10419 43800
rect 10487 43744 10543 43800
rect 8751 43620 8807 43676
rect 8875 43620 8931 43676
rect 8999 43620 9055 43676
rect 9123 43620 9179 43676
rect 9247 43620 9303 43676
rect 9371 43620 9427 43676
rect 9495 43620 9551 43676
rect 9619 43620 9675 43676
rect 9743 43620 9799 43676
rect 9867 43620 9923 43676
rect 9991 43620 10047 43676
rect 10115 43620 10171 43676
rect 10239 43620 10295 43676
rect 10363 43620 10419 43676
rect 10487 43620 10543 43676
rect 8751 43496 8807 43552
rect 8875 43496 8931 43552
rect 8999 43496 9055 43552
rect 9123 43496 9179 43552
rect 9247 43496 9303 43552
rect 9371 43496 9427 43552
rect 9495 43496 9551 43552
rect 9619 43496 9675 43552
rect 9743 43496 9799 43552
rect 9867 43496 9923 43552
rect 9991 43496 10047 43552
rect 10115 43496 10171 43552
rect 10239 43496 10295 43552
rect 10363 43496 10419 43552
rect 10487 43496 10543 43552
rect 8751 43372 8807 43428
rect 8875 43372 8931 43428
rect 8999 43372 9055 43428
rect 9123 43372 9179 43428
rect 9247 43372 9303 43428
rect 9371 43372 9427 43428
rect 9495 43372 9551 43428
rect 9619 43372 9675 43428
rect 9743 43372 9799 43428
rect 9867 43372 9923 43428
rect 9991 43372 10047 43428
rect 10115 43372 10171 43428
rect 10239 43372 10295 43428
rect 10363 43372 10419 43428
rect 10487 43372 10543 43428
rect 8751 43248 8807 43304
rect 8875 43248 8931 43304
rect 8999 43248 9055 43304
rect 9123 43248 9179 43304
rect 9247 43248 9303 43304
rect 9371 43248 9427 43304
rect 9495 43248 9551 43304
rect 9619 43248 9675 43304
rect 9743 43248 9799 43304
rect 9867 43248 9923 43304
rect 9991 43248 10047 43304
rect 10115 43248 10171 43304
rect 10239 43248 10295 43304
rect 10363 43248 10419 43304
rect 10487 43248 10543 43304
rect 12852 44488 12908 44544
rect 12976 44488 13032 44544
rect 13100 44488 13156 44544
rect 13224 44488 13280 44544
rect 13348 44488 13404 44544
rect 13472 44488 13528 44544
rect 13596 44488 13652 44544
rect 13720 44488 13776 44544
rect 13844 44488 13900 44544
rect 12852 44364 12908 44420
rect 12976 44364 13032 44420
rect 13100 44364 13156 44420
rect 13224 44364 13280 44420
rect 13348 44364 13404 44420
rect 13472 44364 13528 44420
rect 13596 44364 13652 44420
rect 13720 44364 13776 44420
rect 13844 44364 13900 44420
rect 12852 44240 12908 44296
rect 12976 44240 13032 44296
rect 13100 44240 13156 44296
rect 13224 44240 13280 44296
rect 13348 44240 13404 44296
rect 13472 44240 13528 44296
rect 13596 44240 13652 44296
rect 13720 44240 13776 44296
rect 13844 44240 13900 44296
rect 12852 44116 12908 44172
rect 12976 44116 13032 44172
rect 13100 44116 13156 44172
rect 13224 44116 13280 44172
rect 13348 44116 13404 44172
rect 13472 44116 13528 44172
rect 13596 44116 13652 44172
rect 13720 44116 13776 44172
rect 13844 44116 13900 44172
rect 12852 43992 12908 44048
rect 12976 43992 13032 44048
rect 13100 43992 13156 44048
rect 13224 43992 13280 44048
rect 13348 43992 13404 44048
rect 13472 43992 13528 44048
rect 13596 43992 13652 44048
rect 13720 43992 13776 44048
rect 13844 43992 13900 44048
rect 12852 43868 12908 43924
rect 12976 43868 13032 43924
rect 13100 43868 13156 43924
rect 13224 43868 13280 43924
rect 13348 43868 13404 43924
rect 13472 43868 13528 43924
rect 13596 43868 13652 43924
rect 13720 43868 13776 43924
rect 13844 43868 13900 43924
rect 12852 43744 12908 43800
rect 12976 43744 13032 43800
rect 13100 43744 13156 43800
rect 13224 43744 13280 43800
rect 13348 43744 13404 43800
rect 13472 43744 13528 43800
rect 13596 43744 13652 43800
rect 13720 43744 13776 43800
rect 13844 43744 13900 43800
rect 12852 43620 12908 43676
rect 12976 43620 13032 43676
rect 13100 43620 13156 43676
rect 13224 43620 13280 43676
rect 13348 43620 13404 43676
rect 13472 43620 13528 43676
rect 13596 43620 13652 43676
rect 13720 43620 13776 43676
rect 13844 43620 13900 43676
rect 12852 43496 12908 43552
rect 12976 43496 13032 43552
rect 13100 43496 13156 43552
rect 13224 43496 13280 43552
rect 13348 43496 13404 43552
rect 13472 43496 13528 43552
rect 13596 43496 13652 43552
rect 13720 43496 13776 43552
rect 13844 43496 13900 43552
rect 12852 43372 12908 43428
rect 12976 43372 13032 43428
rect 13100 43372 13156 43428
rect 13224 43372 13280 43428
rect 13348 43372 13404 43428
rect 13472 43372 13528 43428
rect 13596 43372 13652 43428
rect 13720 43372 13776 43428
rect 13844 43372 13900 43428
rect 12852 43248 12908 43304
rect 12976 43248 13032 43304
rect 13100 43248 13156 43304
rect 13224 43248 13280 43304
rect 13348 43248 13404 43304
rect 13472 43248 13528 43304
rect 13596 43248 13652 43304
rect 13720 43248 13776 43304
rect 13844 43248 13900 43304
rect 6082 43167 6138 43223
rect 5338 43100 5394 43156
rect 6082 43043 6138 43099
rect 5338 42976 5394 43032
rect 5338 42852 5394 42908
rect 5338 42728 5394 42784
rect 5338 42604 5394 42660
rect 5338 42480 5394 42536
rect 5338 42356 5394 42412
rect 5338 42232 5394 42288
rect 5338 42108 5394 42164
rect 5338 41984 5394 42040
rect 5338 41860 5394 41916
rect 5338 41736 5394 41792
rect 5338 41612 5394 41668
rect 4594 41485 4650 41541
rect 4594 41361 4650 41417
rect 4594 41237 4650 41293
rect 4594 41113 4650 41169
rect 4594 40989 4650 41045
rect 4594 40865 4650 40921
rect 4594 40741 4650 40797
rect 4594 40617 4650 40673
rect 4594 40493 4650 40549
rect 4594 40369 4650 40425
rect 4594 40245 4650 40301
rect 4594 40121 4650 40177
rect 4594 39997 4650 40053
rect 4718 41485 4774 41541
rect 5338 41488 5394 41544
rect 5462 42976 5518 43032
rect 5462 42852 5518 42908
rect 5462 42728 5518 42784
rect 5462 42604 5518 42660
rect 5462 42480 5518 42536
rect 5462 42356 5518 42412
rect 5462 42232 5518 42288
rect 5462 42108 5518 42164
rect 5462 41984 5518 42040
rect 5462 41860 5518 41916
rect 5462 41736 5518 41792
rect 5462 41612 5518 41668
rect 5462 41488 5518 41544
rect 4718 41361 4774 41417
rect 4718 41237 4774 41293
rect 4718 41113 4774 41169
rect 4718 40989 4774 41045
rect 4718 40865 4774 40921
rect 4718 40741 4774 40797
rect 4718 40617 4774 40673
rect 4718 40493 4774 40549
rect 4718 40369 4774 40425
rect 4718 40245 4774 40301
rect 4718 40121 4774 40177
rect 4718 39997 4774 40053
rect 4718 39873 4774 39929
rect 4842 41361 4898 41417
rect 5462 41364 5518 41420
rect 5586 42852 5642 42908
rect 7562 42888 7618 42944
rect 7686 42888 7742 42944
rect 7810 42888 7866 42944
rect 7934 42888 7990 42944
rect 8058 42888 8114 42944
rect 8182 42888 8238 42944
rect 8306 42888 8362 42944
rect 8430 42888 8486 42944
rect 8554 42888 8610 42944
rect 5586 42728 5642 42784
rect 5586 42604 5642 42660
rect 5586 42480 5642 42536
rect 5586 42356 5642 42412
rect 5586 42232 5642 42288
rect 5586 42108 5642 42164
rect 5586 41984 5642 42040
rect 5586 41860 5642 41916
rect 5586 41736 5642 41792
rect 5586 41612 5642 41668
rect 5586 41488 5642 41544
rect 5586 41364 5642 41420
rect 4842 41237 4898 41293
rect 4842 41113 4898 41169
rect 4842 40989 4898 41045
rect 4842 40865 4898 40921
rect 4842 40741 4898 40797
rect 4842 40617 4898 40673
rect 4842 40493 4898 40549
rect 4842 40369 4898 40425
rect 4842 40245 4898 40301
rect 4842 40121 4898 40177
rect 4842 39997 4898 40053
rect 4842 39873 4898 39929
rect 4842 39749 4898 39805
rect 4966 41237 5022 41293
rect 5586 41240 5642 41296
rect 5710 42728 5766 42784
rect 7562 42764 7618 42820
rect 7686 42764 7742 42820
rect 7810 42764 7866 42820
rect 7934 42764 7990 42820
rect 8058 42764 8114 42820
rect 8182 42764 8238 42820
rect 8306 42764 8362 42820
rect 8430 42764 8486 42820
rect 8554 42764 8610 42820
rect 5710 42604 5766 42660
rect 5710 42480 5766 42536
rect 5710 42356 5766 42412
rect 5710 42232 5766 42288
rect 5710 42108 5766 42164
rect 5710 41984 5766 42040
rect 5710 41860 5766 41916
rect 5710 41736 5766 41792
rect 5710 41612 5766 41668
rect 5710 41488 5766 41544
rect 5710 41364 5766 41420
rect 5710 41240 5766 41296
rect 4966 41113 5022 41169
rect 4966 40989 5022 41045
rect 4966 40865 5022 40921
rect 4966 40741 5022 40797
rect 4966 40617 5022 40673
rect 4966 40493 5022 40549
rect 4966 40369 5022 40425
rect 4966 40245 5022 40301
rect 4966 40121 5022 40177
rect 4966 39997 5022 40053
rect 4966 39873 5022 39929
rect 4966 39749 5022 39805
rect 4966 39625 5022 39681
rect 5090 41113 5146 41169
rect 5710 41116 5766 41172
rect 5834 42604 5890 42660
rect 7562 42640 7618 42696
rect 7686 42640 7742 42696
rect 7810 42640 7866 42696
rect 7934 42640 7990 42696
rect 8058 42640 8114 42696
rect 8182 42640 8238 42696
rect 8306 42640 8362 42696
rect 8430 42640 8486 42696
rect 8554 42640 8610 42696
rect 5834 42480 5890 42536
rect 5834 42356 5890 42412
rect 5834 42232 5890 42288
rect 5834 42108 5890 42164
rect 5834 41984 5890 42040
rect 5834 41860 5890 41916
rect 5834 41736 5890 41792
rect 5834 41612 5890 41668
rect 5834 41488 5890 41544
rect 5834 41364 5890 41420
rect 5834 41240 5890 41296
rect 5834 41116 5890 41172
rect 5090 40989 5146 41045
rect 5090 40865 5146 40921
rect 5090 40741 5146 40797
rect 5090 40617 5146 40673
rect 5090 40493 5146 40549
rect 5090 40369 5146 40425
rect 5090 40245 5146 40301
rect 5090 40121 5146 40177
rect 5090 39997 5146 40053
rect 5090 39873 5146 39929
rect 5090 39749 5146 39805
rect 5090 39625 5146 39681
rect 5090 39501 5146 39557
rect 5214 40989 5270 41045
rect 5834 40992 5890 41048
rect 5958 42480 6014 42536
rect 7562 42516 7618 42572
rect 7686 42516 7742 42572
rect 7810 42516 7866 42572
rect 7934 42516 7990 42572
rect 8058 42516 8114 42572
rect 8182 42516 8238 42572
rect 8306 42516 8362 42572
rect 8430 42516 8486 42572
rect 8554 42516 8610 42572
rect 5958 42356 6014 42412
rect 5958 42232 6014 42288
rect 5958 42108 6014 42164
rect 5958 41984 6014 42040
rect 5958 41860 6014 41916
rect 5958 41736 6014 41792
rect 5958 41612 6014 41668
rect 5958 41488 6014 41544
rect 5958 41364 6014 41420
rect 5958 41240 6014 41296
rect 5958 41116 6014 41172
rect 5958 40992 6014 41048
rect 5214 40865 5270 40921
rect 5214 40741 5270 40797
rect 5214 40617 5270 40673
rect 5214 40493 5270 40549
rect 5214 40369 5270 40425
rect 5214 40245 5270 40301
rect 5214 40121 5270 40177
rect 5214 39997 5270 40053
rect 5214 39873 5270 39929
rect 5214 39749 5270 39805
rect 5214 39625 5270 39681
rect 5214 39501 5270 39557
rect 5214 39377 5270 39433
rect 5338 40865 5394 40921
rect 5958 40868 6014 40924
rect 6082 42356 6138 42412
rect 6082 42232 6138 42288
rect 6082 42108 6138 42164
rect 6082 41984 6138 42040
rect 6082 41860 6138 41916
rect 6082 41736 6138 41792
rect 6082 41612 6138 41668
rect 7562 42392 7618 42448
rect 7686 42392 7742 42448
rect 7810 42392 7866 42448
rect 7934 42392 7990 42448
rect 8058 42392 8114 42448
rect 8182 42392 8238 42448
rect 8306 42392 8362 42448
rect 8430 42392 8486 42448
rect 8554 42392 8610 42448
rect 7562 42268 7618 42324
rect 7686 42268 7742 42324
rect 7810 42268 7866 42324
rect 7934 42268 7990 42324
rect 8058 42268 8114 42324
rect 8182 42268 8238 42324
rect 8306 42268 8362 42324
rect 8430 42268 8486 42324
rect 8554 42268 8610 42324
rect 7562 42144 7618 42200
rect 7686 42144 7742 42200
rect 7810 42144 7866 42200
rect 7934 42144 7990 42200
rect 8058 42144 8114 42200
rect 8182 42144 8238 42200
rect 8306 42144 8362 42200
rect 8430 42144 8486 42200
rect 8554 42144 8610 42200
rect 7562 42020 7618 42076
rect 7686 42020 7742 42076
rect 7810 42020 7866 42076
rect 7934 42020 7990 42076
rect 8058 42020 8114 42076
rect 8182 42020 8238 42076
rect 8306 42020 8362 42076
rect 8430 42020 8486 42076
rect 8554 42020 8610 42076
rect 7562 41896 7618 41952
rect 7686 41896 7742 41952
rect 7810 41896 7866 41952
rect 7934 41896 7990 41952
rect 8058 41896 8114 41952
rect 8182 41896 8238 41952
rect 8306 41896 8362 41952
rect 8430 41896 8486 41952
rect 8554 41896 8610 41952
rect 7562 41772 7618 41828
rect 7686 41772 7742 41828
rect 7810 41772 7866 41828
rect 7934 41772 7990 41828
rect 8058 41772 8114 41828
rect 8182 41772 8238 41828
rect 8306 41772 8362 41828
rect 8430 41772 8486 41828
rect 8554 41772 8610 41828
rect 7562 41648 7618 41704
rect 7686 41648 7742 41704
rect 7810 41648 7866 41704
rect 7934 41648 7990 41704
rect 8058 41648 8114 41704
rect 8182 41648 8238 41704
rect 8306 41648 8362 41704
rect 8430 41648 8486 41704
rect 8554 41648 8610 41704
rect 10679 42888 10735 42944
rect 10803 42888 10859 42944
rect 10927 42888 10983 42944
rect 11051 42888 11107 42944
rect 11175 42888 11231 42944
rect 11299 42888 11355 42944
rect 11423 42888 11479 42944
rect 11547 42888 11603 42944
rect 11671 42888 11727 42944
rect 11795 42888 11851 42944
rect 11919 42888 11975 42944
rect 12043 42888 12099 42944
rect 12167 42888 12223 42944
rect 12291 42888 12347 42944
rect 12415 42888 12471 42944
rect 10679 42764 10735 42820
rect 10803 42764 10859 42820
rect 10927 42764 10983 42820
rect 11051 42764 11107 42820
rect 11175 42764 11231 42820
rect 11299 42764 11355 42820
rect 11423 42764 11479 42820
rect 11547 42764 11603 42820
rect 11671 42764 11727 42820
rect 11795 42764 11851 42820
rect 11919 42764 11975 42820
rect 12043 42764 12099 42820
rect 12167 42764 12223 42820
rect 12291 42764 12347 42820
rect 12415 42764 12471 42820
rect 10679 42640 10735 42696
rect 10803 42640 10859 42696
rect 10927 42640 10983 42696
rect 11051 42640 11107 42696
rect 11175 42640 11231 42696
rect 11299 42640 11355 42696
rect 11423 42640 11479 42696
rect 11547 42640 11603 42696
rect 11671 42640 11727 42696
rect 11795 42640 11851 42696
rect 11919 42640 11975 42696
rect 12043 42640 12099 42696
rect 12167 42640 12223 42696
rect 12291 42640 12347 42696
rect 12415 42640 12471 42696
rect 10679 42516 10735 42572
rect 10803 42516 10859 42572
rect 10927 42516 10983 42572
rect 11051 42516 11107 42572
rect 11175 42516 11231 42572
rect 11299 42516 11355 42572
rect 11423 42516 11479 42572
rect 11547 42516 11603 42572
rect 11671 42516 11727 42572
rect 11795 42516 11851 42572
rect 11919 42516 11975 42572
rect 12043 42516 12099 42572
rect 12167 42516 12223 42572
rect 12291 42516 12347 42572
rect 12415 42516 12471 42572
rect 10679 42392 10735 42448
rect 10803 42392 10859 42448
rect 10927 42392 10983 42448
rect 11051 42392 11107 42448
rect 11175 42392 11231 42448
rect 11299 42392 11355 42448
rect 11423 42392 11479 42448
rect 11547 42392 11603 42448
rect 11671 42392 11727 42448
rect 11795 42392 11851 42448
rect 11919 42392 11975 42448
rect 12043 42392 12099 42448
rect 12167 42392 12223 42448
rect 12291 42392 12347 42448
rect 12415 42392 12471 42448
rect 10679 42268 10735 42324
rect 10803 42268 10859 42324
rect 10927 42268 10983 42324
rect 11051 42268 11107 42324
rect 11175 42268 11231 42324
rect 11299 42268 11355 42324
rect 11423 42268 11479 42324
rect 11547 42268 11603 42324
rect 11671 42268 11727 42324
rect 11795 42268 11851 42324
rect 11919 42268 11975 42324
rect 12043 42268 12099 42324
rect 12167 42268 12223 42324
rect 12291 42268 12347 42324
rect 12415 42268 12471 42324
rect 10679 42144 10735 42200
rect 10803 42144 10859 42200
rect 10927 42144 10983 42200
rect 11051 42144 11107 42200
rect 11175 42144 11231 42200
rect 11299 42144 11355 42200
rect 11423 42144 11479 42200
rect 11547 42144 11603 42200
rect 11671 42144 11727 42200
rect 11795 42144 11851 42200
rect 11919 42144 11975 42200
rect 12043 42144 12099 42200
rect 12167 42144 12223 42200
rect 12291 42144 12347 42200
rect 12415 42144 12471 42200
rect 10679 42020 10735 42076
rect 10803 42020 10859 42076
rect 10927 42020 10983 42076
rect 11051 42020 11107 42076
rect 11175 42020 11231 42076
rect 11299 42020 11355 42076
rect 11423 42020 11479 42076
rect 11547 42020 11603 42076
rect 11671 42020 11727 42076
rect 11795 42020 11851 42076
rect 11919 42020 11975 42076
rect 12043 42020 12099 42076
rect 12167 42020 12223 42076
rect 12291 42020 12347 42076
rect 12415 42020 12471 42076
rect 10679 41896 10735 41952
rect 10803 41896 10859 41952
rect 10927 41896 10983 41952
rect 11051 41896 11107 41952
rect 11175 41896 11231 41952
rect 11299 41896 11355 41952
rect 11423 41896 11479 41952
rect 11547 41896 11603 41952
rect 11671 41896 11727 41952
rect 11795 41896 11851 41952
rect 11919 41896 11975 41952
rect 12043 41896 12099 41952
rect 12167 41896 12223 41952
rect 12291 41896 12347 41952
rect 12415 41896 12471 41952
rect 10679 41772 10735 41828
rect 10803 41772 10859 41828
rect 10927 41772 10983 41828
rect 11051 41772 11107 41828
rect 11175 41772 11231 41828
rect 11299 41772 11355 41828
rect 11423 41772 11479 41828
rect 11547 41772 11603 41828
rect 11671 41772 11727 41828
rect 11795 41772 11851 41828
rect 11919 41772 11975 41828
rect 12043 41772 12099 41828
rect 12167 41772 12223 41828
rect 12291 41772 12347 41828
rect 12415 41772 12471 41828
rect 10679 41648 10735 41704
rect 10803 41648 10859 41704
rect 10927 41648 10983 41704
rect 11051 41648 11107 41704
rect 11175 41648 11231 41704
rect 11299 41648 11355 41704
rect 11423 41648 11479 41704
rect 11547 41648 11603 41704
rect 11671 41648 11727 41704
rect 11795 41648 11851 41704
rect 11919 41648 11975 41704
rect 12043 41648 12099 41704
rect 12167 41648 12223 41704
rect 12291 41648 12347 41704
rect 12415 41648 12471 41704
rect 6082 41488 6138 41544
rect 6082 41364 6138 41420
rect 6082 41240 6138 41296
rect 6082 41116 6138 41172
rect 6082 40992 6138 41048
rect 6082 40868 6138 40924
rect 5338 40741 5394 40797
rect 5338 40617 5394 40673
rect 5338 40493 5394 40549
rect 5338 40369 5394 40425
rect 5338 40245 5394 40301
rect 5338 40121 5394 40177
rect 5338 39997 5394 40053
rect 5338 39873 5394 39929
rect 5338 39749 5394 39805
rect 5338 39625 5394 39681
rect 5338 39501 5394 39557
rect 5338 39377 5394 39433
rect 5338 39253 5394 39309
rect 5462 40741 5518 40797
rect 6082 40744 6138 40800
rect 7562 41288 7618 41344
rect 7686 41288 7742 41344
rect 7810 41288 7866 41344
rect 7934 41288 7990 41344
rect 8058 41288 8114 41344
rect 8182 41288 8238 41344
rect 8306 41288 8362 41344
rect 8430 41288 8486 41344
rect 8554 41288 8610 41344
rect 7562 41164 7618 41220
rect 7686 41164 7742 41220
rect 7810 41164 7866 41220
rect 7934 41164 7990 41220
rect 8058 41164 8114 41220
rect 8182 41164 8238 41220
rect 8306 41164 8362 41220
rect 8430 41164 8486 41220
rect 8554 41164 8610 41220
rect 7562 41040 7618 41096
rect 7686 41040 7742 41096
rect 7810 41040 7866 41096
rect 7934 41040 7990 41096
rect 8058 41040 8114 41096
rect 8182 41040 8238 41096
rect 8306 41040 8362 41096
rect 8430 41040 8486 41096
rect 8554 41040 8610 41096
rect 7562 40916 7618 40972
rect 7686 40916 7742 40972
rect 7810 40916 7866 40972
rect 7934 40916 7990 40972
rect 8058 40916 8114 40972
rect 8182 40916 8238 40972
rect 8306 40916 8362 40972
rect 8430 40916 8486 40972
rect 8554 40916 8610 40972
rect 7562 40792 7618 40848
rect 7686 40792 7742 40848
rect 7810 40792 7866 40848
rect 7934 40792 7990 40848
rect 8058 40792 8114 40848
rect 8182 40792 8238 40848
rect 8306 40792 8362 40848
rect 8430 40792 8486 40848
rect 8554 40792 8610 40848
rect 5462 40617 5518 40673
rect 5462 40493 5518 40549
rect 5462 40369 5518 40425
rect 5462 40245 5518 40301
rect 5462 40121 5518 40177
rect 5462 39997 5518 40053
rect 5462 39873 5518 39929
rect 5462 39749 5518 39805
rect 5462 39625 5518 39681
rect 5462 39501 5518 39557
rect 5462 39377 5518 39433
rect 5462 39253 5518 39309
rect 5462 39129 5518 39185
rect 5586 40617 5642 40673
rect 7562 40668 7618 40724
rect 7686 40668 7742 40724
rect 7810 40668 7866 40724
rect 7934 40668 7990 40724
rect 8058 40668 8114 40724
rect 8182 40668 8238 40724
rect 8306 40668 8362 40724
rect 8430 40668 8486 40724
rect 8554 40668 8610 40724
rect 5586 40493 5642 40549
rect 5586 40369 5642 40425
rect 5586 40245 5642 40301
rect 5586 40121 5642 40177
rect 5586 39997 5642 40053
rect 5586 39873 5642 39929
rect 5586 39749 5642 39805
rect 5586 39625 5642 39681
rect 5586 39501 5642 39557
rect 5586 39377 5642 39433
rect 5586 39253 5642 39309
rect 5586 39129 5642 39185
rect 5586 39005 5642 39061
rect 5710 40493 5766 40549
rect 7562 40544 7618 40600
rect 7686 40544 7742 40600
rect 7810 40544 7866 40600
rect 7934 40544 7990 40600
rect 8058 40544 8114 40600
rect 8182 40544 8238 40600
rect 8306 40544 8362 40600
rect 8430 40544 8486 40600
rect 8554 40544 8610 40600
rect 5710 40369 5766 40425
rect 5710 40245 5766 40301
rect 5710 40121 5766 40177
rect 5710 39997 5766 40053
rect 5710 39873 5766 39929
rect 5710 39749 5766 39805
rect 5710 39625 5766 39681
rect 5710 39501 5766 39557
rect 5710 39377 5766 39433
rect 5710 39253 5766 39309
rect 5710 39129 5766 39185
rect 5710 39005 5766 39061
rect 5710 38881 5766 38937
rect 5834 40369 5890 40425
rect 7562 40420 7618 40476
rect 7686 40420 7742 40476
rect 7810 40420 7866 40476
rect 7934 40420 7990 40476
rect 8058 40420 8114 40476
rect 8182 40420 8238 40476
rect 8306 40420 8362 40476
rect 8430 40420 8486 40476
rect 8554 40420 8610 40476
rect 5834 40245 5890 40301
rect 5834 40121 5890 40177
rect 5834 39997 5890 40053
rect 5834 39873 5890 39929
rect 5834 39749 5890 39805
rect 5834 39625 5890 39681
rect 5834 39501 5890 39557
rect 5834 39377 5890 39433
rect 5834 39253 5890 39309
rect 5834 39129 5890 39185
rect 5834 39005 5890 39061
rect 5834 38881 5890 38937
rect 5834 38757 5890 38813
rect 5958 40245 6014 40301
rect 7562 40296 7618 40352
rect 7686 40296 7742 40352
rect 7810 40296 7866 40352
rect 7934 40296 7990 40352
rect 8058 40296 8114 40352
rect 8182 40296 8238 40352
rect 8306 40296 8362 40352
rect 8430 40296 8486 40352
rect 8554 40296 8610 40352
rect 5958 40121 6014 40177
rect 5958 39997 6014 40053
rect 5958 39873 6014 39929
rect 5958 39749 6014 39805
rect 5958 39625 6014 39681
rect 5958 39501 6014 39557
rect 5958 39377 6014 39433
rect 5958 39253 6014 39309
rect 5958 39129 6014 39185
rect 5958 39005 6014 39061
rect 5958 38881 6014 38937
rect 5958 38757 6014 38813
rect 5958 38633 6014 38689
rect 6082 40121 6138 40177
rect 6082 39997 6138 40053
rect 7562 40172 7618 40228
rect 7686 40172 7742 40228
rect 7810 40172 7866 40228
rect 7934 40172 7990 40228
rect 8058 40172 8114 40228
rect 8182 40172 8238 40228
rect 8306 40172 8362 40228
rect 8430 40172 8486 40228
rect 8554 40172 8610 40228
rect 7562 40048 7618 40104
rect 7686 40048 7742 40104
rect 7810 40048 7866 40104
rect 7934 40048 7990 40104
rect 8058 40048 8114 40104
rect 8182 40048 8238 40104
rect 8306 40048 8362 40104
rect 8430 40048 8486 40104
rect 8554 40048 8610 40104
rect 10679 41288 10735 41344
rect 10803 41288 10859 41344
rect 10927 41288 10983 41344
rect 11051 41288 11107 41344
rect 11175 41288 11231 41344
rect 11299 41288 11355 41344
rect 11423 41288 11479 41344
rect 11547 41288 11603 41344
rect 11671 41288 11727 41344
rect 11795 41288 11851 41344
rect 11919 41288 11975 41344
rect 12043 41288 12099 41344
rect 12167 41288 12223 41344
rect 12291 41288 12347 41344
rect 12415 41288 12471 41344
rect 10679 41164 10735 41220
rect 10803 41164 10859 41220
rect 10927 41164 10983 41220
rect 11051 41164 11107 41220
rect 11175 41164 11231 41220
rect 11299 41164 11355 41220
rect 11423 41164 11479 41220
rect 11547 41164 11603 41220
rect 11671 41164 11727 41220
rect 11795 41164 11851 41220
rect 11919 41164 11975 41220
rect 12043 41164 12099 41220
rect 12167 41164 12223 41220
rect 12291 41164 12347 41220
rect 12415 41164 12471 41220
rect 10679 41040 10735 41096
rect 10803 41040 10859 41096
rect 10927 41040 10983 41096
rect 11051 41040 11107 41096
rect 11175 41040 11231 41096
rect 11299 41040 11355 41096
rect 11423 41040 11479 41096
rect 11547 41040 11603 41096
rect 11671 41040 11727 41096
rect 11795 41040 11851 41096
rect 11919 41040 11975 41096
rect 12043 41040 12099 41096
rect 12167 41040 12223 41096
rect 12291 41040 12347 41096
rect 12415 41040 12471 41096
rect 10679 40916 10735 40972
rect 10803 40916 10859 40972
rect 10927 40916 10983 40972
rect 11051 40916 11107 40972
rect 11175 40916 11231 40972
rect 11299 40916 11355 40972
rect 11423 40916 11479 40972
rect 11547 40916 11603 40972
rect 11671 40916 11727 40972
rect 11795 40916 11851 40972
rect 11919 40916 11975 40972
rect 12043 40916 12099 40972
rect 12167 40916 12223 40972
rect 12291 40916 12347 40972
rect 12415 40916 12471 40972
rect 10679 40792 10735 40848
rect 10803 40792 10859 40848
rect 10927 40792 10983 40848
rect 11051 40792 11107 40848
rect 11175 40792 11231 40848
rect 11299 40792 11355 40848
rect 11423 40792 11479 40848
rect 11547 40792 11603 40848
rect 11671 40792 11727 40848
rect 11795 40792 11851 40848
rect 11919 40792 11975 40848
rect 12043 40792 12099 40848
rect 12167 40792 12223 40848
rect 12291 40792 12347 40848
rect 12415 40792 12471 40848
rect 10679 40668 10735 40724
rect 10803 40668 10859 40724
rect 10927 40668 10983 40724
rect 11051 40668 11107 40724
rect 11175 40668 11231 40724
rect 11299 40668 11355 40724
rect 11423 40668 11479 40724
rect 11547 40668 11603 40724
rect 11671 40668 11727 40724
rect 11795 40668 11851 40724
rect 11919 40668 11975 40724
rect 12043 40668 12099 40724
rect 12167 40668 12223 40724
rect 12291 40668 12347 40724
rect 12415 40668 12471 40724
rect 10679 40544 10735 40600
rect 10803 40544 10859 40600
rect 10927 40544 10983 40600
rect 11051 40544 11107 40600
rect 11175 40544 11231 40600
rect 11299 40544 11355 40600
rect 11423 40544 11479 40600
rect 11547 40544 11603 40600
rect 11671 40544 11727 40600
rect 11795 40544 11851 40600
rect 11919 40544 11975 40600
rect 12043 40544 12099 40600
rect 12167 40544 12223 40600
rect 12291 40544 12347 40600
rect 12415 40544 12471 40600
rect 10679 40420 10735 40476
rect 10803 40420 10859 40476
rect 10927 40420 10983 40476
rect 11051 40420 11107 40476
rect 11175 40420 11231 40476
rect 11299 40420 11355 40476
rect 11423 40420 11479 40476
rect 11547 40420 11603 40476
rect 11671 40420 11727 40476
rect 11795 40420 11851 40476
rect 11919 40420 11975 40476
rect 12043 40420 12099 40476
rect 12167 40420 12223 40476
rect 12291 40420 12347 40476
rect 12415 40420 12471 40476
rect 10679 40296 10735 40352
rect 10803 40296 10859 40352
rect 10927 40296 10983 40352
rect 11051 40296 11107 40352
rect 11175 40296 11231 40352
rect 11299 40296 11355 40352
rect 11423 40296 11479 40352
rect 11547 40296 11603 40352
rect 11671 40296 11727 40352
rect 11795 40296 11851 40352
rect 11919 40296 11975 40352
rect 12043 40296 12099 40352
rect 12167 40296 12223 40352
rect 12291 40296 12347 40352
rect 12415 40296 12471 40352
rect 10679 40172 10735 40228
rect 10803 40172 10859 40228
rect 10927 40172 10983 40228
rect 11051 40172 11107 40228
rect 11175 40172 11231 40228
rect 11299 40172 11355 40228
rect 11423 40172 11479 40228
rect 11547 40172 11603 40228
rect 11671 40172 11727 40228
rect 11795 40172 11851 40228
rect 11919 40172 11975 40228
rect 12043 40172 12099 40228
rect 12167 40172 12223 40228
rect 12291 40172 12347 40228
rect 12415 40172 12471 40228
rect 10679 40048 10735 40104
rect 10803 40048 10859 40104
rect 10927 40048 10983 40104
rect 11051 40048 11107 40104
rect 11175 40048 11231 40104
rect 11299 40048 11355 40104
rect 11423 40048 11479 40104
rect 11547 40048 11603 40104
rect 11671 40048 11727 40104
rect 11795 40048 11851 40104
rect 11919 40048 11975 40104
rect 12043 40048 12099 40104
rect 12167 40048 12223 40104
rect 12291 40048 12347 40104
rect 12415 40048 12471 40104
rect 6082 39873 6138 39929
rect 6082 39749 6138 39805
rect 6082 39625 6138 39681
rect 6082 39501 6138 39557
rect 6082 39377 6138 39433
rect 6082 39253 6138 39309
rect 6082 39129 6138 39185
rect 6082 39005 6138 39061
rect 6082 38881 6138 38937
rect 6082 38757 6138 38813
rect 6082 38633 6138 38689
rect 6082 38509 6138 38565
rect 7562 39688 7618 39744
rect 7686 39688 7742 39744
rect 7810 39688 7866 39744
rect 7934 39688 7990 39744
rect 8058 39688 8114 39744
rect 8182 39688 8238 39744
rect 8306 39688 8362 39744
rect 8430 39688 8486 39744
rect 8554 39688 8610 39744
rect 7562 39564 7618 39620
rect 7686 39564 7742 39620
rect 7810 39564 7866 39620
rect 7934 39564 7990 39620
rect 8058 39564 8114 39620
rect 8182 39564 8238 39620
rect 8306 39564 8362 39620
rect 8430 39564 8486 39620
rect 8554 39564 8610 39620
rect 7562 39440 7618 39496
rect 7686 39440 7742 39496
rect 7810 39440 7866 39496
rect 7934 39440 7990 39496
rect 8058 39440 8114 39496
rect 8182 39440 8238 39496
rect 8306 39440 8362 39496
rect 8430 39440 8486 39496
rect 8554 39440 8610 39496
rect 7562 39316 7618 39372
rect 7686 39316 7742 39372
rect 7810 39316 7866 39372
rect 7934 39316 7990 39372
rect 8058 39316 8114 39372
rect 8182 39316 8238 39372
rect 8306 39316 8362 39372
rect 8430 39316 8486 39372
rect 8554 39316 8610 39372
rect 7562 39192 7618 39248
rect 7686 39192 7742 39248
rect 7810 39192 7866 39248
rect 7934 39192 7990 39248
rect 8058 39192 8114 39248
rect 8182 39192 8238 39248
rect 8306 39192 8362 39248
rect 8430 39192 8486 39248
rect 8554 39192 8610 39248
rect 7562 39068 7618 39124
rect 7686 39068 7742 39124
rect 7810 39068 7866 39124
rect 7934 39068 7990 39124
rect 8058 39068 8114 39124
rect 8182 39068 8238 39124
rect 8306 39068 8362 39124
rect 8430 39068 8486 39124
rect 8554 39068 8610 39124
rect 7562 38944 7618 39000
rect 7686 38944 7742 39000
rect 7810 38944 7866 39000
rect 7934 38944 7990 39000
rect 8058 38944 8114 39000
rect 8182 38944 8238 39000
rect 8306 38944 8362 39000
rect 8430 38944 8486 39000
rect 8554 38944 8610 39000
rect 7562 38820 7618 38876
rect 7686 38820 7742 38876
rect 7810 38820 7866 38876
rect 7934 38820 7990 38876
rect 8058 38820 8114 38876
rect 8182 38820 8238 38876
rect 8306 38820 8362 38876
rect 8430 38820 8486 38876
rect 8554 38820 8610 38876
rect 7562 38696 7618 38752
rect 7686 38696 7742 38752
rect 7810 38696 7866 38752
rect 7934 38696 7990 38752
rect 8058 38696 8114 38752
rect 8182 38696 8238 38752
rect 8306 38696 8362 38752
rect 8430 38696 8486 38752
rect 8554 38696 8610 38752
rect 7562 38572 7618 38628
rect 7686 38572 7742 38628
rect 7810 38572 7866 38628
rect 7934 38572 7990 38628
rect 8058 38572 8114 38628
rect 8182 38572 8238 38628
rect 8306 38572 8362 38628
rect 8430 38572 8486 38628
rect 8554 38572 8610 38628
rect 7562 38448 7618 38504
rect 7686 38448 7742 38504
rect 7810 38448 7866 38504
rect 7934 38448 7990 38504
rect 8058 38448 8114 38504
rect 8182 38448 8238 38504
rect 8306 38448 8362 38504
rect 8430 38448 8486 38504
rect 8554 38448 8610 38504
rect 10679 39688 10735 39744
rect 10803 39688 10859 39744
rect 10927 39688 10983 39744
rect 11051 39688 11107 39744
rect 11175 39688 11231 39744
rect 11299 39688 11355 39744
rect 11423 39688 11479 39744
rect 11547 39688 11603 39744
rect 11671 39688 11727 39744
rect 11795 39688 11851 39744
rect 11919 39688 11975 39744
rect 12043 39688 12099 39744
rect 12167 39688 12223 39744
rect 12291 39688 12347 39744
rect 12415 39688 12471 39744
rect 10679 39564 10735 39620
rect 10803 39564 10859 39620
rect 10927 39564 10983 39620
rect 11051 39564 11107 39620
rect 11175 39564 11231 39620
rect 11299 39564 11355 39620
rect 11423 39564 11479 39620
rect 11547 39564 11603 39620
rect 11671 39564 11727 39620
rect 11795 39564 11851 39620
rect 11919 39564 11975 39620
rect 12043 39564 12099 39620
rect 12167 39564 12223 39620
rect 12291 39564 12347 39620
rect 12415 39564 12471 39620
rect 10679 39440 10735 39496
rect 10803 39440 10859 39496
rect 10927 39440 10983 39496
rect 11051 39440 11107 39496
rect 11175 39440 11231 39496
rect 11299 39440 11355 39496
rect 11423 39440 11479 39496
rect 11547 39440 11603 39496
rect 11671 39440 11727 39496
rect 11795 39440 11851 39496
rect 11919 39440 11975 39496
rect 12043 39440 12099 39496
rect 12167 39440 12223 39496
rect 12291 39440 12347 39496
rect 12415 39440 12471 39496
rect 10679 39316 10735 39372
rect 10803 39316 10859 39372
rect 10927 39316 10983 39372
rect 11051 39316 11107 39372
rect 11175 39316 11231 39372
rect 11299 39316 11355 39372
rect 11423 39316 11479 39372
rect 11547 39316 11603 39372
rect 11671 39316 11727 39372
rect 11795 39316 11851 39372
rect 11919 39316 11975 39372
rect 12043 39316 12099 39372
rect 12167 39316 12223 39372
rect 12291 39316 12347 39372
rect 12415 39316 12471 39372
rect 10679 39192 10735 39248
rect 10803 39192 10859 39248
rect 10927 39192 10983 39248
rect 11051 39192 11107 39248
rect 11175 39192 11231 39248
rect 11299 39192 11355 39248
rect 11423 39192 11479 39248
rect 11547 39192 11603 39248
rect 11671 39192 11727 39248
rect 11795 39192 11851 39248
rect 11919 39192 11975 39248
rect 12043 39192 12099 39248
rect 12167 39192 12223 39248
rect 12291 39192 12347 39248
rect 12415 39192 12471 39248
rect 10679 39068 10735 39124
rect 10803 39068 10859 39124
rect 10927 39068 10983 39124
rect 11051 39068 11107 39124
rect 11175 39068 11231 39124
rect 11299 39068 11355 39124
rect 11423 39068 11479 39124
rect 11547 39068 11603 39124
rect 11671 39068 11727 39124
rect 11795 39068 11851 39124
rect 11919 39068 11975 39124
rect 12043 39068 12099 39124
rect 12167 39068 12223 39124
rect 12291 39068 12347 39124
rect 12415 39068 12471 39124
rect 10679 38944 10735 39000
rect 10803 38944 10859 39000
rect 10927 38944 10983 39000
rect 11051 38944 11107 39000
rect 11175 38944 11231 39000
rect 11299 38944 11355 39000
rect 11423 38944 11479 39000
rect 11547 38944 11603 39000
rect 11671 38944 11727 39000
rect 11795 38944 11851 39000
rect 11919 38944 11975 39000
rect 12043 38944 12099 39000
rect 12167 38944 12223 39000
rect 12291 38944 12347 39000
rect 12415 38944 12471 39000
rect 10679 38820 10735 38876
rect 10803 38820 10859 38876
rect 10927 38820 10983 38876
rect 11051 38820 11107 38876
rect 11175 38820 11231 38876
rect 11299 38820 11355 38876
rect 11423 38820 11479 38876
rect 11547 38820 11603 38876
rect 11671 38820 11727 38876
rect 11795 38820 11851 38876
rect 11919 38820 11975 38876
rect 12043 38820 12099 38876
rect 12167 38820 12223 38876
rect 12291 38820 12347 38876
rect 12415 38820 12471 38876
rect 10679 38696 10735 38752
rect 10803 38696 10859 38752
rect 10927 38696 10983 38752
rect 11051 38696 11107 38752
rect 11175 38696 11231 38752
rect 11299 38696 11355 38752
rect 11423 38696 11479 38752
rect 11547 38696 11603 38752
rect 11671 38696 11727 38752
rect 11795 38696 11851 38752
rect 11919 38696 11975 38752
rect 12043 38696 12099 38752
rect 12167 38696 12223 38752
rect 12291 38696 12347 38752
rect 12415 38696 12471 38752
rect 10679 38572 10735 38628
rect 10803 38572 10859 38628
rect 10927 38572 10983 38628
rect 11051 38572 11107 38628
rect 11175 38572 11231 38628
rect 11299 38572 11355 38628
rect 11423 38572 11479 38628
rect 11547 38572 11603 38628
rect 11671 38572 11727 38628
rect 11795 38572 11851 38628
rect 11919 38572 11975 38628
rect 12043 38572 12099 38628
rect 12167 38572 12223 38628
rect 12291 38572 12347 38628
rect 12415 38572 12471 38628
rect 10679 38448 10735 38504
rect 10803 38448 10859 38504
rect 10927 38448 10983 38504
rect 11051 38448 11107 38504
rect 11175 38448 11231 38504
rect 11299 38448 11355 38504
rect 11423 38448 11479 38504
rect 11547 38448 11603 38504
rect 11671 38448 11727 38504
rect 11795 38448 11851 38504
rect 11919 38448 11975 38504
rect 12043 38448 12099 38504
rect 12167 38448 12223 38504
rect 12291 38448 12347 38504
rect 12415 38448 12471 38504
rect 2527 36944 2583 37000
rect 2527 36820 2583 36876
rect 2527 36696 2583 36752
rect 2527 36572 2583 36628
rect 2527 36448 2583 36504
rect 2527 36324 2583 36380
rect 2527 36200 2583 36256
rect 2527 36076 2583 36132
rect 2527 35952 2583 36008
rect 2527 35828 2583 35884
rect 2527 35704 2583 35760
rect 2527 35580 2583 35636
rect 2527 35456 2583 35512
rect 2527 35332 2583 35388
rect 2527 35208 2583 35264
rect 2527 35084 2583 35140
rect 2527 34960 2583 35016
rect 2527 34836 2583 34892
rect 2527 34712 2583 34768
rect 2527 34588 2583 34644
rect 2527 34464 2583 34520
rect 2527 34340 2583 34396
rect 2527 34216 2583 34272
rect 2527 34092 2583 34148
rect 2527 33968 2583 34024
rect 2527 33844 2583 33900
rect 1155 33710 1211 33766
rect 2527 33720 2583 33776
rect 1155 33586 1211 33642
rect 1155 33462 1211 33518
rect 1155 33338 1211 33394
rect 1155 33214 1211 33270
rect 1155 33090 1211 33146
rect 1155 32966 1211 33022
rect 1155 32842 1211 32898
rect 1155 32718 1211 32774
rect 1155 32594 1211 32650
rect 1155 32470 1211 32526
rect 1155 32346 1211 32402
rect 1155 32222 1211 32278
rect 1155 32098 1211 32154
rect 1155 31974 1211 32030
rect 1155 31850 1211 31906
rect 1155 31726 1211 31782
rect 1155 31602 1211 31658
rect 1155 31478 1211 31534
rect 1155 31354 1211 31410
rect 1155 31230 1211 31286
rect 1155 31106 1211 31162
rect 1155 30982 1211 31038
rect 1155 30858 1211 30914
rect 1155 30734 1211 30790
rect 1155 30610 1211 30666
rect 1155 30486 1211 30542
rect 1155 30362 1211 30418
rect 1155 30238 1211 30294
rect 1155 30114 1211 30170
rect 1155 29990 1211 30046
rect 1155 29866 1211 29922
rect 1155 29742 1211 29798
rect 1279 33586 1335 33642
rect 2527 33596 2583 33652
rect 1279 33462 1335 33518
rect 1279 33338 1335 33394
rect 1279 33214 1335 33270
rect 1279 33090 1335 33146
rect 1279 32966 1335 33022
rect 1279 32842 1335 32898
rect 1279 32718 1335 32774
rect 1279 32594 1335 32650
rect 1279 32470 1335 32526
rect 1279 32346 1335 32402
rect 1279 32222 1335 32278
rect 1279 32098 1335 32154
rect 1279 31974 1335 32030
rect 1279 31850 1335 31906
rect 1279 31726 1335 31782
rect 1279 31602 1335 31658
rect 1279 31478 1335 31534
rect 1279 31354 1335 31410
rect 1279 31230 1335 31286
rect 1279 31106 1335 31162
rect 1279 30982 1335 31038
rect 1279 30858 1335 30914
rect 1279 30734 1335 30790
rect 1279 30610 1335 30666
rect 1279 30486 1335 30542
rect 1279 30362 1335 30418
rect 1279 30238 1335 30294
rect 1279 30114 1335 30170
rect 1279 29990 1335 30046
rect 1279 29866 1335 29922
rect 1279 29742 1335 29798
rect 1279 29618 1335 29674
rect 1403 33462 1459 33518
rect 2527 33472 2583 33528
rect 1403 33338 1459 33394
rect 1403 33214 1459 33270
rect 1403 33090 1459 33146
rect 1403 32966 1459 33022
rect 1403 32842 1459 32898
rect 1403 32718 1459 32774
rect 1403 32594 1459 32650
rect 1403 32470 1459 32526
rect 1403 32346 1459 32402
rect 1403 32222 1459 32278
rect 1403 32098 1459 32154
rect 1403 31974 1459 32030
rect 1403 31850 1459 31906
rect 1403 31726 1459 31782
rect 1403 31602 1459 31658
rect 1403 31478 1459 31534
rect 1403 31354 1459 31410
rect 1403 31230 1459 31286
rect 1403 31106 1459 31162
rect 1403 30982 1459 31038
rect 1403 30858 1459 30914
rect 1403 30734 1459 30790
rect 1403 30610 1459 30666
rect 1403 30486 1459 30542
rect 1403 30362 1459 30418
rect 1403 30238 1459 30294
rect 1403 30114 1459 30170
rect 1403 29990 1459 30046
rect 1403 29866 1459 29922
rect 1403 29742 1459 29798
rect 1403 29618 1459 29674
rect 1403 29494 1459 29550
rect 1527 33338 1583 33394
rect 2527 33348 2583 33404
rect 1527 33214 1583 33270
rect 1527 33090 1583 33146
rect 1527 32966 1583 33022
rect 1527 32842 1583 32898
rect 1527 32718 1583 32774
rect 1527 32594 1583 32650
rect 1527 32470 1583 32526
rect 1527 32346 1583 32402
rect 1527 32222 1583 32278
rect 1527 32098 1583 32154
rect 1527 31974 1583 32030
rect 1527 31850 1583 31906
rect 1527 31726 1583 31782
rect 1527 31602 1583 31658
rect 1527 31478 1583 31534
rect 1527 31354 1583 31410
rect 1527 31230 1583 31286
rect 1527 31106 1583 31162
rect 1527 30982 1583 31038
rect 1527 30858 1583 30914
rect 1527 30734 1583 30790
rect 1527 30610 1583 30666
rect 1527 30486 1583 30542
rect 1527 30362 1583 30418
rect 1527 30238 1583 30294
rect 1527 30114 1583 30170
rect 1527 29990 1583 30046
rect 1527 29866 1583 29922
rect 1527 29742 1583 29798
rect 1527 29618 1583 29674
rect 1527 29494 1583 29550
rect 1527 29370 1583 29426
rect 1651 33214 1707 33270
rect 2527 33224 2583 33280
rect 1651 33090 1707 33146
rect 1651 32966 1707 33022
rect 1651 32842 1707 32898
rect 1651 32718 1707 32774
rect 1651 32594 1707 32650
rect 1651 32470 1707 32526
rect 1651 32346 1707 32402
rect 1651 32222 1707 32278
rect 1651 32098 1707 32154
rect 1651 31974 1707 32030
rect 1651 31850 1707 31906
rect 1651 31726 1707 31782
rect 1651 31602 1707 31658
rect 1651 31478 1707 31534
rect 1651 31354 1707 31410
rect 1651 31230 1707 31286
rect 1651 31106 1707 31162
rect 1651 30982 1707 31038
rect 1651 30858 1707 30914
rect 1651 30734 1707 30790
rect 1651 30610 1707 30666
rect 1651 30486 1707 30542
rect 1651 30362 1707 30418
rect 1651 30238 1707 30294
rect 1651 30114 1707 30170
rect 1651 29990 1707 30046
rect 1651 29866 1707 29922
rect 1651 29742 1707 29798
rect 1651 29618 1707 29674
rect 1651 29494 1707 29550
rect 1651 29370 1707 29426
rect 1127 29251 1183 29307
rect 1651 29246 1707 29302
rect 1775 33090 1831 33146
rect 2527 33100 2583 33156
rect 1775 32966 1831 33022
rect 1775 32842 1831 32898
rect 1775 32718 1831 32774
rect 1775 32594 1831 32650
rect 1775 32470 1831 32526
rect 1775 32346 1831 32402
rect 1775 32222 1831 32278
rect 1775 32098 1831 32154
rect 1775 31974 1831 32030
rect 1775 31850 1831 31906
rect 1775 31726 1831 31782
rect 1775 31602 1831 31658
rect 1775 31478 1831 31534
rect 1775 31354 1831 31410
rect 1775 31230 1831 31286
rect 1775 31106 1831 31162
rect 1775 30982 1831 31038
rect 1775 30858 1831 30914
rect 1775 30734 1831 30790
rect 1775 30610 1831 30666
rect 1775 30486 1831 30542
rect 1775 30362 1831 30418
rect 1775 30238 1831 30294
rect 1775 30114 1831 30170
rect 1775 29990 1831 30046
rect 1775 29866 1831 29922
rect 1775 29742 1831 29798
rect 1775 29618 1831 29674
rect 1775 29494 1831 29550
rect 1775 29370 1831 29426
rect 1775 29246 1831 29302
rect 1127 29127 1183 29183
rect 1127 29003 1183 29059
rect 1127 28879 1183 28935
rect 1127 28755 1183 28811
rect 1127 28631 1183 28687
rect 1127 28507 1183 28563
rect 1127 28383 1183 28439
rect 1127 28259 1183 28315
rect 1127 28135 1183 28191
rect 1127 28011 1183 28067
rect 1127 27887 1183 27943
rect 1127 27763 1183 27819
rect 1127 27639 1183 27695
rect 1127 27515 1183 27571
rect 1251 29127 1307 29183
rect 1775 29122 1831 29178
rect 1899 32966 1955 33022
rect 2527 32976 2583 33032
rect 2651 36820 2707 36876
rect 2651 36696 2707 36752
rect 2651 36572 2707 36628
rect 2651 36448 2707 36504
rect 2651 36324 2707 36380
rect 2651 36200 2707 36256
rect 2651 36076 2707 36132
rect 2651 35952 2707 36008
rect 2651 35828 2707 35884
rect 2651 35704 2707 35760
rect 2651 35580 2707 35636
rect 2651 35456 2707 35512
rect 2651 35332 2707 35388
rect 2651 35208 2707 35264
rect 2651 35084 2707 35140
rect 2651 34960 2707 35016
rect 2651 34836 2707 34892
rect 2651 34712 2707 34768
rect 2651 34588 2707 34644
rect 2651 34464 2707 34520
rect 2651 34340 2707 34396
rect 2651 34216 2707 34272
rect 2651 34092 2707 34148
rect 2651 33968 2707 34024
rect 2651 33844 2707 33900
rect 2651 33720 2707 33776
rect 2651 33596 2707 33652
rect 2651 33472 2707 33528
rect 2651 33348 2707 33404
rect 2651 33224 2707 33280
rect 2651 33100 2707 33156
rect 2651 32976 2707 33032
rect 1899 32842 1955 32898
rect 1899 32718 1955 32774
rect 1899 32594 1955 32650
rect 1899 32470 1955 32526
rect 1899 32346 1955 32402
rect 1899 32222 1955 32278
rect 1899 32098 1955 32154
rect 1899 31974 1955 32030
rect 1899 31850 1955 31906
rect 1899 31726 1955 31782
rect 1899 31602 1955 31658
rect 1899 31478 1955 31534
rect 1899 31354 1955 31410
rect 1899 31230 1955 31286
rect 1899 31106 1955 31162
rect 1899 30982 1955 31038
rect 1899 30858 1955 30914
rect 1899 30734 1955 30790
rect 1899 30610 1955 30666
rect 1899 30486 1955 30542
rect 1899 30362 1955 30418
rect 1899 30238 1955 30294
rect 1899 30114 1955 30170
rect 1899 29990 1955 30046
rect 1899 29866 1955 29922
rect 1899 29742 1955 29798
rect 1899 29618 1955 29674
rect 1899 29494 1955 29550
rect 1899 29370 1955 29426
rect 1899 29246 1955 29302
rect 1899 29122 1955 29178
rect 1251 29003 1307 29059
rect 1251 28879 1307 28935
rect 1251 28755 1307 28811
rect 1251 28631 1307 28687
rect 1251 28507 1307 28563
rect 1251 28383 1307 28439
rect 1251 28259 1307 28315
rect 1251 28135 1307 28191
rect 1251 28011 1307 28067
rect 1251 27887 1307 27943
rect 1251 27763 1307 27819
rect 1251 27639 1307 27695
rect 1251 27515 1307 27571
rect 1251 27391 1307 27447
rect 1375 29003 1431 29059
rect 1899 28998 1955 29054
rect 2023 32842 2079 32898
rect 2651 32852 2707 32908
rect 2775 36696 2831 36752
rect 2775 36572 2831 36628
rect 2775 36448 2831 36504
rect 2775 36324 2831 36380
rect 2775 36200 2831 36256
rect 2775 36076 2831 36132
rect 2775 35952 2831 36008
rect 2775 35828 2831 35884
rect 2775 35704 2831 35760
rect 2775 35580 2831 35636
rect 2775 35456 2831 35512
rect 2775 35332 2831 35388
rect 2775 35208 2831 35264
rect 2775 35084 2831 35140
rect 2775 34960 2831 35016
rect 2775 34836 2831 34892
rect 2775 34712 2831 34768
rect 2775 34588 2831 34644
rect 2775 34464 2831 34520
rect 2775 34340 2831 34396
rect 2775 34216 2831 34272
rect 2775 34092 2831 34148
rect 2775 33968 2831 34024
rect 2775 33844 2831 33900
rect 2775 33720 2831 33776
rect 2775 33596 2831 33652
rect 2775 33472 2831 33528
rect 2775 33348 2831 33404
rect 2775 33224 2831 33280
rect 2775 33100 2831 33156
rect 2775 32976 2831 33032
rect 2775 32852 2831 32908
rect 2023 32718 2079 32774
rect 2775 32728 2831 32784
rect 2899 36572 2955 36628
rect 2899 36448 2955 36504
rect 2899 36324 2955 36380
rect 2899 36200 2955 36256
rect 2899 36076 2955 36132
rect 2899 35952 2955 36008
rect 2899 35828 2955 35884
rect 2899 35704 2955 35760
rect 2899 35580 2955 35636
rect 2899 35456 2955 35512
rect 2899 35332 2955 35388
rect 2899 35208 2955 35264
rect 2899 35084 2955 35140
rect 2899 34960 2955 35016
rect 2899 34836 2955 34892
rect 2899 34712 2955 34768
rect 2899 34588 2955 34644
rect 2899 34464 2955 34520
rect 2899 34340 2955 34396
rect 2899 34216 2955 34272
rect 2899 34092 2955 34148
rect 2899 33968 2955 34024
rect 2899 33844 2955 33900
rect 2899 33720 2955 33776
rect 2899 33596 2955 33652
rect 2899 33472 2955 33528
rect 2899 33348 2955 33404
rect 2899 33224 2955 33280
rect 2899 33100 2955 33156
rect 2899 32976 2955 33032
rect 2899 32852 2955 32908
rect 2899 32728 2955 32784
rect 2023 32594 2079 32650
rect 2899 32604 2955 32660
rect 3023 36448 3079 36504
rect 3023 36324 3079 36380
rect 3023 36200 3079 36256
rect 3023 36076 3079 36132
rect 3023 35952 3079 36008
rect 3023 35828 3079 35884
rect 3023 35704 3079 35760
rect 3023 35580 3079 35636
rect 3023 35456 3079 35512
rect 3023 35332 3079 35388
rect 3023 35208 3079 35264
rect 3023 35084 3079 35140
rect 3023 34960 3079 35016
rect 3023 34836 3079 34892
rect 3023 34712 3079 34768
rect 3023 34588 3079 34644
rect 3023 34464 3079 34520
rect 3023 34340 3079 34396
rect 3023 34216 3079 34272
rect 3023 34092 3079 34148
rect 3023 33968 3079 34024
rect 3023 33844 3079 33900
rect 3023 33720 3079 33776
rect 3023 33596 3079 33652
rect 3023 33472 3079 33528
rect 3023 33348 3079 33404
rect 3023 33224 3079 33280
rect 3023 33100 3079 33156
rect 3023 32976 3079 33032
rect 3023 32852 3079 32908
rect 3023 32728 3079 32784
rect 3023 32604 3079 32660
rect 2023 32470 2079 32526
rect 3023 32480 3079 32536
rect 3147 36324 3203 36380
rect 3147 36200 3203 36256
rect 3147 36076 3203 36132
rect 3147 35952 3203 36008
rect 3147 35828 3203 35884
rect 3147 35704 3203 35760
rect 3147 35580 3203 35636
rect 3147 35456 3203 35512
rect 3147 35332 3203 35388
rect 3147 35208 3203 35264
rect 3147 35084 3203 35140
rect 3147 34960 3203 35016
rect 3147 34836 3203 34892
rect 3147 34712 3203 34768
rect 3147 34588 3203 34644
rect 3147 34464 3203 34520
rect 3147 34340 3203 34396
rect 3147 34216 3203 34272
rect 3147 34092 3203 34148
rect 3147 33968 3203 34024
rect 3147 33844 3203 33900
rect 3147 33720 3203 33776
rect 3147 33596 3203 33652
rect 3147 33472 3203 33528
rect 3147 33348 3203 33404
rect 3147 33224 3203 33280
rect 3147 33100 3203 33156
rect 3147 32976 3203 33032
rect 3147 32852 3203 32908
rect 3147 32728 3203 32784
rect 3147 32604 3203 32660
rect 3147 32480 3203 32536
rect 2023 32346 2079 32402
rect 3147 32356 3203 32412
rect 3271 36200 3327 36256
rect 3271 36076 3327 36132
rect 3271 35952 3327 36008
rect 3271 35828 3327 35884
rect 3271 35704 3327 35760
rect 3271 35580 3327 35636
rect 3271 35456 3327 35512
rect 3271 35332 3327 35388
rect 3271 35208 3327 35264
rect 3271 35084 3327 35140
rect 3271 34960 3327 35016
rect 3271 34836 3327 34892
rect 3271 34712 3327 34768
rect 3271 34588 3327 34644
rect 3271 34464 3327 34520
rect 3271 34340 3327 34396
rect 3271 34216 3327 34272
rect 3271 34092 3327 34148
rect 3271 33968 3327 34024
rect 3271 33844 3327 33900
rect 3271 33720 3327 33776
rect 3271 33596 3327 33652
rect 3271 33472 3327 33528
rect 3271 33348 3327 33404
rect 3271 33224 3327 33280
rect 3271 33100 3327 33156
rect 3271 32976 3327 33032
rect 3271 32852 3327 32908
rect 3271 32728 3327 32784
rect 3271 32604 3327 32660
rect 3271 32480 3327 32536
rect 3271 32356 3327 32412
rect 2023 32222 2079 32278
rect 3271 32232 3327 32288
rect 3395 36076 3451 36132
rect 3395 35952 3451 36008
rect 3395 35828 3451 35884
rect 3395 35704 3451 35760
rect 3395 35580 3451 35636
rect 3395 35456 3451 35512
rect 3395 35332 3451 35388
rect 3395 35208 3451 35264
rect 3395 35084 3451 35140
rect 3395 34960 3451 35016
rect 3395 34836 3451 34892
rect 3395 34712 3451 34768
rect 3395 34588 3451 34644
rect 3395 34464 3451 34520
rect 3395 34340 3451 34396
rect 3395 34216 3451 34272
rect 3395 34092 3451 34148
rect 3395 33968 3451 34024
rect 3395 33844 3451 33900
rect 3395 33720 3451 33776
rect 3395 33596 3451 33652
rect 3395 33472 3451 33528
rect 3395 33348 3451 33404
rect 3395 33224 3451 33280
rect 3395 33100 3451 33156
rect 3395 32976 3451 33032
rect 3395 32852 3451 32908
rect 3395 32728 3451 32784
rect 3395 32604 3451 32660
rect 3395 32480 3451 32536
rect 3395 32356 3451 32412
rect 3395 32232 3451 32288
rect 2023 32098 2079 32154
rect 3395 32108 3451 32164
rect 3519 35890 3575 35946
rect 3519 35766 3575 35822
rect 3519 35642 3575 35698
rect 3519 35518 3575 35574
rect 3519 35394 3575 35450
rect 3519 35270 3575 35326
rect 3519 35146 3575 35202
rect 3519 35022 3575 35078
rect 3519 34898 3575 34954
rect 3519 34774 3575 34830
rect 3519 34650 3575 34706
rect 3519 34526 3575 34582
rect 3519 34402 3575 34458
rect 3519 34278 3575 34334
rect 3519 34154 3575 34210
rect 3519 34030 3575 34086
rect 3519 33906 3575 33962
rect 3519 33782 3575 33838
rect 3519 33658 3575 33714
rect 3519 33534 3575 33590
rect 3519 33410 3575 33466
rect 3519 33286 3575 33342
rect 3519 33162 3575 33218
rect 3519 33038 3575 33094
rect 3519 32914 3575 32970
rect 3519 32790 3575 32846
rect 3519 32666 3575 32722
rect 3519 32542 3575 32598
rect 3519 32418 3575 32474
rect 3519 32294 3575 32350
rect 3519 32170 3575 32226
rect 3519 32046 3575 32102
rect 3643 35757 3699 35813
rect 3643 35633 3699 35689
rect 3643 35509 3699 35565
rect 3643 35385 3699 35441
rect 3643 35261 3699 35317
rect 3643 35137 3699 35193
rect 3643 35013 3699 35069
rect 3643 34889 3699 34945
rect 3643 34765 3699 34821
rect 3643 34641 3699 34697
rect 3643 34517 3699 34573
rect 3643 34393 3699 34449
rect 3643 34269 3699 34325
rect 3643 34145 3699 34201
rect 3643 34021 3699 34077
rect 3643 33897 3699 33953
rect 3643 33773 3699 33829
rect 3643 33649 3699 33705
rect 3643 33525 3699 33581
rect 3643 33401 3699 33457
rect 3643 33277 3699 33333
rect 3643 33153 3699 33209
rect 3643 33029 3699 33085
rect 3643 32905 3699 32961
rect 3643 32781 3699 32837
rect 3643 32657 3699 32713
rect 3643 32533 3699 32589
rect 3643 32409 3699 32465
rect 3643 32285 3699 32341
rect 3643 32161 3699 32217
rect 3643 32037 3699 32093
rect 3767 35654 3823 35710
rect 3767 35530 3823 35586
rect 3767 35406 3823 35462
rect 3767 35282 3823 35338
rect 3767 35158 3823 35214
rect 3767 35034 3823 35090
rect 3767 34910 3823 34966
rect 3767 34786 3823 34842
rect 3767 34662 3823 34718
rect 3767 34538 3823 34594
rect 3767 34414 3823 34470
rect 3767 34290 3823 34346
rect 3767 34166 3823 34222
rect 3767 34042 3823 34098
rect 3767 33918 3823 33974
rect 3767 33794 3823 33850
rect 3767 33670 3823 33726
rect 3767 33546 3823 33602
rect 3767 33422 3823 33478
rect 3767 33298 3823 33354
rect 3767 33174 3823 33230
rect 3767 33050 3823 33106
rect 3767 32926 3823 32982
rect 3767 32802 3823 32858
rect 3767 32678 3823 32734
rect 3767 32554 3823 32610
rect 3767 32430 3823 32486
rect 3767 32306 3823 32362
rect 3767 32182 3823 32238
rect 3767 32058 3823 32114
rect 3891 35550 3947 35606
rect 3891 35426 3947 35482
rect 3891 35302 3947 35358
rect 3891 35178 3947 35234
rect 3891 35054 3947 35110
rect 3891 34930 3947 34986
rect 3891 34806 3947 34862
rect 3891 34682 3947 34738
rect 3891 34558 3947 34614
rect 3891 34434 3947 34490
rect 3891 34310 3947 34366
rect 3891 34186 3947 34242
rect 3891 34062 3947 34118
rect 3891 33938 3947 33994
rect 3891 33814 3947 33870
rect 3891 33690 3947 33746
rect 3891 33566 3947 33622
rect 3891 33442 3947 33498
rect 3891 33318 3947 33374
rect 3891 33194 3947 33250
rect 3891 33070 3947 33126
rect 3891 32946 3947 33002
rect 3891 32822 3947 32878
rect 3891 32698 3947 32754
rect 3891 32574 3947 32630
rect 3891 32450 3947 32506
rect 3891 32326 3947 32382
rect 3891 32202 3947 32258
rect 3891 32078 3947 32134
rect 4015 35479 4071 35535
rect 4015 35355 4071 35411
rect 4015 35231 4071 35287
rect 4015 35107 4071 35163
rect 4015 34983 4071 35039
rect 4015 34859 4071 34915
rect 4015 34735 4071 34791
rect 4015 34611 4071 34667
rect 4015 34487 4071 34543
rect 4015 34363 4071 34419
rect 4015 34239 4071 34295
rect 4015 34115 4071 34171
rect 4015 33991 4071 34047
rect 4015 33867 4071 33923
rect 4015 33743 4071 33799
rect 4015 33619 4071 33675
rect 4015 33495 4071 33551
rect 4015 33371 4071 33427
rect 4015 33247 4071 33303
rect 4015 33123 4071 33179
rect 4015 32999 4071 33055
rect 4015 32875 4071 32931
rect 4015 32751 4071 32807
rect 4015 32627 4071 32683
rect 4015 32503 4071 32559
rect 4015 32379 4071 32435
rect 4015 32255 4071 32311
rect 4015 32131 4071 32187
rect 2023 31974 2079 32030
rect 4015 32007 4071 32063
rect 4139 35361 4195 35417
rect 4139 35237 4195 35293
rect 14767 36570 14823 36572
rect 14767 36518 14769 36570
rect 14769 36518 14821 36570
rect 14821 36518 14823 36570
rect 14767 36462 14823 36518
rect 14767 36410 14769 36462
rect 14769 36410 14821 36462
rect 14821 36410 14823 36462
rect 14767 36354 14823 36410
rect 14767 36302 14769 36354
rect 14769 36302 14821 36354
rect 14821 36302 14823 36354
rect 14767 36246 14823 36302
rect 14767 36194 14769 36246
rect 14769 36194 14821 36246
rect 14821 36194 14823 36246
rect 14767 36138 14823 36194
rect 14767 36086 14769 36138
rect 14769 36086 14821 36138
rect 14821 36086 14823 36138
rect 14767 36030 14823 36086
rect 14767 35978 14769 36030
rect 14769 35978 14821 36030
rect 14821 35978 14823 36030
rect 14767 35922 14823 35978
rect 14767 35870 14769 35922
rect 14769 35870 14821 35922
rect 14821 35870 14823 35922
rect 14767 35814 14823 35870
rect 14767 35762 14769 35814
rect 14769 35762 14821 35814
rect 14821 35762 14823 35814
rect 14767 35706 14823 35762
rect 14767 35654 14769 35706
rect 14769 35654 14821 35706
rect 14821 35654 14823 35706
rect 14767 35598 14823 35654
rect 14767 35546 14769 35598
rect 14769 35546 14821 35598
rect 14821 35546 14823 35598
rect 14767 35490 14823 35546
rect 14767 35438 14769 35490
rect 14769 35438 14821 35490
rect 14821 35438 14823 35490
rect 14767 35382 14823 35438
rect 14767 35330 14769 35382
rect 14769 35330 14821 35382
rect 14821 35330 14823 35382
rect 14767 35274 14823 35330
rect 14767 35222 14769 35274
rect 14769 35222 14821 35274
rect 14821 35222 14823 35274
rect 14767 35220 14823 35222
rect 4139 35113 4195 35169
rect 4139 34989 4195 35045
rect 4139 34865 4195 34921
rect 4139 34741 4195 34797
rect 4139 34617 4195 34673
rect 4139 34493 4195 34549
rect 4139 34369 4195 34425
rect 4139 34245 4195 34301
rect 4139 34121 4195 34177
rect 4139 33997 4195 34053
rect 4139 33873 4195 33929
rect 4139 33749 4195 33805
rect 4139 33625 4195 33681
rect 4139 33501 4195 33557
rect 4139 33377 4195 33433
rect 4139 33253 4195 33309
rect 4139 33129 4195 33185
rect 4139 33005 4195 33061
rect 4139 32881 4195 32937
rect 4139 32757 4195 32813
rect 4139 32633 4195 32689
rect 4139 32509 4195 32565
rect 4139 32385 4195 32441
rect 4139 32261 4195 32317
rect 4139 32137 4195 32193
rect 4139 32013 4195 32069
rect 6368 34894 6424 34950
rect 6492 34894 6548 34950
rect 6616 34894 6672 34950
rect 6740 34894 6796 34950
rect 6864 34894 6920 34950
rect 6988 34894 7044 34950
rect 7112 34894 7168 34950
rect 7236 34894 7292 34950
rect 7360 34894 7416 34950
rect 6368 34770 6424 34826
rect 6492 34770 6548 34826
rect 6616 34770 6672 34826
rect 6740 34770 6796 34826
rect 6864 34770 6920 34826
rect 6988 34770 7044 34826
rect 7112 34770 7168 34826
rect 7236 34770 7292 34826
rect 7360 34770 7416 34826
rect 6368 34646 6424 34702
rect 6492 34646 6548 34702
rect 6616 34646 6672 34702
rect 6740 34646 6796 34702
rect 6864 34646 6920 34702
rect 6988 34646 7044 34702
rect 7112 34646 7168 34702
rect 7236 34646 7292 34702
rect 7360 34646 7416 34702
rect 6368 34522 6424 34578
rect 6492 34522 6548 34578
rect 6616 34522 6672 34578
rect 6740 34522 6796 34578
rect 6864 34522 6920 34578
rect 6988 34522 7044 34578
rect 7112 34522 7168 34578
rect 7236 34522 7292 34578
rect 7360 34522 7416 34578
rect 6368 34398 6424 34454
rect 6492 34398 6548 34454
rect 6616 34398 6672 34454
rect 6740 34398 6796 34454
rect 6864 34398 6920 34454
rect 6988 34398 7044 34454
rect 7112 34398 7168 34454
rect 7236 34398 7292 34454
rect 7360 34398 7416 34454
rect 6368 34274 6424 34330
rect 6492 34274 6548 34330
rect 6616 34274 6672 34330
rect 6740 34274 6796 34330
rect 6864 34274 6920 34330
rect 6988 34274 7044 34330
rect 7112 34274 7168 34330
rect 7236 34274 7292 34330
rect 7360 34274 7416 34330
rect 6368 34150 6424 34206
rect 6492 34150 6548 34206
rect 6616 34150 6672 34206
rect 6740 34150 6796 34206
rect 6864 34150 6920 34206
rect 6988 34150 7044 34206
rect 7112 34150 7168 34206
rect 7236 34150 7292 34206
rect 7360 34150 7416 34206
rect 6368 34026 6424 34082
rect 6492 34026 6548 34082
rect 6616 34026 6672 34082
rect 6740 34026 6796 34082
rect 6864 34026 6920 34082
rect 6988 34026 7044 34082
rect 7112 34026 7168 34082
rect 7236 34026 7292 34082
rect 7360 34026 7416 34082
rect 6368 33902 6424 33958
rect 6492 33902 6548 33958
rect 6616 33902 6672 33958
rect 6740 33902 6796 33958
rect 6864 33902 6920 33958
rect 6988 33902 7044 33958
rect 7112 33902 7168 33958
rect 7236 33902 7292 33958
rect 7360 33902 7416 33958
rect 6368 33778 6424 33834
rect 6492 33778 6548 33834
rect 6616 33778 6672 33834
rect 6740 33778 6796 33834
rect 6864 33778 6920 33834
rect 6988 33778 7044 33834
rect 7112 33778 7168 33834
rect 7236 33778 7292 33834
rect 7360 33778 7416 33834
rect 6368 33654 6424 33710
rect 6492 33654 6548 33710
rect 6616 33654 6672 33710
rect 6740 33654 6796 33710
rect 6864 33654 6920 33710
rect 6988 33654 7044 33710
rect 7112 33654 7168 33710
rect 7236 33654 7292 33710
rect 7360 33654 7416 33710
rect 6368 33530 6424 33586
rect 6492 33530 6548 33586
rect 6616 33530 6672 33586
rect 6740 33530 6796 33586
rect 6864 33530 6920 33586
rect 6988 33530 7044 33586
rect 7112 33530 7168 33586
rect 7236 33530 7292 33586
rect 7360 33530 7416 33586
rect 6368 33406 6424 33462
rect 6492 33406 6548 33462
rect 6616 33406 6672 33462
rect 6740 33406 6796 33462
rect 6864 33406 6920 33462
rect 6988 33406 7044 33462
rect 7112 33406 7168 33462
rect 7236 33406 7292 33462
rect 7360 33406 7416 33462
rect 6368 33282 6424 33338
rect 6492 33282 6548 33338
rect 6616 33282 6672 33338
rect 6740 33282 6796 33338
rect 6864 33282 6920 33338
rect 6988 33282 7044 33338
rect 7112 33282 7168 33338
rect 7236 33282 7292 33338
rect 7360 33282 7416 33338
rect 6368 33158 6424 33214
rect 6492 33158 6548 33214
rect 6616 33158 6672 33214
rect 6740 33158 6796 33214
rect 6864 33158 6920 33214
rect 6988 33158 7044 33214
rect 7112 33158 7168 33214
rect 7236 33158 7292 33214
rect 7360 33158 7416 33214
rect 6368 33034 6424 33090
rect 6492 33034 6548 33090
rect 6616 33034 6672 33090
rect 6740 33034 6796 33090
rect 6864 33034 6920 33090
rect 6988 33034 7044 33090
rect 7112 33034 7168 33090
rect 7236 33034 7292 33090
rect 7360 33034 7416 33090
rect 6368 32910 6424 32966
rect 6492 32910 6548 32966
rect 6616 32910 6672 32966
rect 6740 32910 6796 32966
rect 6864 32910 6920 32966
rect 6988 32910 7044 32966
rect 7112 32910 7168 32966
rect 7236 32910 7292 32966
rect 7360 32910 7416 32966
rect 6368 32786 6424 32842
rect 6492 32786 6548 32842
rect 6616 32786 6672 32842
rect 6740 32786 6796 32842
rect 6864 32786 6920 32842
rect 6988 32786 7044 32842
rect 7112 32786 7168 32842
rect 7236 32786 7292 32842
rect 7360 32786 7416 32842
rect 6368 32662 6424 32718
rect 6492 32662 6548 32718
rect 6616 32662 6672 32718
rect 6740 32662 6796 32718
rect 6864 32662 6920 32718
rect 6988 32662 7044 32718
rect 7112 32662 7168 32718
rect 7236 32662 7292 32718
rect 7360 32662 7416 32718
rect 6368 32538 6424 32594
rect 6492 32538 6548 32594
rect 6616 32538 6672 32594
rect 6740 32538 6796 32594
rect 6864 32538 6920 32594
rect 6988 32538 7044 32594
rect 7112 32538 7168 32594
rect 7236 32538 7292 32594
rect 7360 32538 7416 32594
rect 6368 32414 6424 32470
rect 6492 32414 6548 32470
rect 6616 32414 6672 32470
rect 6740 32414 6796 32470
rect 6864 32414 6920 32470
rect 6988 32414 7044 32470
rect 7112 32414 7168 32470
rect 7236 32414 7292 32470
rect 7360 32414 7416 32470
rect 6368 32290 6424 32346
rect 6492 32290 6548 32346
rect 6616 32290 6672 32346
rect 6740 32290 6796 32346
rect 6864 32290 6920 32346
rect 6988 32290 7044 32346
rect 7112 32290 7168 32346
rect 7236 32290 7292 32346
rect 7360 32290 7416 32346
rect 6368 32166 6424 32222
rect 6492 32166 6548 32222
rect 6616 32166 6672 32222
rect 6740 32166 6796 32222
rect 6864 32166 6920 32222
rect 6988 32166 7044 32222
rect 7112 32166 7168 32222
rect 7236 32166 7292 32222
rect 7360 32166 7416 32222
rect 6368 32042 6424 32098
rect 6492 32042 6548 32098
rect 6616 32042 6672 32098
rect 6740 32042 6796 32098
rect 6864 32042 6920 32098
rect 6988 32042 7044 32098
rect 7112 32042 7168 32098
rect 7236 32042 7292 32098
rect 7360 32042 7416 32098
rect 8751 34894 8807 34950
rect 8875 34894 8931 34950
rect 8999 34894 9055 34950
rect 9123 34894 9179 34950
rect 9247 34894 9303 34950
rect 9371 34894 9427 34950
rect 9495 34894 9551 34950
rect 9619 34894 9675 34950
rect 9743 34894 9799 34950
rect 9867 34894 9923 34950
rect 9991 34894 10047 34950
rect 10115 34894 10171 34950
rect 10239 34894 10295 34950
rect 10363 34894 10419 34950
rect 10487 34894 10543 34950
rect 8751 34770 8807 34826
rect 8875 34770 8931 34826
rect 8999 34770 9055 34826
rect 9123 34770 9179 34826
rect 9247 34770 9303 34826
rect 9371 34770 9427 34826
rect 9495 34770 9551 34826
rect 9619 34770 9675 34826
rect 9743 34770 9799 34826
rect 9867 34770 9923 34826
rect 9991 34770 10047 34826
rect 10115 34770 10171 34826
rect 10239 34770 10295 34826
rect 10363 34770 10419 34826
rect 10487 34770 10543 34826
rect 8751 34646 8807 34702
rect 8875 34646 8931 34702
rect 8999 34646 9055 34702
rect 9123 34646 9179 34702
rect 9247 34646 9303 34702
rect 9371 34646 9427 34702
rect 9495 34646 9551 34702
rect 9619 34646 9675 34702
rect 9743 34646 9799 34702
rect 9867 34646 9923 34702
rect 9991 34646 10047 34702
rect 10115 34646 10171 34702
rect 10239 34646 10295 34702
rect 10363 34646 10419 34702
rect 10487 34646 10543 34702
rect 8751 34522 8807 34578
rect 8875 34522 8931 34578
rect 8999 34522 9055 34578
rect 9123 34522 9179 34578
rect 9247 34522 9303 34578
rect 9371 34522 9427 34578
rect 9495 34522 9551 34578
rect 9619 34522 9675 34578
rect 9743 34522 9799 34578
rect 9867 34522 9923 34578
rect 9991 34522 10047 34578
rect 10115 34522 10171 34578
rect 10239 34522 10295 34578
rect 10363 34522 10419 34578
rect 10487 34522 10543 34578
rect 8751 34398 8807 34454
rect 8875 34398 8931 34454
rect 8999 34398 9055 34454
rect 9123 34398 9179 34454
rect 9247 34398 9303 34454
rect 9371 34398 9427 34454
rect 9495 34398 9551 34454
rect 9619 34398 9675 34454
rect 9743 34398 9799 34454
rect 9867 34398 9923 34454
rect 9991 34398 10047 34454
rect 10115 34398 10171 34454
rect 10239 34398 10295 34454
rect 10363 34398 10419 34454
rect 10487 34398 10543 34454
rect 8751 34274 8807 34330
rect 8875 34274 8931 34330
rect 8999 34274 9055 34330
rect 9123 34274 9179 34330
rect 9247 34274 9303 34330
rect 9371 34274 9427 34330
rect 9495 34274 9551 34330
rect 9619 34274 9675 34330
rect 9743 34274 9799 34330
rect 9867 34274 9923 34330
rect 9991 34274 10047 34330
rect 10115 34274 10171 34330
rect 10239 34274 10295 34330
rect 10363 34274 10419 34330
rect 10487 34274 10543 34330
rect 8751 34150 8807 34206
rect 8875 34150 8931 34206
rect 8999 34150 9055 34206
rect 9123 34150 9179 34206
rect 9247 34150 9303 34206
rect 9371 34150 9427 34206
rect 9495 34150 9551 34206
rect 9619 34150 9675 34206
rect 9743 34150 9799 34206
rect 9867 34150 9923 34206
rect 9991 34150 10047 34206
rect 10115 34150 10171 34206
rect 10239 34150 10295 34206
rect 10363 34150 10419 34206
rect 10487 34150 10543 34206
rect 8751 34026 8807 34082
rect 8875 34026 8931 34082
rect 8999 34026 9055 34082
rect 9123 34026 9179 34082
rect 9247 34026 9303 34082
rect 9371 34026 9427 34082
rect 9495 34026 9551 34082
rect 9619 34026 9675 34082
rect 9743 34026 9799 34082
rect 9867 34026 9923 34082
rect 9991 34026 10047 34082
rect 10115 34026 10171 34082
rect 10239 34026 10295 34082
rect 10363 34026 10419 34082
rect 10487 34026 10543 34082
rect 8751 33902 8807 33958
rect 8875 33902 8931 33958
rect 8999 33902 9055 33958
rect 9123 33902 9179 33958
rect 9247 33902 9303 33958
rect 9371 33902 9427 33958
rect 9495 33902 9551 33958
rect 9619 33902 9675 33958
rect 9743 33902 9799 33958
rect 9867 33902 9923 33958
rect 9991 33902 10047 33958
rect 10115 33902 10171 33958
rect 10239 33902 10295 33958
rect 10363 33902 10419 33958
rect 10487 33902 10543 33958
rect 8751 33778 8807 33834
rect 8875 33778 8931 33834
rect 8999 33778 9055 33834
rect 9123 33778 9179 33834
rect 9247 33778 9303 33834
rect 9371 33778 9427 33834
rect 9495 33778 9551 33834
rect 9619 33778 9675 33834
rect 9743 33778 9799 33834
rect 9867 33778 9923 33834
rect 9991 33778 10047 33834
rect 10115 33778 10171 33834
rect 10239 33778 10295 33834
rect 10363 33778 10419 33834
rect 10487 33778 10543 33834
rect 8751 33654 8807 33710
rect 8875 33654 8931 33710
rect 8999 33654 9055 33710
rect 9123 33654 9179 33710
rect 9247 33654 9303 33710
rect 9371 33654 9427 33710
rect 9495 33654 9551 33710
rect 9619 33654 9675 33710
rect 9743 33654 9799 33710
rect 9867 33654 9923 33710
rect 9991 33654 10047 33710
rect 10115 33654 10171 33710
rect 10239 33654 10295 33710
rect 10363 33654 10419 33710
rect 10487 33654 10543 33710
rect 8751 33530 8807 33586
rect 8875 33530 8931 33586
rect 8999 33530 9055 33586
rect 9123 33530 9179 33586
rect 9247 33530 9303 33586
rect 9371 33530 9427 33586
rect 9495 33530 9551 33586
rect 9619 33530 9675 33586
rect 9743 33530 9799 33586
rect 9867 33530 9923 33586
rect 9991 33530 10047 33586
rect 10115 33530 10171 33586
rect 10239 33530 10295 33586
rect 10363 33530 10419 33586
rect 10487 33530 10543 33586
rect 8751 33406 8807 33462
rect 8875 33406 8931 33462
rect 8999 33406 9055 33462
rect 9123 33406 9179 33462
rect 9247 33406 9303 33462
rect 9371 33406 9427 33462
rect 9495 33406 9551 33462
rect 9619 33406 9675 33462
rect 9743 33406 9799 33462
rect 9867 33406 9923 33462
rect 9991 33406 10047 33462
rect 10115 33406 10171 33462
rect 10239 33406 10295 33462
rect 10363 33406 10419 33462
rect 10487 33406 10543 33462
rect 8751 33282 8807 33338
rect 8875 33282 8931 33338
rect 8999 33282 9055 33338
rect 9123 33282 9179 33338
rect 9247 33282 9303 33338
rect 9371 33282 9427 33338
rect 9495 33282 9551 33338
rect 9619 33282 9675 33338
rect 9743 33282 9799 33338
rect 9867 33282 9923 33338
rect 9991 33282 10047 33338
rect 10115 33282 10171 33338
rect 10239 33282 10295 33338
rect 10363 33282 10419 33338
rect 10487 33282 10543 33338
rect 8751 33158 8807 33214
rect 8875 33158 8931 33214
rect 8999 33158 9055 33214
rect 9123 33158 9179 33214
rect 9247 33158 9303 33214
rect 9371 33158 9427 33214
rect 9495 33158 9551 33214
rect 9619 33158 9675 33214
rect 9743 33158 9799 33214
rect 9867 33158 9923 33214
rect 9991 33158 10047 33214
rect 10115 33158 10171 33214
rect 10239 33158 10295 33214
rect 10363 33158 10419 33214
rect 10487 33158 10543 33214
rect 8751 33034 8807 33090
rect 8875 33034 8931 33090
rect 8999 33034 9055 33090
rect 9123 33034 9179 33090
rect 9247 33034 9303 33090
rect 9371 33034 9427 33090
rect 9495 33034 9551 33090
rect 9619 33034 9675 33090
rect 9743 33034 9799 33090
rect 9867 33034 9923 33090
rect 9991 33034 10047 33090
rect 10115 33034 10171 33090
rect 10239 33034 10295 33090
rect 10363 33034 10419 33090
rect 10487 33034 10543 33090
rect 8751 32910 8807 32966
rect 8875 32910 8931 32966
rect 8999 32910 9055 32966
rect 9123 32910 9179 32966
rect 9247 32910 9303 32966
rect 9371 32910 9427 32966
rect 9495 32910 9551 32966
rect 9619 32910 9675 32966
rect 9743 32910 9799 32966
rect 9867 32910 9923 32966
rect 9991 32910 10047 32966
rect 10115 32910 10171 32966
rect 10239 32910 10295 32966
rect 10363 32910 10419 32966
rect 10487 32910 10543 32966
rect 8751 32786 8807 32842
rect 8875 32786 8931 32842
rect 8999 32786 9055 32842
rect 9123 32786 9179 32842
rect 9247 32786 9303 32842
rect 9371 32786 9427 32842
rect 9495 32786 9551 32842
rect 9619 32786 9675 32842
rect 9743 32786 9799 32842
rect 9867 32786 9923 32842
rect 9991 32786 10047 32842
rect 10115 32786 10171 32842
rect 10239 32786 10295 32842
rect 10363 32786 10419 32842
rect 10487 32786 10543 32842
rect 8751 32662 8807 32718
rect 8875 32662 8931 32718
rect 8999 32662 9055 32718
rect 9123 32662 9179 32718
rect 9247 32662 9303 32718
rect 9371 32662 9427 32718
rect 9495 32662 9551 32718
rect 9619 32662 9675 32718
rect 9743 32662 9799 32718
rect 9867 32662 9923 32718
rect 9991 32662 10047 32718
rect 10115 32662 10171 32718
rect 10239 32662 10295 32718
rect 10363 32662 10419 32718
rect 10487 32662 10543 32718
rect 8751 32538 8807 32594
rect 8875 32538 8931 32594
rect 8999 32538 9055 32594
rect 9123 32538 9179 32594
rect 9247 32538 9303 32594
rect 9371 32538 9427 32594
rect 9495 32538 9551 32594
rect 9619 32538 9675 32594
rect 9743 32538 9799 32594
rect 9867 32538 9923 32594
rect 9991 32538 10047 32594
rect 10115 32538 10171 32594
rect 10239 32538 10295 32594
rect 10363 32538 10419 32594
rect 10487 32538 10543 32594
rect 8751 32414 8807 32470
rect 8875 32414 8931 32470
rect 8999 32414 9055 32470
rect 9123 32414 9179 32470
rect 9247 32414 9303 32470
rect 9371 32414 9427 32470
rect 9495 32414 9551 32470
rect 9619 32414 9675 32470
rect 9743 32414 9799 32470
rect 9867 32414 9923 32470
rect 9991 32414 10047 32470
rect 10115 32414 10171 32470
rect 10239 32414 10295 32470
rect 10363 32414 10419 32470
rect 10487 32414 10543 32470
rect 8751 32290 8807 32346
rect 8875 32290 8931 32346
rect 8999 32290 9055 32346
rect 9123 32290 9179 32346
rect 9247 32290 9303 32346
rect 9371 32290 9427 32346
rect 9495 32290 9551 32346
rect 9619 32290 9675 32346
rect 9743 32290 9799 32346
rect 9867 32290 9923 32346
rect 9991 32290 10047 32346
rect 10115 32290 10171 32346
rect 10239 32290 10295 32346
rect 10363 32290 10419 32346
rect 10487 32290 10543 32346
rect 8751 32166 8807 32222
rect 8875 32166 8931 32222
rect 8999 32166 9055 32222
rect 9123 32166 9179 32222
rect 9247 32166 9303 32222
rect 9371 32166 9427 32222
rect 9495 32166 9551 32222
rect 9619 32166 9675 32222
rect 9743 32166 9799 32222
rect 9867 32166 9923 32222
rect 9991 32166 10047 32222
rect 10115 32166 10171 32222
rect 10239 32166 10295 32222
rect 10363 32166 10419 32222
rect 10487 32166 10543 32222
rect 8751 32042 8807 32098
rect 8875 32042 8931 32098
rect 8999 32042 9055 32098
rect 9123 32042 9179 32098
rect 9247 32042 9303 32098
rect 9371 32042 9427 32098
rect 9495 32042 9551 32098
rect 9619 32042 9675 32098
rect 9743 32042 9799 32098
rect 9867 32042 9923 32098
rect 9991 32042 10047 32098
rect 10115 32042 10171 32098
rect 10239 32042 10295 32098
rect 10363 32042 10419 32098
rect 10487 32042 10543 32098
rect 12852 34894 12908 34950
rect 12976 34894 13032 34950
rect 13100 34894 13156 34950
rect 13224 34894 13280 34950
rect 13348 34894 13404 34950
rect 13472 34894 13528 34950
rect 13596 34894 13652 34950
rect 13720 34894 13776 34950
rect 13844 34894 13900 34950
rect 12852 34770 12908 34826
rect 12976 34770 13032 34826
rect 13100 34770 13156 34826
rect 13224 34770 13280 34826
rect 13348 34770 13404 34826
rect 13472 34770 13528 34826
rect 13596 34770 13652 34826
rect 13720 34770 13776 34826
rect 13844 34770 13900 34826
rect 12852 34646 12908 34702
rect 12976 34646 13032 34702
rect 13100 34646 13156 34702
rect 13224 34646 13280 34702
rect 13348 34646 13404 34702
rect 13472 34646 13528 34702
rect 13596 34646 13652 34702
rect 13720 34646 13776 34702
rect 13844 34646 13900 34702
rect 12852 34522 12908 34578
rect 12976 34522 13032 34578
rect 13100 34522 13156 34578
rect 13224 34522 13280 34578
rect 13348 34522 13404 34578
rect 13472 34522 13528 34578
rect 13596 34522 13652 34578
rect 13720 34522 13776 34578
rect 13844 34522 13900 34578
rect 12852 34398 12908 34454
rect 12976 34398 13032 34454
rect 13100 34398 13156 34454
rect 13224 34398 13280 34454
rect 13348 34398 13404 34454
rect 13472 34398 13528 34454
rect 13596 34398 13652 34454
rect 13720 34398 13776 34454
rect 13844 34398 13900 34454
rect 12852 34274 12908 34330
rect 12976 34274 13032 34330
rect 13100 34274 13156 34330
rect 13224 34274 13280 34330
rect 13348 34274 13404 34330
rect 13472 34274 13528 34330
rect 13596 34274 13652 34330
rect 13720 34274 13776 34330
rect 13844 34274 13900 34330
rect 12852 34150 12908 34206
rect 12976 34150 13032 34206
rect 13100 34150 13156 34206
rect 13224 34150 13280 34206
rect 13348 34150 13404 34206
rect 13472 34150 13528 34206
rect 13596 34150 13652 34206
rect 13720 34150 13776 34206
rect 13844 34150 13900 34206
rect 12852 34026 12908 34082
rect 12976 34026 13032 34082
rect 13100 34026 13156 34082
rect 13224 34026 13280 34082
rect 13348 34026 13404 34082
rect 13472 34026 13528 34082
rect 13596 34026 13652 34082
rect 13720 34026 13776 34082
rect 13844 34026 13900 34082
rect 12852 33902 12908 33958
rect 12976 33902 13032 33958
rect 13100 33902 13156 33958
rect 13224 33902 13280 33958
rect 13348 33902 13404 33958
rect 13472 33902 13528 33958
rect 13596 33902 13652 33958
rect 13720 33902 13776 33958
rect 13844 33902 13900 33958
rect 12852 33778 12908 33834
rect 12976 33778 13032 33834
rect 13100 33778 13156 33834
rect 13224 33778 13280 33834
rect 13348 33778 13404 33834
rect 13472 33778 13528 33834
rect 13596 33778 13652 33834
rect 13720 33778 13776 33834
rect 13844 33778 13900 33834
rect 12852 33654 12908 33710
rect 12976 33654 13032 33710
rect 13100 33654 13156 33710
rect 13224 33654 13280 33710
rect 13348 33654 13404 33710
rect 13472 33654 13528 33710
rect 13596 33654 13652 33710
rect 13720 33654 13776 33710
rect 13844 33654 13900 33710
rect 12852 33530 12908 33586
rect 12976 33530 13032 33586
rect 13100 33530 13156 33586
rect 13224 33530 13280 33586
rect 13348 33530 13404 33586
rect 13472 33530 13528 33586
rect 13596 33530 13652 33586
rect 13720 33530 13776 33586
rect 13844 33530 13900 33586
rect 12852 33406 12908 33462
rect 12976 33406 13032 33462
rect 13100 33406 13156 33462
rect 13224 33406 13280 33462
rect 13348 33406 13404 33462
rect 13472 33406 13528 33462
rect 13596 33406 13652 33462
rect 13720 33406 13776 33462
rect 13844 33406 13900 33462
rect 12852 33282 12908 33338
rect 12976 33282 13032 33338
rect 13100 33282 13156 33338
rect 13224 33282 13280 33338
rect 13348 33282 13404 33338
rect 13472 33282 13528 33338
rect 13596 33282 13652 33338
rect 13720 33282 13776 33338
rect 13844 33282 13900 33338
rect 12852 33158 12908 33214
rect 12976 33158 13032 33214
rect 13100 33158 13156 33214
rect 13224 33158 13280 33214
rect 13348 33158 13404 33214
rect 13472 33158 13528 33214
rect 13596 33158 13652 33214
rect 13720 33158 13776 33214
rect 13844 33158 13900 33214
rect 12852 33034 12908 33090
rect 12976 33034 13032 33090
rect 13100 33034 13156 33090
rect 13224 33034 13280 33090
rect 13348 33034 13404 33090
rect 13472 33034 13528 33090
rect 13596 33034 13652 33090
rect 13720 33034 13776 33090
rect 13844 33034 13900 33090
rect 12852 32910 12908 32966
rect 12976 32910 13032 32966
rect 13100 32910 13156 32966
rect 13224 32910 13280 32966
rect 13348 32910 13404 32966
rect 13472 32910 13528 32966
rect 13596 32910 13652 32966
rect 13720 32910 13776 32966
rect 13844 32910 13900 32966
rect 12852 32786 12908 32842
rect 12976 32786 13032 32842
rect 13100 32786 13156 32842
rect 13224 32786 13280 32842
rect 13348 32786 13404 32842
rect 13472 32786 13528 32842
rect 13596 32786 13652 32842
rect 13720 32786 13776 32842
rect 13844 32786 13900 32842
rect 12852 32662 12908 32718
rect 12976 32662 13032 32718
rect 13100 32662 13156 32718
rect 13224 32662 13280 32718
rect 13348 32662 13404 32718
rect 13472 32662 13528 32718
rect 13596 32662 13652 32718
rect 13720 32662 13776 32718
rect 13844 32662 13900 32718
rect 12852 32538 12908 32594
rect 12976 32538 13032 32594
rect 13100 32538 13156 32594
rect 13224 32538 13280 32594
rect 13348 32538 13404 32594
rect 13472 32538 13528 32594
rect 13596 32538 13652 32594
rect 13720 32538 13776 32594
rect 13844 32538 13900 32594
rect 12852 32414 12908 32470
rect 12976 32414 13032 32470
rect 13100 32414 13156 32470
rect 13224 32414 13280 32470
rect 13348 32414 13404 32470
rect 13472 32414 13528 32470
rect 13596 32414 13652 32470
rect 13720 32414 13776 32470
rect 13844 32414 13900 32470
rect 12852 32290 12908 32346
rect 12976 32290 13032 32346
rect 13100 32290 13156 32346
rect 13224 32290 13280 32346
rect 13348 32290 13404 32346
rect 13472 32290 13528 32346
rect 13596 32290 13652 32346
rect 13720 32290 13776 32346
rect 13844 32290 13900 32346
rect 12852 32166 12908 32222
rect 12976 32166 13032 32222
rect 13100 32166 13156 32222
rect 13224 32166 13280 32222
rect 13348 32166 13404 32222
rect 13472 32166 13528 32222
rect 13596 32166 13652 32222
rect 13720 32166 13776 32222
rect 13844 32166 13900 32222
rect 12852 32042 12908 32098
rect 12976 32042 13032 32098
rect 13100 32042 13156 32098
rect 13224 32042 13280 32098
rect 13348 32042 13404 32098
rect 13472 32042 13528 32098
rect 13596 32042 13652 32098
rect 13720 32042 13776 32098
rect 13844 32042 13900 32098
rect 2023 31850 2079 31906
rect 2023 31726 2079 31782
rect 2023 31602 2079 31658
rect 2023 31478 2079 31534
rect 2023 31354 2079 31410
rect 2023 31230 2079 31286
rect 2023 31106 2079 31162
rect 2023 30982 2079 31038
rect 2023 30858 2079 30914
rect 2023 30734 2079 30790
rect 2023 30610 2079 30666
rect 2023 30486 2079 30542
rect 2023 30362 2079 30418
rect 2023 30238 2079 30294
rect 2023 30114 2079 30170
rect 2023 29990 2079 30046
rect 2023 29866 2079 29922
rect 2023 29742 2079 29798
rect 2023 29618 2079 29674
rect 2023 29494 2079 29550
rect 2023 29370 2079 29426
rect 2023 29246 2079 29302
rect 2023 29122 2079 29178
rect 2023 28998 2079 29054
rect 1375 28879 1431 28935
rect 1375 28755 1431 28811
rect 1375 28631 1431 28687
rect 1375 28507 1431 28563
rect 1375 28383 1431 28439
rect 1375 28259 1431 28315
rect 1375 28135 1431 28191
rect 1375 28011 1431 28067
rect 1375 27887 1431 27943
rect 1375 27763 1431 27819
rect 1375 27639 1431 27695
rect 1375 27515 1431 27571
rect 1375 27391 1431 27447
rect 1375 27267 1431 27323
rect 1499 28866 1555 28922
rect 2023 28874 2079 28930
rect 4435 31694 4491 31750
rect 4559 31694 4615 31750
rect 4683 31694 4739 31750
rect 4807 31694 4863 31750
rect 4931 31694 4987 31750
rect 5055 31694 5111 31750
rect 5179 31694 5235 31750
rect 5303 31694 5359 31750
rect 5427 31694 5483 31750
rect 5551 31694 5607 31750
rect 5675 31694 5731 31750
rect 5799 31694 5855 31750
rect 5923 31694 5979 31750
rect 6047 31694 6103 31750
rect 6171 31694 6227 31750
rect 4435 31570 4491 31626
rect 4559 31570 4615 31626
rect 4683 31570 4739 31626
rect 4807 31570 4863 31626
rect 4931 31570 4987 31626
rect 5055 31570 5111 31626
rect 5179 31570 5235 31626
rect 5303 31570 5359 31626
rect 5427 31570 5483 31626
rect 5551 31570 5607 31626
rect 5675 31570 5731 31626
rect 5799 31570 5855 31626
rect 5923 31570 5979 31626
rect 6047 31570 6103 31626
rect 6171 31570 6227 31626
rect 4435 31446 4491 31502
rect 4559 31446 4615 31502
rect 4683 31446 4739 31502
rect 4807 31446 4863 31502
rect 4931 31446 4987 31502
rect 5055 31446 5111 31502
rect 5179 31446 5235 31502
rect 5303 31446 5359 31502
rect 5427 31446 5483 31502
rect 5551 31446 5607 31502
rect 5675 31446 5731 31502
rect 5799 31446 5855 31502
rect 5923 31446 5979 31502
rect 6047 31446 6103 31502
rect 6171 31446 6227 31502
rect 4435 31322 4491 31378
rect 4559 31322 4615 31378
rect 4683 31322 4739 31378
rect 4807 31322 4863 31378
rect 4931 31322 4987 31378
rect 5055 31322 5111 31378
rect 5179 31322 5235 31378
rect 5303 31322 5359 31378
rect 5427 31322 5483 31378
rect 5551 31322 5607 31378
rect 5675 31322 5731 31378
rect 5799 31322 5855 31378
rect 5923 31322 5979 31378
rect 6047 31322 6103 31378
rect 6171 31322 6227 31378
rect 4435 31198 4491 31254
rect 4559 31198 4615 31254
rect 4683 31198 4739 31254
rect 4807 31198 4863 31254
rect 4931 31198 4987 31254
rect 5055 31198 5111 31254
rect 5179 31198 5235 31254
rect 5303 31198 5359 31254
rect 5427 31198 5483 31254
rect 5551 31198 5607 31254
rect 5675 31198 5731 31254
rect 5799 31198 5855 31254
rect 5923 31198 5979 31254
rect 6047 31198 6103 31254
rect 6171 31198 6227 31254
rect 4435 31074 4491 31130
rect 4559 31074 4615 31130
rect 4683 31074 4739 31130
rect 4807 31074 4863 31130
rect 4931 31074 4987 31130
rect 5055 31074 5111 31130
rect 5179 31074 5235 31130
rect 5303 31074 5359 31130
rect 5427 31074 5483 31130
rect 5551 31074 5607 31130
rect 5675 31074 5731 31130
rect 5799 31074 5855 31130
rect 5923 31074 5979 31130
rect 6047 31074 6103 31130
rect 6171 31074 6227 31130
rect 4435 30950 4491 31006
rect 4559 30950 4615 31006
rect 4683 30950 4739 31006
rect 4807 30950 4863 31006
rect 4931 30950 4987 31006
rect 5055 30950 5111 31006
rect 5179 30950 5235 31006
rect 5303 30950 5359 31006
rect 5427 30950 5483 31006
rect 5551 30950 5607 31006
rect 5675 30950 5731 31006
rect 5799 30950 5855 31006
rect 5923 30950 5979 31006
rect 6047 30950 6103 31006
rect 6171 30950 6227 31006
rect 4435 30826 4491 30882
rect 4559 30826 4615 30882
rect 4683 30826 4739 30882
rect 4807 30826 4863 30882
rect 4931 30826 4987 30882
rect 5055 30826 5111 30882
rect 5179 30826 5235 30882
rect 5303 30826 5359 30882
rect 5427 30826 5483 30882
rect 5551 30826 5607 30882
rect 5675 30826 5731 30882
rect 5799 30826 5855 30882
rect 5923 30826 5979 30882
rect 6047 30826 6103 30882
rect 6171 30826 6227 30882
rect 4435 30702 4491 30758
rect 4559 30702 4615 30758
rect 4683 30702 4739 30758
rect 4807 30702 4863 30758
rect 4931 30702 4987 30758
rect 5055 30702 5111 30758
rect 5179 30702 5235 30758
rect 5303 30702 5359 30758
rect 5427 30702 5483 30758
rect 5551 30702 5607 30758
rect 5675 30702 5731 30758
rect 5799 30702 5855 30758
rect 5923 30702 5979 30758
rect 6047 30702 6103 30758
rect 6171 30702 6227 30758
rect 4435 30578 4491 30634
rect 4559 30578 4615 30634
rect 4683 30578 4739 30634
rect 4807 30578 4863 30634
rect 4931 30578 4987 30634
rect 5055 30578 5111 30634
rect 5179 30578 5235 30634
rect 5303 30578 5359 30634
rect 5427 30578 5483 30634
rect 5551 30578 5607 30634
rect 5675 30578 5731 30634
rect 5799 30578 5855 30634
rect 5923 30578 5979 30634
rect 6047 30578 6103 30634
rect 6171 30578 6227 30634
rect 4435 30454 4491 30510
rect 4559 30454 4615 30510
rect 4683 30454 4739 30510
rect 4807 30454 4863 30510
rect 4931 30454 4987 30510
rect 5055 30454 5111 30510
rect 5179 30454 5235 30510
rect 5303 30454 5359 30510
rect 5427 30454 5483 30510
rect 5551 30454 5607 30510
rect 5675 30454 5731 30510
rect 5799 30454 5855 30510
rect 5923 30454 5979 30510
rect 6047 30454 6103 30510
rect 6171 30454 6227 30510
rect 4435 30330 4491 30386
rect 4559 30330 4615 30386
rect 4683 30330 4739 30386
rect 4807 30330 4863 30386
rect 4931 30330 4987 30386
rect 5055 30330 5111 30386
rect 5179 30330 5235 30386
rect 5303 30330 5359 30386
rect 5427 30330 5483 30386
rect 5551 30330 5607 30386
rect 5675 30330 5731 30386
rect 5799 30330 5855 30386
rect 5923 30330 5979 30386
rect 6047 30330 6103 30386
rect 6171 30330 6227 30386
rect 4435 30206 4491 30262
rect 4559 30206 4615 30262
rect 4683 30206 4739 30262
rect 4807 30206 4863 30262
rect 4931 30206 4987 30262
rect 5055 30206 5111 30262
rect 5179 30206 5235 30262
rect 5303 30206 5359 30262
rect 5427 30206 5483 30262
rect 5551 30206 5607 30262
rect 5675 30206 5731 30262
rect 5799 30206 5855 30262
rect 5923 30206 5979 30262
rect 6047 30206 6103 30262
rect 6171 30206 6227 30262
rect 4435 30082 4491 30138
rect 4559 30082 4615 30138
rect 4683 30082 4739 30138
rect 4807 30082 4863 30138
rect 4931 30082 4987 30138
rect 5055 30082 5111 30138
rect 5179 30082 5235 30138
rect 5303 30082 5359 30138
rect 5427 30082 5483 30138
rect 5551 30082 5607 30138
rect 5675 30082 5731 30138
rect 5799 30082 5855 30138
rect 5923 30082 5979 30138
rect 6047 30082 6103 30138
rect 6171 30082 6227 30138
rect 4435 29958 4491 30014
rect 4559 29958 4615 30014
rect 4683 29958 4739 30014
rect 4807 29958 4863 30014
rect 4931 29958 4987 30014
rect 5055 29958 5111 30014
rect 5179 29958 5235 30014
rect 5303 29958 5359 30014
rect 5427 29958 5483 30014
rect 5551 29958 5607 30014
rect 5675 29958 5731 30014
rect 5799 29958 5855 30014
rect 5923 29958 5979 30014
rect 6047 29958 6103 30014
rect 6171 29958 6227 30014
rect 4435 29834 4491 29890
rect 4559 29834 4615 29890
rect 4683 29834 4739 29890
rect 4807 29834 4863 29890
rect 4931 29834 4987 29890
rect 5055 29834 5111 29890
rect 5179 29834 5235 29890
rect 5303 29834 5359 29890
rect 5427 29834 5483 29890
rect 5551 29834 5607 29890
rect 5675 29834 5731 29890
rect 5799 29834 5855 29890
rect 5923 29834 5979 29890
rect 6047 29834 6103 29890
rect 6171 29834 6227 29890
rect 4435 29710 4491 29766
rect 4559 29710 4615 29766
rect 4683 29710 4739 29766
rect 4807 29710 4863 29766
rect 4931 29710 4987 29766
rect 5055 29710 5111 29766
rect 5179 29710 5235 29766
rect 5303 29710 5359 29766
rect 5427 29710 5483 29766
rect 5551 29710 5607 29766
rect 5675 29710 5731 29766
rect 5799 29710 5855 29766
rect 5923 29710 5979 29766
rect 6047 29710 6103 29766
rect 6171 29710 6227 29766
rect 4435 29586 4491 29642
rect 4559 29586 4615 29642
rect 4683 29586 4739 29642
rect 4807 29586 4863 29642
rect 4931 29586 4987 29642
rect 5055 29586 5111 29642
rect 5179 29586 5235 29642
rect 5303 29586 5359 29642
rect 5427 29586 5483 29642
rect 5551 29586 5607 29642
rect 5675 29586 5731 29642
rect 5799 29586 5855 29642
rect 5923 29586 5979 29642
rect 6047 29586 6103 29642
rect 6171 29586 6227 29642
rect 4435 29462 4491 29518
rect 4559 29462 4615 29518
rect 4683 29462 4739 29518
rect 4807 29462 4863 29518
rect 4931 29462 4987 29518
rect 5055 29462 5111 29518
rect 5179 29462 5235 29518
rect 5303 29462 5359 29518
rect 5427 29462 5483 29518
rect 5551 29462 5607 29518
rect 5675 29462 5731 29518
rect 5799 29462 5855 29518
rect 5923 29462 5979 29518
rect 6047 29462 6103 29518
rect 6171 29462 6227 29518
rect 4435 29338 4491 29394
rect 4559 29338 4615 29394
rect 4683 29338 4739 29394
rect 4807 29338 4863 29394
rect 4931 29338 4987 29394
rect 5055 29338 5111 29394
rect 5179 29338 5235 29394
rect 5303 29338 5359 29394
rect 5427 29338 5483 29394
rect 5551 29338 5607 29394
rect 5675 29338 5731 29394
rect 5799 29338 5855 29394
rect 5923 29338 5979 29394
rect 6047 29338 6103 29394
rect 6171 29338 6227 29394
rect 4435 29214 4491 29270
rect 4559 29214 4615 29270
rect 4683 29214 4739 29270
rect 4807 29214 4863 29270
rect 4931 29214 4987 29270
rect 5055 29214 5111 29270
rect 5179 29214 5235 29270
rect 5303 29214 5359 29270
rect 5427 29214 5483 29270
rect 5551 29214 5607 29270
rect 5675 29214 5731 29270
rect 5799 29214 5855 29270
rect 5923 29214 5979 29270
rect 6047 29214 6103 29270
rect 6171 29214 6227 29270
rect 4435 29090 4491 29146
rect 4559 29090 4615 29146
rect 4683 29090 4739 29146
rect 4807 29090 4863 29146
rect 4931 29090 4987 29146
rect 5055 29090 5111 29146
rect 5179 29090 5235 29146
rect 5303 29090 5359 29146
rect 5427 29090 5483 29146
rect 5551 29090 5607 29146
rect 5675 29090 5731 29146
rect 5799 29090 5855 29146
rect 5923 29090 5979 29146
rect 6047 29090 6103 29146
rect 6171 29090 6227 29146
rect 4435 28966 4491 29022
rect 4559 28966 4615 29022
rect 4683 28966 4739 29022
rect 4807 28966 4863 29022
rect 4931 28966 4987 29022
rect 5055 28966 5111 29022
rect 5179 28966 5235 29022
rect 5303 28966 5359 29022
rect 5427 28966 5483 29022
rect 5551 28966 5607 29022
rect 5675 28966 5731 29022
rect 5799 28966 5855 29022
rect 5923 28966 5979 29022
rect 6047 28966 6103 29022
rect 6171 28966 6227 29022
rect 4435 28842 4491 28898
rect 4559 28842 4615 28898
rect 4683 28842 4739 28898
rect 4807 28842 4863 28898
rect 4931 28842 4987 28898
rect 5055 28842 5111 28898
rect 5179 28842 5235 28898
rect 5303 28842 5359 28898
rect 5427 28842 5483 28898
rect 5551 28842 5607 28898
rect 5675 28842 5731 28898
rect 5799 28842 5855 28898
rect 5923 28842 5979 28898
rect 6047 28842 6103 28898
rect 6171 28842 6227 28898
rect 7562 31694 7618 31750
rect 7686 31694 7742 31750
rect 7810 31694 7866 31750
rect 7934 31694 7990 31750
rect 8058 31694 8114 31750
rect 8182 31694 8238 31750
rect 8306 31694 8362 31750
rect 8430 31694 8486 31750
rect 8554 31694 8610 31750
rect 7562 31570 7618 31626
rect 7686 31570 7742 31626
rect 7810 31570 7866 31626
rect 7934 31570 7990 31626
rect 8058 31570 8114 31626
rect 8182 31570 8238 31626
rect 8306 31570 8362 31626
rect 8430 31570 8486 31626
rect 8554 31570 8610 31626
rect 7562 31446 7618 31502
rect 7686 31446 7742 31502
rect 7810 31446 7866 31502
rect 7934 31446 7990 31502
rect 8058 31446 8114 31502
rect 8182 31446 8238 31502
rect 8306 31446 8362 31502
rect 8430 31446 8486 31502
rect 8554 31446 8610 31502
rect 7562 31322 7618 31378
rect 7686 31322 7742 31378
rect 7810 31322 7866 31378
rect 7934 31322 7990 31378
rect 8058 31322 8114 31378
rect 8182 31322 8238 31378
rect 8306 31322 8362 31378
rect 8430 31322 8486 31378
rect 8554 31322 8610 31378
rect 7562 31198 7618 31254
rect 7686 31198 7742 31254
rect 7810 31198 7866 31254
rect 7934 31198 7990 31254
rect 8058 31198 8114 31254
rect 8182 31198 8238 31254
rect 8306 31198 8362 31254
rect 8430 31198 8486 31254
rect 8554 31198 8610 31254
rect 7562 31074 7618 31130
rect 7686 31074 7742 31130
rect 7810 31074 7866 31130
rect 7934 31074 7990 31130
rect 8058 31074 8114 31130
rect 8182 31074 8238 31130
rect 8306 31074 8362 31130
rect 8430 31074 8486 31130
rect 8554 31074 8610 31130
rect 7562 30950 7618 31006
rect 7686 30950 7742 31006
rect 7810 30950 7866 31006
rect 7934 30950 7990 31006
rect 8058 30950 8114 31006
rect 8182 30950 8238 31006
rect 8306 30950 8362 31006
rect 8430 30950 8486 31006
rect 8554 30950 8610 31006
rect 7562 30826 7618 30882
rect 7686 30826 7742 30882
rect 7810 30826 7866 30882
rect 7934 30826 7990 30882
rect 8058 30826 8114 30882
rect 8182 30826 8238 30882
rect 8306 30826 8362 30882
rect 8430 30826 8486 30882
rect 8554 30826 8610 30882
rect 7562 30702 7618 30758
rect 7686 30702 7742 30758
rect 7810 30702 7866 30758
rect 7934 30702 7990 30758
rect 8058 30702 8114 30758
rect 8182 30702 8238 30758
rect 8306 30702 8362 30758
rect 8430 30702 8486 30758
rect 8554 30702 8610 30758
rect 7562 30578 7618 30634
rect 7686 30578 7742 30634
rect 7810 30578 7866 30634
rect 7934 30578 7990 30634
rect 8058 30578 8114 30634
rect 8182 30578 8238 30634
rect 8306 30578 8362 30634
rect 8430 30578 8486 30634
rect 8554 30578 8610 30634
rect 7562 30454 7618 30510
rect 7686 30454 7742 30510
rect 7810 30454 7866 30510
rect 7934 30454 7990 30510
rect 8058 30454 8114 30510
rect 8182 30454 8238 30510
rect 8306 30454 8362 30510
rect 8430 30454 8486 30510
rect 8554 30454 8610 30510
rect 7562 30330 7618 30386
rect 7686 30330 7742 30386
rect 7810 30330 7866 30386
rect 7934 30330 7990 30386
rect 8058 30330 8114 30386
rect 8182 30330 8238 30386
rect 8306 30330 8362 30386
rect 8430 30330 8486 30386
rect 8554 30330 8610 30386
rect 7562 30206 7618 30262
rect 7686 30206 7742 30262
rect 7810 30206 7866 30262
rect 7934 30206 7990 30262
rect 8058 30206 8114 30262
rect 8182 30206 8238 30262
rect 8306 30206 8362 30262
rect 8430 30206 8486 30262
rect 8554 30206 8610 30262
rect 7562 30082 7618 30138
rect 7686 30082 7742 30138
rect 7810 30082 7866 30138
rect 7934 30082 7990 30138
rect 8058 30082 8114 30138
rect 8182 30082 8238 30138
rect 8306 30082 8362 30138
rect 8430 30082 8486 30138
rect 8554 30082 8610 30138
rect 7562 29958 7618 30014
rect 7686 29958 7742 30014
rect 7810 29958 7866 30014
rect 7934 29958 7990 30014
rect 8058 29958 8114 30014
rect 8182 29958 8238 30014
rect 8306 29958 8362 30014
rect 8430 29958 8486 30014
rect 8554 29958 8610 30014
rect 7562 29834 7618 29890
rect 7686 29834 7742 29890
rect 7810 29834 7866 29890
rect 7934 29834 7990 29890
rect 8058 29834 8114 29890
rect 8182 29834 8238 29890
rect 8306 29834 8362 29890
rect 8430 29834 8486 29890
rect 8554 29834 8610 29890
rect 7562 29710 7618 29766
rect 7686 29710 7742 29766
rect 7810 29710 7866 29766
rect 7934 29710 7990 29766
rect 8058 29710 8114 29766
rect 8182 29710 8238 29766
rect 8306 29710 8362 29766
rect 8430 29710 8486 29766
rect 8554 29710 8610 29766
rect 7562 29586 7618 29642
rect 7686 29586 7742 29642
rect 7810 29586 7866 29642
rect 7934 29586 7990 29642
rect 8058 29586 8114 29642
rect 8182 29586 8238 29642
rect 8306 29586 8362 29642
rect 8430 29586 8486 29642
rect 8554 29586 8610 29642
rect 7562 29462 7618 29518
rect 7686 29462 7742 29518
rect 7810 29462 7866 29518
rect 7934 29462 7990 29518
rect 8058 29462 8114 29518
rect 8182 29462 8238 29518
rect 8306 29462 8362 29518
rect 8430 29462 8486 29518
rect 8554 29462 8610 29518
rect 7562 29338 7618 29394
rect 7686 29338 7742 29394
rect 7810 29338 7866 29394
rect 7934 29338 7990 29394
rect 8058 29338 8114 29394
rect 8182 29338 8238 29394
rect 8306 29338 8362 29394
rect 8430 29338 8486 29394
rect 8554 29338 8610 29394
rect 7562 29214 7618 29270
rect 7686 29214 7742 29270
rect 7810 29214 7866 29270
rect 7934 29214 7990 29270
rect 8058 29214 8114 29270
rect 8182 29214 8238 29270
rect 8306 29214 8362 29270
rect 8430 29214 8486 29270
rect 8554 29214 8610 29270
rect 7562 29090 7618 29146
rect 7686 29090 7742 29146
rect 7810 29090 7866 29146
rect 7934 29090 7990 29146
rect 8058 29090 8114 29146
rect 8182 29090 8238 29146
rect 8306 29090 8362 29146
rect 8430 29090 8486 29146
rect 8554 29090 8610 29146
rect 7562 28966 7618 29022
rect 7686 28966 7742 29022
rect 7810 28966 7866 29022
rect 7934 28966 7990 29022
rect 8058 28966 8114 29022
rect 8182 28966 8238 29022
rect 8306 28966 8362 29022
rect 8430 28966 8486 29022
rect 8554 28966 8610 29022
rect 7562 28842 7618 28898
rect 7686 28842 7742 28898
rect 7810 28842 7866 28898
rect 7934 28842 7990 28898
rect 8058 28842 8114 28898
rect 8182 28842 8238 28898
rect 8306 28842 8362 28898
rect 8430 28842 8486 28898
rect 8554 28842 8610 28898
rect 10679 31694 10735 31750
rect 10803 31694 10859 31750
rect 10927 31694 10983 31750
rect 11051 31694 11107 31750
rect 11175 31694 11231 31750
rect 11299 31694 11355 31750
rect 11423 31694 11479 31750
rect 11547 31694 11603 31750
rect 11671 31694 11727 31750
rect 11795 31694 11851 31750
rect 11919 31694 11975 31750
rect 12043 31694 12099 31750
rect 12167 31694 12223 31750
rect 12291 31694 12347 31750
rect 12415 31694 12471 31750
rect 10679 31570 10735 31626
rect 10803 31570 10859 31626
rect 10927 31570 10983 31626
rect 11051 31570 11107 31626
rect 11175 31570 11231 31626
rect 11299 31570 11355 31626
rect 11423 31570 11479 31626
rect 11547 31570 11603 31626
rect 11671 31570 11727 31626
rect 11795 31570 11851 31626
rect 11919 31570 11975 31626
rect 12043 31570 12099 31626
rect 12167 31570 12223 31626
rect 12291 31570 12347 31626
rect 12415 31570 12471 31626
rect 10679 31446 10735 31502
rect 10803 31446 10859 31502
rect 10927 31446 10983 31502
rect 11051 31446 11107 31502
rect 11175 31446 11231 31502
rect 11299 31446 11355 31502
rect 11423 31446 11479 31502
rect 11547 31446 11603 31502
rect 11671 31446 11727 31502
rect 11795 31446 11851 31502
rect 11919 31446 11975 31502
rect 12043 31446 12099 31502
rect 12167 31446 12223 31502
rect 12291 31446 12347 31502
rect 12415 31446 12471 31502
rect 10679 31322 10735 31378
rect 10803 31322 10859 31378
rect 10927 31322 10983 31378
rect 11051 31322 11107 31378
rect 11175 31322 11231 31378
rect 11299 31322 11355 31378
rect 11423 31322 11479 31378
rect 11547 31322 11603 31378
rect 11671 31322 11727 31378
rect 11795 31322 11851 31378
rect 11919 31322 11975 31378
rect 12043 31322 12099 31378
rect 12167 31322 12223 31378
rect 12291 31322 12347 31378
rect 12415 31322 12471 31378
rect 10679 31198 10735 31254
rect 10803 31198 10859 31254
rect 10927 31198 10983 31254
rect 11051 31198 11107 31254
rect 11175 31198 11231 31254
rect 11299 31198 11355 31254
rect 11423 31198 11479 31254
rect 11547 31198 11603 31254
rect 11671 31198 11727 31254
rect 11795 31198 11851 31254
rect 11919 31198 11975 31254
rect 12043 31198 12099 31254
rect 12167 31198 12223 31254
rect 12291 31198 12347 31254
rect 12415 31198 12471 31254
rect 10679 31074 10735 31130
rect 10803 31074 10859 31130
rect 10927 31074 10983 31130
rect 11051 31074 11107 31130
rect 11175 31074 11231 31130
rect 11299 31074 11355 31130
rect 11423 31074 11479 31130
rect 11547 31074 11603 31130
rect 11671 31074 11727 31130
rect 11795 31074 11851 31130
rect 11919 31074 11975 31130
rect 12043 31074 12099 31130
rect 12167 31074 12223 31130
rect 12291 31074 12347 31130
rect 12415 31074 12471 31130
rect 10679 30950 10735 31006
rect 10803 30950 10859 31006
rect 10927 30950 10983 31006
rect 11051 30950 11107 31006
rect 11175 30950 11231 31006
rect 11299 30950 11355 31006
rect 11423 30950 11479 31006
rect 11547 30950 11603 31006
rect 11671 30950 11727 31006
rect 11795 30950 11851 31006
rect 11919 30950 11975 31006
rect 12043 30950 12099 31006
rect 12167 30950 12223 31006
rect 12291 30950 12347 31006
rect 12415 30950 12471 31006
rect 10679 30826 10735 30882
rect 10803 30826 10859 30882
rect 10927 30826 10983 30882
rect 11051 30826 11107 30882
rect 11175 30826 11231 30882
rect 11299 30826 11355 30882
rect 11423 30826 11479 30882
rect 11547 30826 11603 30882
rect 11671 30826 11727 30882
rect 11795 30826 11851 30882
rect 11919 30826 11975 30882
rect 12043 30826 12099 30882
rect 12167 30826 12223 30882
rect 12291 30826 12347 30882
rect 12415 30826 12471 30882
rect 10679 30702 10735 30758
rect 10803 30702 10859 30758
rect 10927 30702 10983 30758
rect 11051 30702 11107 30758
rect 11175 30702 11231 30758
rect 11299 30702 11355 30758
rect 11423 30702 11479 30758
rect 11547 30702 11603 30758
rect 11671 30702 11727 30758
rect 11795 30702 11851 30758
rect 11919 30702 11975 30758
rect 12043 30702 12099 30758
rect 12167 30702 12223 30758
rect 12291 30702 12347 30758
rect 12415 30702 12471 30758
rect 10679 30578 10735 30634
rect 10803 30578 10859 30634
rect 10927 30578 10983 30634
rect 11051 30578 11107 30634
rect 11175 30578 11231 30634
rect 11299 30578 11355 30634
rect 11423 30578 11479 30634
rect 11547 30578 11603 30634
rect 11671 30578 11727 30634
rect 11795 30578 11851 30634
rect 11919 30578 11975 30634
rect 12043 30578 12099 30634
rect 12167 30578 12223 30634
rect 12291 30578 12347 30634
rect 12415 30578 12471 30634
rect 10679 30454 10735 30510
rect 10803 30454 10859 30510
rect 10927 30454 10983 30510
rect 11051 30454 11107 30510
rect 11175 30454 11231 30510
rect 11299 30454 11355 30510
rect 11423 30454 11479 30510
rect 11547 30454 11603 30510
rect 11671 30454 11727 30510
rect 11795 30454 11851 30510
rect 11919 30454 11975 30510
rect 12043 30454 12099 30510
rect 12167 30454 12223 30510
rect 12291 30454 12347 30510
rect 12415 30454 12471 30510
rect 10679 30330 10735 30386
rect 10803 30330 10859 30386
rect 10927 30330 10983 30386
rect 11051 30330 11107 30386
rect 11175 30330 11231 30386
rect 11299 30330 11355 30386
rect 11423 30330 11479 30386
rect 11547 30330 11603 30386
rect 11671 30330 11727 30386
rect 11795 30330 11851 30386
rect 11919 30330 11975 30386
rect 12043 30330 12099 30386
rect 12167 30330 12223 30386
rect 12291 30330 12347 30386
rect 12415 30330 12471 30386
rect 10679 30206 10735 30262
rect 10803 30206 10859 30262
rect 10927 30206 10983 30262
rect 11051 30206 11107 30262
rect 11175 30206 11231 30262
rect 11299 30206 11355 30262
rect 11423 30206 11479 30262
rect 11547 30206 11603 30262
rect 11671 30206 11727 30262
rect 11795 30206 11851 30262
rect 11919 30206 11975 30262
rect 12043 30206 12099 30262
rect 12167 30206 12223 30262
rect 12291 30206 12347 30262
rect 12415 30206 12471 30262
rect 10679 30082 10735 30138
rect 10803 30082 10859 30138
rect 10927 30082 10983 30138
rect 11051 30082 11107 30138
rect 11175 30082 11231 30138
rect 11299 30082 11355 30138
rect 11423 30082 11479 30138
rect 11547 30082 11603 30138
rect 11671 30082 11727 30138
rect 11795 30082 11851 30138
rect 11919 30082 11975 30138
rect 12043 30082 12099 30138
rect 12167 30082 12223 30138
rect 12291 30082 12347 30138
rect 12415 30082 12471 30138
rect 10679 29958 10735 30014
rect 10803 29958 10859 30014
rect 10927 29958 10983 30014
rect 11051 29958 11107 30014
rect 11175 29958 11231 30014
rect 11299 29958 11355 30014
rect 11423 29958 11479 30014
rect 11547 29958 11603 30014
rect 11671 29958 11727 30014
rect 11795 29958 11851 30014
rect 11919 29958 11975 30014
rect 12043 29958 12099 30014
rect 12167 29958 12223 30014
rect 12291 29958 12347 30014
rect 12415 29958 12471 30014
rect 10679 29834 10735 29890
rect 10803 29834 10859 29890
rect 10927 29834 10983 29890
rect 11051 29834 11107 29890
rect 11175 29834 11231 29890
rect 11299 29834 11355 29890
rect 11423 29834 11479 29890
rect 11547 29834 11603 29890
rect 11671 29834 11727 29890
rect 11795 29834 11851 29890
rect 11919 29834 11975 29890
rect 12043 29834 12099 29890
rect 12167 29834 12223 29890
rect 12291 29834 12347 29890
rect 12415 29834 12471 29890
rect 10679 29710 10735 29766
rect 10803 29710 10859 29766
rect 10927 29710 10983 29766
rect 11051 29710 11107 29766
rect 11175 29710 11231 29766
rect 11299 29710 11355 29766
rect 11423 29710 11479 29766
rect 11547 29710 11603 29766
rect 11671 29710 11727 29766
rect 11795 29710 11851 29766
rect 11919 29710 11975 29766
rect 12043 29710 12099 29766
rect 12167 29710 12223 29766
rect 12291 29710 12347 29766
rect 12415 29710 12471 29766
rect 10679 29586 10735 29642
rect 10803 29586 10859 29642
rect 10927 29586 10983 29642
rect 11051 29586 11107 29642
rect 11175 29586 11231 29642
rect 11299 29586 11355 29642
rect 11423 29586 11479 29642
rect 11547 29586 11603 29642
rect 11671 29586 11727 29642
rect 11795 29586 11851 29642
rect 11919 29586 11975 29642
rect 12043 29586 12099 29642
rect 12167 29586 12223 29642
rect 12291 29586 12347 29642
rect 12415 29586 12471 29642
rect 10679 29462 10735 29518
rect 10803 29462 10859 29518
rect 10927 29462 10983 29518
rect 11051 29462 11107 29518
rect 11175 29462 11231 29518
rect 11299 29462 11355 29518
rect 11423 29462 11479 29518
rect 11547 29462 11603 29518
rect 11671 29462 11727 29518
rect 11795 29462 11851 29518
rect 11919 29462 11975 29518
rect 12043 29462 12099 29518
rect 12167 29462 12223 29518
rect 12291 29462 12347 29518
rect 12415 29462 12471 29518
rect 10679 29338 10735 29394
rect 10803 29338 10859 29394
rect 10927 29338 10983 29394
rect 11051 29338 11107 29394
rect 11175 29338 11231 29394
rect 11299 29338 11355 29394
rect 11423 29338 11479 29394
rect 11547 29338 11603 29394
rect 11671 29338 11727 29394
rect 11795 29338 11851 29394
rect 11919 29338 11975 29394
rect 12043 29338 12099 29394
rect 12167 29338 12223 29394
rect 12291 29338 12347 29394
rect 12415 29338 12471 29394
rect 10679 29214 10735 29270
rect 10803 29214 10859 29270
rect 10927 29214 10983 29270
rect 11051 29214 11107 29270
rect 11175 29214 11231 29270
rect 11299 29214 11355 29270
rect 11423 29214 11479 29270
rect 11547 29214 11603 29270
rect 11671 29214 11727 29270
rect 11795 29214 11851 29270
rect 11919 29214 11975 29270
rect 12043 29214 12099 29270
rect 12167 29214 12223 29270
rect 12291 29214 12347 29270
rect 12415 29214 12471 29270
rect 10679 29090 10735 29146
rect 10803 29090 10859 29146
rect 10927 29090 10983 29146
rect 11051 29090 11107 29146
rect 11175 29090 11231 29146
rect 11299 29090 11355 29146
rect 11423 29090 11479 29146
rect 11547 29090 11603 29146
rect 11671 29090 11727 29146
rect 11795 29090 11851 29146
rect 11919 29090 11975 29146
rect 12043 29090 12099 29146
rect 12167 29090 12223 29146
rect 12291 29090 12347 29146
rect 12415 29090 12471 29146
rect 10679 28966 10735 29022
rect 10803 28966 10859 29022
rect 10927 28966 10983 29022
rect 11051 28966 11107 29022
rect 11175 28966 11231 29022
rect 11299 28966 11355 29022
rect 11423 28966 11479 29022
rect 11547 28966 11603 29022
rect 11671 28966 11727 29022
rect 11795 28966 11851 29022
rect 11919 28966 11975 29022
rect 12043 28966 12099 29022
rect 12167 28966 12223 29022
rect 12291 28966 12347 29022
rect 12415 28966 12471 29022
rect 10679 28842 10735 28898
rect 10803 28842 10859 28898
rect 10927 28842 10983 28898
rect 11051 28842 11107 28898
rect 11175 28842 11231 28898
rect 11299 28842 11355 28898
rect 11423 28842 11479 28898
rect 11547 28842 11603 28898
rect 11671 28842 11727 28898
rect 11795 28842 11851 28898
rect 11919 28842 11975 28898
rect 12043 28842 12099 28898
rect 12167 28842 12223 28898
rect 12291 28842 12347 28898
rect 12415 28842 12471 28898
rect 1499 28742 1555 28798
rect 1499 28618 1555 28674
rect 1499 28494 1555 28550
rect 1499 28370 1555 28426
rect 1499 28246 1555 28302
rect 1499 28122 1555 28178
rect 1499 27998 1555 28054
rect 1499 27874 1555 27930
rect 1499 27750 1555 27806
rect 1499 27626 1555 27682
rect 1499 27502 1555 27558
rect 1499 27378 1555 27434
rect 1499 27254 1555 27310
rect 1623 28752 1679 28808
rect 1623 28628 1679 28684
rect 1623 28504 1679 28560
rect 1623 28380 1679 28436
rect 1623 28256 1679 28312
rect 1623 28132 1679 28188
rect 1623 28008 1679 28064
rect 1623 27884 1679 27940
rect 1623 27760 1679 27816
rect 1623 27636 1679 27692
rect 1623 27512 1679 27568
rect 1623 27388 1679 27444
rect 1623 27264 1679 27320
rect 1747 28597 1803 28653
rect 1747 28473 1803 28529
rect 1747 28349 1803 28405
rect 1747 28225 1803 28281
rect 1747 28101 1803 28157
rect 1747 27977 1803 28033
rect 1747 27853 1803 27909
rect 1747 27729 1803 27785
rect 1747 27605 1803 27661
rect 1747 27481 1803 27537
rect 1747 27357 1803 27413
rect 1747 27233 1803 27289
rect 1871 28483 1927 28539
rect 1871 28359 1927 28415
rect 1871 28235 1927 28291
rect 1871 28111 1927 28167
rect 1871 27987 1927 28043
rect 1871 27863 1927 27919
rect 1871 27739 1927 27795
rect 1871 27615 1927 27671
rect 1871 27491 1927 27547
rect 1871 27367 1927 27423
rect 1871 27243 1927 27299
rect 1995 28481 2051 28537
rect 1995 28357 2051 28413
rect 1995 28233 2051 28289
rect 1995 28109 2051 28165
rect 1995 27985 2051 28041
rect 1995 27861 2051 27917
rect 1995 27737 2051 27793
rect 1995 27613 2051 27669
rect 1995 27489 2051 27545
rect 1995 27365 2051 27421
rect 1995 27241 2051 27297
rect 4435 28488 4491 28544
rect 4559 28488 4615 28544
rect 4683 28488 4739 28544
rect 4807 28488 4863 28544
rect 4931 28488 4987 28544
rect 5055 28488 5111 28544
rect 5179 28488 5235 28544
rect 5303 28488 5359 28544
rect 5427 28488 5483 28544
rect 5551 28488 5607 28544
rect 5675 28488 5731 28544
rect 5799 28488 5855 28544
rect 5923 28488 5979 28544
rect 6047 28488 6103 28544
rect 6171 28488 6227 28544
rect 4435 28364 4491 28420
rect 4559 28364 4615 28420
rect 4683 28364 4739 28420
rect 4807 28364 4863 28420
rect 4931 28364 4987 28420
rect 5055 28364 5111 28420
rect 5179 28364 5235 28420
rect 5303 28364 5359 28420
rect 5427 28364 5483 28420
rect 5551 28364 5607 28420
rect 5675 28364 5731 28420
rect 5799 28364 5855 28420
rect 5923 28364 5979 28420
rect 6047 28364 6103 28420
rect 6171 28364 6227 28420
rect 4435 28240 4491 28296
rect 4559 28240 4615 28296
rect 4683 28240 4739 28296
rect 4807 28240 4863 28296
rect 4931 28240 4987 28296
rect 5055 28240 5111 28296
rect 5179 28240 5235 28296
rect 5303 28240 5359 28296
rect 5427 28240 5483 28296
rect 5551 28240 5607 28296
rect 5675 28240 5731 28296
rect 5799 28240 5855 28296
rect 5923 28240 5979 28296
rect 6047 28240 6103 28296
rect 6171 28240 6227 28296
rect 4435 28116 4491 28172
rect 4559 28116 4615 28172
rect 4683 28116 4739 28172
rect 4807 28116 4863 28172
rect 4931 28116 4987 28172
rect 5055 28116 5111 28172
rect 5179 28116 5235 28172
rect 5303 28116 5359 28172
rect 5427 28116 5483 28172
rect 5551 28116 5607 28172
rect 5675 28116 5731 28172
rect 5799 28116 5855 28172
rect 5923 28116 5979 28172
rect 6047 28116 6103 28172
rect 6171 28116 6227 28172
rect 4435 27992 4491 28048
rect 4559 27992 4615 28048
rect 4683 27992 4739 28048
rect 4807 27992 4863 28048
rect 4931 27992 4987 28048
rect 5055 27992 5111 28048
rect 5179 27992 5235 28048
rect 5303 27992 5359 28048
rect 5427 27992 5483 28048
rect 5551 27992 5607 28048
rect 5675 27992 5731 28048
rect 5799 27992 5855 28048
rect 5923 27992 5979 28048
rect 6047 27992 6103 28048
rect 6171 27992 6227 28048
rect 4435 27868 4491 27924
rect 4559 27868 4615 27924
rect 4683 27868 4739 27924
rect 4807 27868 4863 27924
rect 4931 27868 4987 27924
rect 5055 27868 5111 27924
rect 5179 27868 5235 27924
rect 5303 27868 5359 27924
rect 5427 27868 5483 27924
rect 5551 27868 5607 27924
rect 5675 27868 5731 27924
rect 5799 27868 5855 27924
rect 5923 27868 5979 27924
rect 6047 27868 6103 27924
rect 6171 27868 6227 27924
rect 4435 27744 4491 27800
rect 4559 27744 4615 27800
rect 4683 27744 4739 27800
rect 4807 27744 4863 27800
rect 4931 27744 4987 27800
rect 5055 27744 5111 27800
rect 5179 27744 5235 27800
rect 5303 27744 5359 27800
rect 5427 27744 5483 27800
rect 5551 27744 5607 27800
rect 5675 27744 5731 27800
rect 5799 27744 5855 27800
rect 5923 27744 5979 27800
rect 6047 27744 6103 27800
rect 6171 27744 6227 27800
rect 4435 27620 4491 27676
rect 4559 27620 4615 27676
rect 4683 27620 4739 27676
rect 4807 27620 4863 27676
rect 4931 27620 4987 27676
rect 5055 27620 5111 27676
rect 5179 27620 5235 27676
rect 5303 27620 5359 27676
rect 5427 27620 5483 27676
rect 5551 27620 5607 27676
rect 5675 27620 5731 27676
rect 5799 27620 5855 27676
rect 5923 27620 5979 27676
rect 6047 27620 6103 27676
rect 6171 27620 6227 27676
rect 4435 27496 4491 27552
rect 4559 27496 4615 27552
rect 4683 27496 4739 27552
rect 4807 27496 4863 27552
rect 4931 27496 4987 27552
rect 5055 27496 5111 27552
rect 5179 27496 5235 27552
rect 5303 27496 5359 27552
rect 5427 27496 5483 27552
rect 5551 27496 5607 27552
rect 5675 27496 5731 27552
rect 5799 27496 5855 27552
rect 5923 27496 5979 27552
rect 6047 27496 6103 27552
rect 6171 27496 6227 27552
rect 4435 27372 4491 27428
rect 4559 27372 4615 27428
rect 4683 27372 4739 27428
rect 4807 27372 4863 27428
rect 4931 27372 4987 27428
rect 5055 27372 5111 27428
rect 5179 27372 5235 27428
rect 5303 27372 5359 27428
rect 5427 27372 5483 27428
rect 5551 27372 5607 27428
rect 5675 27372 5731 27428
rect 5799 27372 5855 27428
rect 5923 27372 5979 27428
rect 6047 27372 6103 27428
rect 6171 27372 6227 27428
rect 4435 27248 4491 27304
rect 4559 27248 4615 27304
rect 4683 27248 4739 27304
rect 4807 27248 4863 27304
rect 4931 27248 4987 27304
rect 5055 27248 5111 27304
rect 5179 27248 5235 27304
rect 5303 27248 5359 27304
rect 5427 27248 5483 27304
rect 5551 27248 5607 27304
rect 5675 27248 5731 27304
rect 5799 27248 5855 27304
rect 5923 27248 5979 27304
rect 6047 27248 6103 27304
rect 6171 27248 6227 27304
rect 7562 28488 7618 28544
rect 7686 28488 7742 28544
rect 7810 28488 7866 28544
rect 7934 28488 7990 28544
rect 8058 28488 8114 28544
rect 8182 28488 8238 28544
rect 8306 28488 8362 28544
rect 8430 28488 8486 28544
rect 8554 28488 8610 28544
rect 7562 28364 7618 28420
rect 7686 28364 7742 28420
rect 7810 28364 7866 28420
rect 7934 28364 7990 28420
rect 8058 28364 8114 28420
rect 8182 28364 8238 28420
rect 8306 28364 8362 28420
rect 8430 28364 8486 28420
rect 8554 28364 8610 28420
rect 7562 28240 7618 28296
rect 7686 28240 7742 28296
rect 7810 28240 7866 28296
rect 7934 28240 7990 28296
rect 8058 28240 8114 28296
rect 8182 28240 8238 28296
rect 8306 28240 8362 28296
rect 8430 28240 8486 28296
rect 8554 28240 8610 28296
rect 7562 28116 7618 28172
rect 7686 28116 7742 28172
rect 7810 28116 7866 28172
rect 7934 28116 7990 28172
rect 8058 28116 8114 28172
rect 8182 28116 8238 28172
rect 8306 28116 8362 28172
rect 8430 28116 8486 28172
rect 8554 28116 8610 28172
rect 7562 27992 7618 28048
rect 7686 27992 7742 28048
rect 7810 27992 7866 28048
rect 7934 27992 7990 28048
rect 8058 27992 8114 28048
rect 8182 27992 8238 28048
rect 8306 27992 8362 28048
rect 8430 27992 8486 28048
rect 8554 27992 8610 28048
rect 7562 27868 7618 27924
rect 7686 27868 7742 27924
rect 7810 27868 7866 27924
rect 7934 27868 7990 27924
rect 8058 27868 8114 27924
rect 8182 27868 8238 27924
rect 8306 27868 8362 27924
rect 8430 27868 8486 27924
rect 8554 27868 8610 27924
rect 7562 27744 7618 27800
rect 7686 27744 7742 27800
rect 7810 27744 7866 27800
rect 7934 27744 7990 27800
rect 8058 27744 8114 27800
rect 8182 27744 8238 27800
rect 8306 27744 8362 27800
rect 8430 27744 8486 27800
rect 8554 27744 8610 27800
rect 7562 27620 7618 27676
rect 7686 27620 7742 27676
rect 7810 27620 7866 27676
rect 7934 27620 7990 27676
rect 8058 27620 8114 27676
rect 8182 27620 8238 27676
rect 8306 27620 8362 27676
rect 8430 27620 8486 27676
rect 8554 27620 8610 27676
rect 7562 27496 7618 27552
rect 7686 27496 7742 27552
rect 7810 27496 7866 27552
rect 7934 27496 7990 27552
rect 8058 27496 8114 27552
rect 8182 27496 8238 27552
rect 8306 27496 8362 27552
rect 8430 27496 8486 27552
rect 8554 27496 8610 27552
rect 7562 27372 7618 27428
rect 7686 27372 7742 27428
rect 7810 27372 7866 27428
rect 7934 27372 7990 27428
rect 8058 27372 8114 27428
rect 8182 27372 8238 27428
rect 8306 27372 8362 27428
rect 8430 27372 8486 27428
rect 8554 27372 8610 27428
rect 7562 27248 7618 27304
rect 7686 27248 7742 27304
rect 7810 27248 7866 27304
rect 7934 27248 7990 27304
rect 8058 27248 8114 27304
rect 8182 27248 8238 27304
rect 8306 27248 8362 27304
rect 8430 27248 8486 27304
rect 8554 27248 8610 27304
rect 10679 28488 10735 28544
rect 10803 28488 10859 28544
rect 10927 28488 10983 28544
rect 11051 28488 11107 28544
rect 11175 28488 11231 28544
rect 11299 28488 11355 28544
rect 11423 28488 11479 28544
rect 11547 28488 11603 28544
rect 11671 28488 11727 28544
rect 11795 28488 11851 28544
rect 11919 28488 11975 28544
rect 12043 28488 12099 28544
rect 12167 28488 12223 28544
rect 12291 28488 12347 28544
rect 12415 28488 12471 28544
rect 10679 28364 10735 28420
rect 10803 28364 10859 28420
rect 10927 28364 10983 28420
rect 11051 28364 11107 28420
rect 11175 28364 11231 28420
rect 11299 28364 11355 28420
rect 11423 28364 11479 28420
rect 11547 28364 11603 28420
rect 11671 28364 11727 28420
rect 11795 28364 11851 28420
rect 11919 28364 11975 28420
rect 12043 28364 12099 28420
rect 12167 28364 12223 28420
rect 12291 28364 12347 28420
rect 12415 28364 12471 28420
rect 10679 28240 10735 28296
rect 10803 28240 10859 28296
rect 10927 28240 10983 28296
rect 11051 28240 11107 28296
rect 11175 28240 11231 28296
rect 11299 28240 11355 28296
rect 11423 28240 11479 28296
rect 11547 28240 11603 28296
rect 11671 28240 11727 28296
rect 11795 28240 11851 28296
rect 11919 28240 11975 28296
rect 12043 28240 12099 28296
rect 12167 28240 12223 28296
rect 12291 28240 12347 28296
rect 12415 28240 12471 28296
rect 10679 28116 10735 28172
rect 10803 28116 10859 28172
rect 10927 28116 10983 28172
rect 11051 28116 11107 28172
rect 11175 28116 11231 28172
rect 11299 28116 11355 28172
rect 11423 28116 11479 28172
rect 11547 28116 11603 28172
rect 11671 28116 11727 28172
rect 11795 28116 11851 28172
rect 11919 28116 11975 28172
rect 12043 28116 12099 28172
rect 12167 28116 12223 28172
rect 12291 28116 12347 28172
rect 12415 28116 12471 28172
rect 10679 27992 10735 28048
rect 10803 27992 10859 28048
rect 10927 27992 10983 28048
rect 11051 27992 11107 28048
rect 11175 27992 11231 28048
rect 11299 27992 11355 28048
rect 11423 27992 11479 28048
rect 11547 27992 11603 28048
rect 11671 27992 11727 28048
rect 11795 27992 11851 28048
rect 11919 27992 11975 28048
rect 12043 27992 12099 28048
rect 12167 27992 12223 28048
rect 12291 27992 12347 28048
rect 12415 27992 12471 28048
rect 10679 27868 10735 27924
rect 10803 27868 10859 27924
rect 10927 27868 10983 27924
rect 11051 27868 11107 27924
rect 11175 27868 11231 27924
rect 11299 27868 11355 27924
rect 11423 27868 11479 27924
rect 11547 27868 11603 27924
rect 11671 27868 11727 27924
rect 11795 27868 11851 27924
rect 11919 27868 11975 27924
rect 12043 27868 12099 27924
rect 12167 27868 12223 27924
rect 12291 27868 12347 27924
rect 12415 27868 12471 27924
rect 10679 27744 10735 27800
rect 10803 27744 10859 27800
rect 10927 27744 10983 27800
rect 11051 27744 11107 27800
rect 11175 27744 11231 27800
rect 11299 27744 11355 27800
rect 11423 27744 11479 27800
rect 11547 27744 11603 27800
rect 11671 27744 11727 27800
rect 11795 27744 11851 27800
rect 11919 27744 11975 27800
rect 12043 27744 12099 27800
rect 12167 27744 12223 27800
rect 12291 27744 12347 27800
rect 12415 27744 12471 27800
rect 10679 27620 10735 27676
rect 10803 27620 10859 27676
rect 10927 27620 10983 27676
rect 11051 27620 11107 27676
rect 11175 27620 11231 27676
rect 11299 27620 11355 27676
rect 11423 27620 11479 27676
rect 11547 27620 11603 27676
rect 11671 27620 11727 27676
rect 11795 27620 11851 27676
rect 11919 27620 11975 27676
rect 12043 27620 12099 27676
rect 12167 27620 12223 27676
rect 12291 27620 12347 27676
rect 12415 27620 12471 27676
rect 10679 27496 10735 27552
rect 10803 27496 10859 27552
rect 10927 27496 10983 27552
rect 11051 27496 11107 27552
rect 11175 27496 11231 27552
rect 11299 27496 11355 27552
rect 11423 27496 11479 27552
rect 11547 27496 11603 27552
rect 11671 27496 11727 27552
rect 11795 27496 11851 27552
rect 11919 27496 11975 27552
rect 12043 27496 12099 27552
rect 12167 27496 12223 27552
rect 12291 27496 12347 27552
rect 12415 27496 12471 27552
rect 10679 27372 10735 27428
rect 10803 27372 10859 27428
rect 10927 27372 10983 27428
rect 11051 27372 11107 27428
rect 11175 27372 11231 27428
rect 11299 27372 11355 27428
rect 11423 27372 11479 27428
rect 11547 27372 11603 27428
rect 11671 27372 11727 27428
rect 11795 27372 11851 27428
rect 11919 27372 11975 27428
rect 12043 27372 12099 27428
rect 12167 27372 12223 27428
rect 12291 27372 12347 27428
rect 12415 27372 12471 27428
rect 10679 27248 10735 27304
rect 10803 27248 10859 27304
rect 10927 27248 10983 27304
rect 11051 27248 11107 27304
rect 11175 27248 11231 27304
rect 11299 27248 11355 27304
rect 11423 27248 11479 27304
rect 11547 27248 11603 27304
rect 11671 27248 11727 27304
rect 11795 27248 11851 27304
rect 11919 27248 11975 27304
rect 12043 27248 12099 27304
rect 12167 27248 12223 27304
rect 12291 27248 12347 27304
rect 12415 27248 12471 27304
rect 2507 26888 2563 26944
rect 2631 26888 2687 26944
rect 2755 26888 2811 26944
rect 2879 26888 2935 26944
rect 3003 26888 3059 26944
rect 3127 26888 3183 26944
rect 3251 26888 3307 26944
rect 3375 26888 3431 26944
rect 3499 26888 3555 26944
rect 3623 26888 3679 26944
rect 3747 26888 3803 26944
rect 3871 26888 3927 26944
rect 3995 26888 4051 26944
rect 4119 26888 4175 26944
rect 4243 26888 4299 26944
rect 2507 26764 2563 26820
rect 2631 26764 2687 26820
rect 2755 26764 2811 26820
rect 2879 26764 2935 26820
rect 3003 26764 3059 26820
rect 3127 26764 3183 26820
rect 3251 26764 3307 26820
rect 3375 26764 3431 26820
rect 3499 26764 3555 26820
rect 3623 26764 3679 26820
rect 3747 26764 3803 26820
rect 3871 26764 3927 26820
rect 3995 26764 4051 26820
rect 4119 26764 4175 26820
rect 4243 26764 4299 26820
rect 2507 26640 2563 26696
rect 2631 26640 2687 26696
rect 2755 26640 2811 26696
rect 2879 26640 2935 26696
rect 3003 26640 3059 26696
rect 3127 26640 3183 26696
rect 3251 26640 3307 26696
rect 3375 26640 3431 26696
rect 3499 26640 3555 26696
rect 3623 26640 3679 26696
rect 3747 26640 3803 26696
rect 3871 26640 3927 26696
rect 3995 26640 4051 26696
rect 4119 26640 4175 26696
rect 4243 26640 4299 26696
rect 2507 26516 2563 26572
rect 2631 26516 2687 26572
rect 2755 26516 2811 26572
rect 2879 26516 2935 26572
rect 3003 26516 3059 26572
rect 3127 26516 3183 26572
rect 3251 26516 3307 26572
rect 3375 26516 3431 26572
rect 3499 26516 3555 26572
rect 3623 26516 3679 26572
rect 3747 26516 3803 26572
rect 3871 26516 3927 26572
rect 3995 26516 4051 26572
rect 4119 26516 4175 26572
rect 4243 26516 4299 26572
rect 2507 26392 2563 26448
rect 2631 26392 2687 26448
rect 2755 26392 2811 26448
rect 2879 26392 2935 26448
rect 3003 26392 3059 26448
rect 3127 26392 3183 26448
rect 3251 26392 3307 26448
rect 3375 26392 3431 26448
rect 3499 26392 3555 26448
rect 3623 26392 3679 26448
rect 3747 26392 3803 26448
rect 3871 26392 3927 26448
rect 3995 26392 4051 26448
rect 4119 26392 4175 26448
rect 4243 26392 4299 26448
rect 2507 26268 2563 26324
rect 2631 26268 2687 26324
rect 2755 26268 2811 26324
rect 2879 26268 2935 26324
rect 3003 26268 3059 26324
rect 3127 26268 3183 26324
rect 3251 26268 3307 26324
rect 3375 26268 3431 26324
rect 3499 26268 3555 26324
rect 3623 26268 3679 26324
rect 3747 26268 3803 26324
rect 3871 26268 3927 26324
rect 3995 26268 4051 26324
rect 4119 26268 4175 26324
rect 4243 26268 4299 26324
rect 2507 26144 2563 26200
rect 2631 26144 2687 26200
rect 2755 26144 2811 26200
rect 2879 26144 2935 26200
rect 3003 26144 3059 26200
rect 3127 26144 3183 26200
rect 3251 26144 3307 26200
rect 3375 26144 3431 26200
rect 3499 26144 3555 26200
rect 3623 26144 3679 26200
rect 3747 26144 3803 26200
rect 3871 26144 3927 26200
rect 3995 26144 4051 26200
rect 4119 26144 4175 26200
rect 4243 26144 4299 26200
rect 2507 26020 2563 26076
rect 2631 26020 2687 26076
rect 2755 26020 2811 26076
rect 2879 26020 2935 26076
rect 3003 26020 3059 26076
rect 3127 26020 3183 26076
rect 3251 26020 3307 26076
rect 3375 26020 3431 26076
rect 3499 26020 3555 26076
rect 3623 26020 3679 26076
rect 3747 26020 3803 26076
rect 3871 26020 3927 26076
rect 3995 26020 4051 26076
rect 4119 26020 4175 26076
rect 4243 26020 4299 26076
rect 2507 25896 2563 25952
rect 2631 25896 2687 25952
rect 2755 25896 2811 25952
rect 2879 25896 2935 25952
rect 3003 25896 3059 25952
rect 3127 25896 3183 25952
rect 3251 25896 3307 25952
rect 3375 25896 3431 25952
rect 3499 25896 3555 25952
rect 3623 25896 3679 25952
rect 3747 25896 3803 25952
rect 3871 25896 3927 25952
rect 3995 25896 4051 25952
rect 4119 25896 4175 25952
rect 4243 25896 4299 25952
rect 2507 25772 2563 25828
rect 2631 25772 2687 25828
rect 2755 25772 2811 25828
rect 2879 25772 2935 25828
rect 3003 25772 3059 25828
rect 3127 25772 3183 25828
rect 3251 25772 3307 25828
rect 3375 25772 3431 25828
rect 3499 25772 3555 25828
rect 3623 25772 3679 25828
rect 3747 25772 3803 25828
rect 3871 25772 3927 25828
rect 3995 25772 4051 25828
rect 4119 25772 4175 25828
rect 4243 25772 4299 25828
rect 2507 25648 2563 25704
rect 2631 25648 2687 25704
rect 2755 25648 2811 25704
rect 2879 25648 2935 25704
rect 3003 25648 3059 25704
rect 3127 25648 3183 25704
rect 3251 25648 3307 25704
rect 3375 25648 3431 25704
rect 3499 25648 3555 25704
rect 3623 25648 3679 25704
rect 3747 25648 3803 25704
rect 3871 25648 3927 25704
rect 3995 25648 4051 25704
rect 4119 25648 4175 25704
rect 4243 25648 4299 25704
rect 6368 26888 6424 26944
rect 6492 26888 6548 26944
rect 6616 26888 6672 26944
rect 6740 26888 6796 26944
rect 6864 26888 6920 26944
rect 6988 26888 7044 26944
rect 7112 26888 7168 26944
rect 7236 26888 7292 26944
rect 7360 26888 7416 26944
rect 6368 26764 6424 26820
rect 6492 26764 6548 26820
rect 6616 26764 6672 26820
rect 6740 26764 6796 26820
rect 6864 26764 6920 26820
rect 6988 26764 7044 26820
rect 7112 26764 7168 26820
rect 7236 26764 7292 26820
rect 7360 26764 7416 26820
rect 6368 26640 6424 26696
rect 6492 26640 6548 26696
rect 6616 26640 6672 26696
rect 6740 26640 6796 26696
rect 6864 26640 6920 26696
rect 6988 26640 7044 26696
rect 7112 26640 7168 26696
rect 7236 26640 7292 26696
rect 7360 26640 7416 26696
rect 6368 26516 6424 26572
rect 6492 26516 6548 26572
rect 6616 26516 6672 26572
rect 6740 26516 6796 26572
rect 6864 26516 6920 26572
rect 6988 26516 7044 26572
rect 7112 26516 7168 26572
rect 7236 26516 7292 26572
rect 7360 26516 7416 26572
rect 6368 26392 6424 26448
rect 6492 26392 6548 26448
rect 6616 26392 6672 26448
rect 6740 26392 6796 26448
rect 6864 26392 6920 26448
rect 6988 26392 7044 26448
rect 7112 26392 7168 26448
rect 7236 26392 7292 26448
rect 7360 26392 7416 26448
rect 6368 26268 6424 26324
rect 6492 26268 6548 26324
rect 6616 26268 6672 26324
rect 6740 26268 6796 26324
rect 6864 26268 6920 26324
rect 6988 26268 7044 26324
rect 7112 26268 7168 26324
rect 7236 26268 7292 26324
rect 7360 26268 7416 26324
rect 6368 26144 6424 26200
rect 6492 26144 6548 26200
rect 6616 26144 6672 26200
rect 6740 26144 6796 26200
rect 6864 26144 6920 26200
rect 6988 26144 7044 26200
rect 7112 26144 7168 26200
rect 7236 26144 7292 26200
rect 7360 26144 7416 26200
rect 6368 26020 6424 26076
rect 6492 26020 6548 26076
rect 6616 26020 6672 26076
rect 6740 26020 6796 26076
rect 6864 26020 6920 26076
rect 6988 26020 7044 26076
rect 7112 26020 7168 26076
rect 7236 26020 7292 26076
rect 7360 26020 7416 26076
rect 6368 25896 6424 25952
rect 6492 25896 6548 25952
rect 6616 25896 6672 25952
rect 6740 25896 6796 25952
rect 6864 25896 6920 25952
rect 6988 25896 7044 25952
rect 7112 25896 7168 25952
rect 7236 25896 7292 25952
rect 7360 25896 7416 25952
rect 6368 25772 6424 25828
rect 6492 25772 6548 25828
rect 6616 25772 6672 25828
rect 6740 25772 6796 25828
rect 6864 25772 6920 25828
rect 6988 25772 7044 25828
rect 7112 25772 7168 25828
rect 7236 25772 7292 25828
rect 7360 25772 7416 25828
rect 6368 25648 6424 25704
rect 6492 25648 6548 25704
rect 6616 25648 6672 25704
rect 6740 25648 6796 25704
rect 6864 25648 6920 25704
rect 6988 25648 7044 25704
rect 7112 25648 7168 25704
rect 7236 25648 7292 25704
rect 7360 25648 7416 25704
rect 8751 26888 8807 26944
rect 8875 26888 8931 26944
rect 8999 26888 9055 26944
rect 9123 26888 9179 26944
rect 9247 26888 9303 26944
rect 9371 26888 9427 26944
rect 9495 26888 9551 26944
rect 9619 26888 9675 26944
rect 9743 26888 9799 26944
rect 9867 26888 9923 26944
rect 9991 26888 10047 26944
rect 10115 26888 10171 26944
rect 10239 26888 10295 26944
rect 10363 26888 10419 26944
rect 10487 26888 10543 26944
rect 8751 26764 8807 26820
rect 8875 26764 8931 26820
rect 8999 26764 9055 26820
rect 9123 26764 9179 26820
rect 9247 26764 9303 26820
rect 9371 26764 9427 26820
rect 9495 26764 9551 26820
rect 9619 26764 9675 26820
rect 9743 26764 9799 26820
rect 9867 26764 9923 26820
rect 9991 26764 10047 26820
rect 10115 26764 10171 26820
rect 10239 26764 10295 26820
rect 10363 26764 10419 26820
rect 10487 26764 10543 26820
rect 8751 26640 8807 26696
rect 8875 26640 8931 26696
rect 8999 26640 9055 26696
rect 9123 26640 9179 26696
rect 9247 26640 9303 26696
rect 9371 26640 9427 26696
rect 9495 26640 9551 26696
rect 9619 26640 9675 26696
rect 9743 26640 9799 26696
rect 9867 26640 9923 26696
rect 9991 26640 10047 26696
rect 10115 26640 10171 26696
rect 10239 26640 10295 26696
rect 10363 26640 10419 26696
rect 10487 26640 10543 26696
rect 8751 26516 8807 26572
rect 8875 26516 8931 26572
rect 8999 26516 9055 26572
rect 9123 26516 9179 26572
rect 9247 26516 9303 26572
rect 9371 26516 9427 26572
rect 9495 26516 9551 26572
rect 9619 26516 9675 26572
rect 9743 26516 9799 26572
rect 9867 26516 9923 26572
rect 9991 26516 10047 26572
rect 10115 26516 10171 26572
rect 10239 26516 10295 26572
rect 10363 26516 10419 26572
rect 10487 26516 10543 26572
rect 8751 26392 8807 26448
rect 8875 26392 8931 26448
rect 8999 26392 9055 26448
rect 9123 26392 9179 26448
rect 9247 26392 9303 26448
rect 9371 26392 9427 26448
rect 9495 26392 9551 26448
rect 9619 26392 9675 26448
rect 9743 26392 9799 26448
rect 9867 26392 9923 26448
rect 9991 26392 10047 26448
rect 10115 26392 10171 26448
rect 10239 26392 10295 26448
rect 10363 26392 10419 26448
rect 10487 26392 10543 26448
rect 8751 26268 8807 26324
rect 8875 26268 8931 26324
rect 8999 26268 9055 26324
rect 9123 26268 9179 26324
rect 9247 26268 9303 26324
rect 9371 26268 9427 26324
rect 9495 26268 9551 26324
rect 9619 26268 9675 26324
rect 9743 26268 9799 26324
rect 9867 26268 9923 26324
rect 9991 26268 10047 26324
rect 10115 26268 10171 26324
rect 10239 26268 10295 26324
rect 10363 26268 10419 26324
rect 10487 26268 10543 26324
rect 8751 26144 8807 26200
rect 8875 26144 8931 26200
rect 8999 26144 9055 26200
rect 9123 26144 9179 26200
rect 9247 26144 9303 26200
rect 9371 26144 9427 26200
rect 9495 26144 9551 26200
rect 9619 26144 9675 26200
rect 9743 26144 9799 26200
rect 9867 26144 9923 26200
rect 9991 26144 10047 26200
rect 10115 26144 10171 26200
rect 10239 26144 10295 26200
rect 10363 26144 10419 26200
rect 10487 26144 10543 26200
rect 8751 26020 8807 26076
rect 8875 26020 8931 26076
rect 8999 26020 9055 26076
rect 9123 26020 9179 26076
rect 9247 26020 9303 26076
rect 9371 26020 9427 26076
rect 9495 26020 9551 26076
rect 9619 26020 9675 26076
rect 9743 26020 9799 26076
rect 9867 26020 9923 26076
rect 9991 26020 10047 26076
rect 10115 26020 10171 26076
rect 10239 26020 10295 26076
rect 10363 26020 10419 26076
rect 10487 26020 10543 26076
rect 8751 25896 8807 25952
rect 8875 25896 8931 25952
rect 8999 25896 9055 25952
rect 9123 25896 9179 25952
rect 9247 25896 9303 25952
rect 9371 25896 9427 25952
rect 9495 25896 9551 25952
rect 9619 25896 9675 25952
rect 9743 25896 9799 25952
rect 9867 25896 9923 25952
rect 9991 25896 10047 25952
rect 10115 25896 10171 25952
rect 10239 25896 10295 25952
rect 10363 25896 10419 25952
rect 10487 25896 10543 25952
rect 8751 25772 8807 25828
rect 8875 25772 8931 25828
rect 8999 25772 9055 25828
rect 9123 25772 9179 25828
rect 9247 25772 9303 25828
rect 9371 25772 9427 25828
rect 9495 25772 9551 25828
rect 9619 25772 9675 25828
rect 9743 25772 9799 25828
rect 9867 25772 9923 25828
rect 9991 25772 10047 25828
rect 10115 25772 10171 25828
rect 10239 25772 10295 25828
rect 10363 25772 10419 25828
rect 10487 25772 10543 25828
rect 8751 25648 8807 25704
rect 8875 25648 8931 25704
rect 8999 25648 9055 25704
rect 9123 25648 9179 25704
rect 9247 25648 9303 25704
rect 9371 25648 9427 25704
rect 9495 25648 9551 25704
rect 9619 25648 9675 25704
rect 9743 25648 9799 25704
rect 9867 25648 9923 25704
rect 9991 25648 10047 25704
rect 10115 25648 10171 25704
rect 10239 25648 10295 25704
rect 10363 25648 10419 25704
rect 10487 25648 10543 25704
rect 12852 26888 12908 26944
rect 12976 26888 13032 26944
rect 13100 26888 13156 26944
rect 13224 26888 13280 26944
rect 13348 26888 13404 26944
rect 13472 26888 13528 26944
rect 13596 26888 13652 26944
rect 13720 26888 13776 26944
rect 13844 26888 13900 26944
rect 12852 26764 12908 26820
rect 12976 26764 13032 26820
rect 13100 26764 13156 26820
rect 13224 26764 13280 26820
rect 13348 26764 13404 26820
rect 13472 26764 13528 26820
rect 13596 26764 13652 26820
rect 13720 26764 13776 26820
rect 13844 26764 13900 26820
rect 12852 26640 12908 26696
rect 12976 26640 13032 26696
rect 13100 26640 13156 26696
rect 13224 26640 13280 26696
rect 13348 26640 13404 26696
rect 13472 26640 13528 26696
rect 13596 26640 13652 26696
rect 13720 26640 13776 26696
rect 13844 26640 13900 26696
rect 12852 26516 12908 26572
rect 12976 26516 13032 26572
rect 13100 26516 13156 26572
rect 13224 26516 13280 26572
rect 13348 26516 13404 26572
rect 13472 26516 13528 26572
rect 13596 26516 13652 26572
rect 13720 26516 13776 26572
rect 13844 26516 13900 26572
rect 12852 26392 12908 26448
rect 12976 26392 13032 26448
rect 13100 26392 13156 26448
rect 13224 26392 13280 26448
rect 13348 26392 13404 26448
rect 13472 26392 13528 26448
rect 13596 26392 13652 26448
rect 13720 26392 13776 26448
rect 13844 26392 13900 26448
rect 12852 26268 12908 26324
rect 12976 26268 13032 26324
rect 13100 26268 13156 26324
rect 13224 26268 13280 26324
rect 13348 26268 13404 26324
rect 13472 26268 13528 26324
rect 13596 26268 13652 26324
rect 13720 26268 13776 26324
rect 13844 26268 13900 26324
rect 12852 26144 12908 26200
rect 12976 26144 13032 26200
rect 13100 26144 13156 26200
rect 13224 26144 13280 26200
rect 13348 26144 13404 26200
rect 13472 26144 13528 26200
rect 13596 26144 13652 26200
rect 13720 26144 13776 26200
rect 13844 26144 13900 26200
rect 12852 26020 12908 26076
rect 12976 26020 13032 26076
rect 13100 26020 13156 26076
rect 13224 26020 13280 26076
rect 13348 26020 13404 26076
rect 13472 26020 13528 26076
rect 13596 26020 13652 26076
rect 13720 26020 13776 26076
rect 13844 26020 13900 26076
rect 12852 25896 12908 25952
rect 12976 25896 13032 25952
rect 13100 25896 13156 25952
rect 13224 25896 13280 25952
rect 13348 25896 13404 25952
rect 13472 25896 13528 25952
rect 13596 25896 13652 25952
rect 13720 25896 13776 25952
rect 13844 25896 13900 25952
rect 12852 25772 12908 25828
rect 12976 25772 13032 25828
rect 13100 25772 13156 25828
rect 13224 25772 13280 25828
rect 13348 25772 13404 25828
rect 13472 25772 13528 25828
rect 13596 25772 13652 25828
rect 13720 25772 13776 25828
rect 13844 25772 13900 25828
rect 12852 25648 12908 25704
rect 12976 25648 13032 25704
rect 13100 25648 13156 25704
rect 13224 25648 13280 25704
rect 13348 25648 13404 25704
rect 13472 25648 13528 25704
rect 13596 25648 13652 25704
rect 13720 25648 13776 25704
rect 13844 25648 13900 25704
rect 1078 25294 1134 25350
rect 1202 25294 1258 25350
rect 1326 25294 1382 25350
rect 1450 25294 1506 25350
rect 1574 25294 1630 25350
rect 1698 25294 1754 25350
rect 1822 25294 1878 25350
rect 1946 25294 2002 25350
rect 2070 25294 2126 25350
rect 1078 25170 1134 25226
rect 1202 25170 1258 25226
rect 1326 25170 1382 25226
rect 1450 25170 1506 25226
rect 1574 25170 1630 25226
rect 1698 25170 1754 25226
rect 1822 25170 1878 25226
rect 1946 25170 2002 25226
rect 2070 25170 2126 25226
rect 1078 25046 1134 25102
rect 1202 25046 1258 25102
rect 1326 25046 1382 25102
rect 1450 25046 1506 25102
rect 1574 25046 1630 25102
rect 1698 25046 1754 25102
rect 1822 25046 1878 25102
rect 1946 25046 2002 25102
rect 2070 25046 2126 25102
rect 1078 24922 1134 24978
rect 1202 24922 1258 24978
rect 1326 24922 1382 24978
rect 1450 24922 1506 24978
rect 1574 24922 1630 24978
rect 1698 24922 1754 24978
rect 1822 24922 1878 24978
rect 1946 24922 2002 24978
rect 2070 24922 2126 24978
rect 1078 24798 1134 24854
rect 1202 24798 1258 24854
rect 1326 24798 1382 24854
rect 1450 24798 1506 24854
rect 1574 24798 1630 24854
rect 1698 24798 1754 24854
rect 1822 24798 1878 24854
rect 1946 24798 2002 24854
rect 2070 24798 2126 24854
rect 1078 24674 1134 24730
rect 1202 24674 1258 24730
rect 1326 24674 1382 24730
rect 1450 24674 1506 24730
rect 1574 24674 1630 24730
rect 1698 24674 1754 24730
rect 1822 24674 1878 24730
rect 1946 24674 2002 24730
rect 2070 24674 2126 24730
rect 1078 24550 1134 24606
rect 1202 24550 1258 24606
rect 1326 24550 1382 24606
rect 1450 24550 1506 24606
rect 1574 24550 1630 24606
rect 1698 24550 1754 24606
rect 1822 24550 1878 24606
rect 1946 24550 2002 24606
rect 2070 24550 2126 24606
rect 1078 24426 1134 24482
rect 1202 24426 1258 24482
rect 1326 24426 1382 24482
rect 1450 24426 1506 24482
rect 1574 24426 1630 24482
rect 1698 24426 1754 24482
rect 1822 24426 1878 24482
rect 1946 24426 2002 24482
rect 2070 24426 2126 24482
rect 1078 24302 1134 24358
rect 1202 24302 1258 24358
rect 1326 24302 1382 24358
rect 1450 24302 1506 24358
rect 1574 24302 1630 24358
rect 1698 24302 1754 24358
rect 1822 24302 1878 24358
rect 1946 24302 2002 24358
rect 2070 24302 2126 24358
rect 1078 24178 1134 24234
rect 1202 24178 1258 24234
rect 1326 24178 1382 24234
rect 1450 24178 1506 24234
rect 1574 24178 1630 24234
rect 1698 24178 1754 24234
rect 1822 24178 1878 24234
rect 1946 24178 2002 24234
rect 2070 24178 2126 24234
rect 1078 24054 1134 24110
rect 1202 24054 1258 24110
rect 1326 24054 1382 24110
rect 1450 24054 1506 24110
rect 1574 24054 1630 24110
rect 1698 24054 1754 24110
rect 1822 24054 1878 24110
rect 1946 24054 2002 24110
rect 2070 24054 2126 24110
rect 1078 23930 1134 23986
rect 1202 23930 1258 23986
rect 1326 23930 1382 23986
rect 1450 23930 1506 23986
rect 1574 23930 1630 23986
rect 1698 23930 1754 23986
rect 1822 23930 1878 23986
rect 1946 23930 2002 23986
rect 2070 23930 2126 23986
rect 1078 23806 1134 23862
rect 1202 23806 1258 23862
rect 1326 23806 1382 23862
rect 1450 23806 1506 23862
rect 1574 23806 1630 23862
rect 1698 23806 1754 23862
rect 1822 23806 1878 23862
rect 1946 23806 2002 23862
rect 2070 23806 2126 23862
rect 1078 23682 1134 23738
rect 1202 23682 1258 23738
rect 1326 23682 1382 23738
rect 1450 23682 1506 23738
rect 1574 23682 1630 23738
rect 1698 23682 1754 23738
rect 1822 23682 1878 23738
rect 1946 23682 2002 23738
rect 2070 23682 2126 23738
rect 1078 23558 1134 23614
rect 1202 23558 1258 23614
rect 1326 23558 1382 23614
rect 1450 23558 1506 23614
rect 1574 23558 1630 23614
rect 1698 23558 1754 23614
rect 1822 23558 1878 23614
rect 1946 23558 2002 23614
rect 2070 23558 2126 23614
rect 1078 23434 1134 23490
rect 1202 23434 1258 23490
rect 1326 23434 1382 23490
rect 1450 23434 1506 23490
rect 1574 23434 1630 23490
rect 1698 23434 1754 23490
rect 1822 23434 1878 23490
rect 1946 23434 2002 23490
rect 2070 23434 2126 23490
rect 1078 23310 1134 23366
rect 1202 23310 1258 23366
rect 1326 23310 1382 23366
rect 1450 23310 1506 23366
rect 1574 23310 1630 23366
rect 1698 23310 1754 23366
rect 1822 23310 1878 23366
rect 1946 23310 2002 23366
rect 2070 23310 2126 23366
rect 1078 23186 1134 23242
rect 1202 23186 1258 23242
rect 1326 23186 1382 23242
rect 1450 23186 1506 23242
rect 1574 23186 1630 23242
rect 1698 23186 1754 23242
rect 1822 23186 1878 23242
rect 1946 23186 2002 23242
rect 2070 23186 2126 23242
rect 1078 23062 1134 23118
rect 1202 23062 1258 23118
rect 1326 23062 1382 23118
rect 1450 23062 1506 23118
rect 1574 23062 1630 23118
rect 1698 23062 1754 23118
rect 1822 23062 1878 23118
rect 1946 23062 2002 23118
rect 2070 23062 2126 23118
rect 1078 22938 1134 22994
rect 1202 22938 1258 22994
rect 1326 22938 1382 22994
rect 1450 22938 1506 22994
rect 1574 22938 1630 22994
rect 1698 22938 1754 22994
rect 1822 22938 1878 22994
rect 1946 22938 2002 22994
rect 2070 22938 2126 22994
rect 1078 22814 1134 22870
rect 1202 22814 1258 22870
rect 1326 22814 1382 22870
rect 1450 22814 1506 22870
rect 1574 22814 1630 22870
rect 1698 22814 1754 22870
rect 1822 22814 1878 22870
rect 1946 22814 2002 22870
rect 2070 22814 2126 22870
rect 1078 22690 1134 22746
rect 1202 22690 1258 22746
rect 1326 22690 1382 22746
rect 1450 22690 1506 22746
rect 1574 22690 1630 22746
rect 1698 22690 1754 22746
rect 1822 22690 1878 22746
rect 1946 22690 2002 22746
rect 2070 22690 2126 22746
rect 1078 22566 1134 22622
rect 1202 22566 1258 22622
rect 1326 22566 1382 22622
rect 1450 22566 1506 22622
rect 1574 22566 1630 22622
rect 1698 22566 1754 22622
rect 1822 22566 1878 22622
rect 1946 22566 2002 22622
rect 2070 22566 2126 22622
rect 1078 22442 1134 22498
rect 1202 22442 1258 22498
rect 1326 22442 1382 22498
rect 1450 22442 1506 22498
rect 1574 22442 1630 22498
rect 1698 22442 1754 22498
rect 1822 22442 1878 22498
rect 1946 22442 2002 22498
rect 2070 22442 2126 22498
rect 4435 25294 4491 25350
rect 4559 25294 4615 25350
rect 4683 25294 4739 25350
rect 4807 25294 4863 25350
rect 4931 25294 4987 25350
rect 5055 25294 5111 25350
rect 5179 25294 5235 25350
rect 5303 25294 5359 25350
rect 5427 25294 5483 25350
rect 5551 25294 5607 25350
rect 5675 25294 5731 25350
rect 5799 25294 5855 25350
rect 5923 25294 5979 25350
rect 6047 25294 6103 25350
rect 6171 25294 6227 25350
rect 4435 25170 4491 25226
rect 4559 25170 4615 25226
rect 4683 25170 4739 25226
rect 4807 25170 4863 25226
rect 4931 25170 4987 25226
rect 5055 25170 5111 25226
rect 5179 25170 5235 25226
rect 5303 25170 5359 25226
rect 5427 25170 5483 25226
rect 5551 25170 5607 25226
rect 5675 25170 5731 25226
rect 5799 25170 5855 25226
rect 5923 25170 5979 25226
rect 6047 25170 6103 25226
rect 6171 25170 6227 25226
rect 4435 25046 4491 25102
rect 4559 25046 4615 25102
rect 4683 25046 4739 25102
rect 4807 25046 4863 25102
rect 4931 25046 4987 25102
rect 5055 25046 5111 25102
rect 5179 25046 5235 25102
rect 5303 25046 5359 25102
rect 5427 25046 5483 25102
rect 5551 25046 5607 25102
rect 5675 25046 5731 25102
rect 5799 25046 5855 25102
rect 5923 25046 5979 25102
rect 6047 25046 6103 25102
rect 6171 25046 6227 25102
rect 4435 24922 4491 24978
rect 4559 24922 4615 24978
rect 4683 24922 4739 24978
rect 4807 24922 4863 24978
rect 4931 24922 4987 24978
rect 5055 24922 5111 24978
rect 5179 24922 5235 24978
rect 5303 24922 5359 24978
rect 5427 24922 5483 24978
rect 5551 24922 5607 24978
rect 5675 24922 5731 24978
rect 5799 24922 5855 24978
rect 5923 24922 5979 24978
rect 6047 24922 6103 24978
rect 6171 24922 6227 24978
rect 4435 24798 4491 24854
rect 4559 24798 4615 24854
rect 4683 24798 4739 24854
rect 4807 24798 4863 24854
rect 4931 24798 4987 24854
rect 5055 24798 5111 24854
rect 5179 24798 5235 24854
rect 5303 24798 5359 24854
rect 5427 24798 5483 24854
rect 5551 24798 5607 24854
rect 5675 24798 5731 24854
rect 5799 24798 5855 24854
rect 5923 24798 5979 24854
rect 6047 24798 6103 24854
rect 6171 24798 6227 24854
rect 4435 24674 4491 24730
rect 4559 24674 4615 24730
rect 4683 24674 4739 24730
rect 4807 24674 4863 24730
rect 4931 24674 4987 24730
rect 5055 24674 5111 24730
rect 5179 24674 5235 24730
rect 5303 24674 5359 24730
rect 5427 24674 5483 24730
rect 5551 24674 5607 24730
rect 5675 24674 5731 24730
rect 5799 24674 5855 24730
rect 5923 24674 5979 24730
rect 6047 24674 6103 24730
rect 6171 24674 6227 24730
rect 4435 24550 4491 24606
rect 4559 24550 4615 24606
rect 4683 24550 4739 24606
rect 4807 24550 4863 24606
rect 4931 24550 4987 24606
rect 5055 24550 5111 24606
rect 5179 24550 5235 24606
rect 5303 24550 5359 24606
rect 5427 24550 5483 24606
rect 5551 24550 5607 24606
rect 5675 24550 5731 24606
rect 5799 24550 5855 24606
rect 5923 24550 5979 24606
rect 6047 24550 6103 24606
rect 6171 24550 6227 24606
rect 4435 24426 4491 24482
rect 4559 24426 4615 24482
rect 4683 24426 4739 24482
rect 4807 24426 4863 24482
rect 4931 24426 4987 24482
rect 5055 24426 5111 24482
rect 5179 24426 5235 24482
rect 5303 24426 5359 24482
rect 5427 24426 5483 24482
rect 5551 24426 5607 24482
rect 5675 24426 5731 24482
rect 5799 24426 5855 24482
rect 5923 24426 5979 24482
rect 6047 24426 6103 24482
rect 6171 24426 6227 24482
rect 4435 24302 4491 24358
rect 4559 24302 4615 24358
rect 4683 24302 4739 24358
rect 4807 24302 4863 24358
rect 4931 24302 4987 24358
rect 5055 24302 5111 24358
rect 5179 24302 5235 24358
rect 5303 24302 5359 24358
rect 5427 24302 5483 24358
rect 5551 24302 5607 24358
rect 5675 24302 5731 24358
rect 5799 24302 5855 24358
rect 5923 24302 5979 24358
rect 6047 24302 6103 24358
rect 6171 24302 6227 24358
rect 4435 24178 4491 24234
rect 4559 24178 4615 24234
rect 4683 24178 4739 24234
rect 4807 24178 4863 24234
rect 4931 24178 4987 24234
rect 5055 24178 5111 24234
rect 5179 24178 5235 24234
rect 5303 24178 5359 24234
rect 5427 24178 5483 24234
rect 5551 24178 5607 24234
rect 5675 24178 5731 24234
rect 5799 24178 5855 24234
rect 5923 24178 5979 24234
rect 6047 24178 6103 24234
rect 6171 24178 6227 24234
rect 4435 24054 4491 24110
rect 4559 24054 4615 24110
rect 4683 24054 4739 24110
rect 4807 24054 4863 24110
rect 4931 24054 4987 24110
rect 5055 24054 5111 24110
rect 5179 24054 5235 24110
rect 5303 24054 5359 24110
rect 5427 24054 5483 24110
rect 5551 24054 5607 24110
rect 5675 24054 5731 24110
rect 5799 24054 5855 24110
rect 5923 24054 5979 24110
rect 6047 24054 6103 24110
rect 6171 24054 6227 24110
rect 4435 23930 4491 23986
rect 4559 23930 4615 23986
rect 4683 23930 4739 23986
rect 4807 23930 4863 23986
rect 4931 23930 4987 23986
rect 5055 23930 5111 23986
rect 5179 23930 5235 23986
rect 5303 23930 5359 23986
rect 5427 23930 5483 23986
rect 5551 23930 5607 23986
rect 5675 23930 5731 23986
rect 5799 23930 5855 23986
rect 5923 23930 5979 23986
rect 6047 23930 6103 23986
rect 6171 23930 6227 23986
rect 4435 23806 4491 23862
rect 4559 23806 4615 23862
rect 4683 23806 4739 23862
rect 4807 23806 4863 23862
rect 4931 23806 4987 23862
rect 5055 23806 5111 23862
rect 5179 23806 5235 23862
rect 5303 23806 5359 23862
rect 5427 23806 5483 23862
rect 5551 23806 5607 23862
rect 5675 23806 5731 23862
rect 5799 23806 5855 23862
rect 5923 23806 5979 23862
rect 6047 23806 6103 23862
rect 6171 23806 6227 23862
rect 4435 23682 4491 23738
rect 4559 23682 4615 23738
rect 4683 23682 4739 23738
rect 4807 23682 4863 23738
rect 4931 23682 4987 23738
rect 5055 23682 5111 23738
rect 5179 23682 5235 23738
rect 5303 23682 5359 23738
rect 5427 23682 5483 23738
rect 5551 23682 5607 23738
rect 5675 23682 5731 23738
rect 5799 23682 5855 23738
rect 5923 23682 5979 23738
rect 6047 23682 6103 23738
rect 6171 23682 6227 23738
rect 4435 23558 4491 23614
rect 4559 23558 4615 23614
rect 4683 23558 4739 23614
rect 4807 23558 4863 23614
rect 4931 23558 4987 23614
rect 5055 23558 5111 23614
rect 5179 23558 5235 23614
rect 5303 23558 5359 23614
rect 5427 23558 5483 23614
rect 5551 23558 5607 23614
rect 5675 23558 5731 23614
rect 5799 23558 5855 23614
rect 5923 23558 5979 23614
rect 6047 23558 6103 23614
rect 6171 23558 6227 23614
rect 4435 23434 4491 23490
rect 4559 23434 4615 23490
rect 4683 23434 4739 23490
rect 4807 23434 4863 23490
rect 4931 23434 4987 23490
rect 5055 23434 5111 23490
rect 5179 23434 5235 23490
rect 5303 23434 5359 23490
rect 5427 23434 5483 23490
rect 5551 23434 5607 23490
rect 5675 23434 5731 23490
rect 5799 23434 5855 23490
rect 5923 23434 5979 23490
rect 6047 23434 6103 23490
rect 6171 23434 6227 23490
rect 4435 23310 4491 23366
rect 4559 23310 4615 23366
rect 4683 23310 4739 23366
rect 4807 23310 4863 23366
rect 4931 23310 4987 23366
rect 5055 23310 5111 23366
rect 5179 23310 5235 23366
rect 5303 23310 5359 23366
rect 5427 23310 5483 23366
rect 5551 23310 5607 23366
rect 5675 23310 5731 23366
rect 5799 23310 5855 23366
rect 5923 23310 5979 23366
rect 6047 23310 6103 23366
rect 6171 23310 6227 23366
rect 4435 23186 4491 23242
rect 4559 23186 4615 23242
rect 4683 23186 4739 23242
rect 4807 23186 4863 23242
rect 4931 23186 4987 23242
rect 5055 23186 5111 23242
rect 5179 23186 5235 23242
rect 5303 23186 5359 23242
rect 5427 23186 5483 23242
rect 5551 23186 5607 23242
rect 5675 23186 5731 23242
rect 5799 23186 5855 23242
rect 5923 23186 5979 23242
rect 6047 23186 6103 23242
rect 6171 23186 6227 23242
rect 4435 23062 4491 23118
rect 4559 23062 4615 23118
rect 4683 23062 4739 23118
rect 4807 23062 4863 23118
rect 4931 23062 4987 23118
rect 5055 23062 5111 23118
rect 5179 23062 5235 23118
rect 5303 23062 5359 23118
rect 5427 23062 5483 23118
rect 5551 23062 5607 23118
rect 5675 23062 5731 23118
rect 5799 23062 5855 23118
rect 5923 23062 5979 23118
rect 6047 23062 6103 23118
rect 6171 23062 6227 23118
rect 4435 22938 4491 22994
rect 4559 22938 4615 22994
rect 4683 22938 4739 22994
rect 4807 22938 4863 22994
rect 4931 22938 4987 22994
rect 5055 22938 5111 22994
rect 5179 22938 5235 22994
rect 5303 22938 5359 22994
rect 5427 22938 5483 22994
rect 5551 22938 5607 22994
rect 5675 22938 5731 22994
rect 5799 22938 5855 22994
rect 5923 22938 5979 22994
rect 6047 22938 6103 22994
rect 6171 22938 6227 22994
rect 4435 22814 4491 22870
rect 4559 22814 4615 22870
rect 4683 22814 4739 22870
rect 4807 22814 4863 22870
rect 4931 22814 4987 22870
rect 5055 22814 5111 22870
rect 5179 22814 5235 22870
rect 5303 22814 5359 22870
rect 5427 22814 5483 22870
rect 5551 22814 5607 22870
rect 5675 22814 5731 22870
rect 5799 22814 5855 22870
rect 5923 22814 5979 22870
rect 6047 22814 6103 22870
rect 6171 22814 6227 22870
rect 4435 22690 4491 22746
rect 4559 22690 4615 22746
rect 4683 22690 4739 22746
rect 4807 22690 4863 22746
rect 4931 22690 4987 22746
rect 5055 22690 5111 22746
rect 5179 22690 5235 22746
rect 5303 22690 5359 22746
rect 5427 22690 5483 22746
rect 5551 22690 5607 22746
rect 5675 22690 5731 22746
rect 5799 22690 5855 22746
rect 5923 22690 5979 22746
rect 6047 22690 6103 22746
rect 6171 22690 6227 22746
rect 4435 22566 4491 22622
rect 4559 22566 4615 22622
rect 4683 22566 4739 22622
rect 4807 22566 4863 22622
rect 4931 22566 4987 22622
rect 5055 22566 5111 22622
rect 5179 22566 5235 22622
rect 5303 22566 5359 22622
rect 5427 22566 5483 22622
rect 5551 22566 5607 22622
rect 5675 22566 5731 22622
rect 5799 22566 5855 22622
rect 5923 22566 5979 22622
rect 6047 22566 6103 22622
rect 6171 22566 6227 22622
rect 4435 22442 4491 22498
rect 4559 22442 4615 22498
rect 4683 22442 4739 22498
rect 4807 22442 4863 22498
rect 4931 22442 4987 22498
rect 5055 22442 5111 22498
rect 5179 22442 5235 22498
rect 5303 22442 5359 22498
rect 5427 22442 5483 22498
rect 5551 22442 5607 22498
rect 5675 22442 5731 22498
rect 5799 22442 5855 22498
rect 5923 22442 5979 22498
rect 6047 22442 6103 22498
rect 6171 22442 6227 22498
rect 7562 25294 7618 25350
rect 7686 25294 7742 25350
rect 7810 25294 7866 25350
rect 7934 25294 7990 25350
rect 8058 25294 8114 25350
rect 8182 25294 8238 25350
rect 8306 25294 8362 25350
rect 8430 25294 8486 25350
rect 8554 25294 8610 25350
rect 7562 25170 7618 25226
rect 7686 25170 7742 25226
rect 7810 25170 7866 25226
rect 7934 25170 7990 25226
rect 8058 25170 8114 25226
rect 8182 25170 8238 25226
rect 8306 25170 8362 25226
rect 8430 25170 8486 25226
rect 8554 25170 8610 25226
rect 7562 25046 7618 25102
rect 7686 25046 7742 25102
rect 7810 25046 7866 25102
rect 7934 25046 7990 25102
rect 8058 25046 8114 25102
rect 8182 25046 8238 25102
rect 8306 25046 8362 25102
rect 8430 25046 8486 25102
rect 8554 25046 8610 25102
rect 7562 24922 7618 24978
rect 7686 24922 7742 24978
rect 7810 24922 7866 24978
rect 7934 24922 7990 24978
rect 8058 24922 8114 24978
rect 8182 24922 8238 24978
rect 8306 24922 8362 24978
rect 8430 24922 8486 24978
rect 8554 24922 8610 24978
rect 7562 24798 7618 24854
rect 7686 24798 7742 24854
rect 7810 24798 7866 24854
rect 7934 24798 7990 24854
rect 8058 24798 8114 24854
rect 8182 24798 8238 24854
rect 8306 24798 8362 24854
rect 8430 24798 8486 24854
rect 8554 24798 8610 24854
rect 7562 24674 7618 24730
rect 7686 24674 7742 24730
rect 7810 24674 7866 24730
rect 7934 24674 7990 24730
rect 8058 24674 8114 24730
rect 8182 24674 8238 24730
rect 8306 24674 8362 24730
rect 8430 24674 8486 24730
rect 8554 24674 8610 24730
rect 7562 24550 7618 24606
rect 7686 24550 7742 24606
rect 7810 24550 7866 24606
rect 7934 24550 7990 24606
rect 8058 24550 8114 24606
rect 8182 24550 8238 24606
rect 8306 24550 8362 24606
rect 8430 24550 8486 24606
rect 8554 24550 8610 24606
rect 7562 24426 7618 24482
rect 7686 24426 7742 24482
rect 7810 24426 7866 24482
rect 7934 24426 7990 24482
rect 8058 24426 8114 24482
rect 8182 24426 8238 24482
rect 8306 24426 8362 24482
rect 8430 24426 8486 24482
rect 8554 24426 8610 24482
rect 7562 24302 7618 24358
rect 7686 24302 7742 24358
rect 7810 24302 7866 24358
rect 7934 24302 7990 24358
rect 8058 24302 8114 24358
rect 8182 24302 8238 24358
rect 8306 24302 8362 24358
rect 8430 24302 8486 24358
rect 8554 24302 8610 24358
rect 7562 24178 7618 24234
rect 7686 24178 7742 24234
rect 7810 24178 7866 24234
rect 7934 24178 7990 24234
rect 8058 24178 8114 24234
rect 8182 24178 8238 24234
rect 8306 24178 8362 24234
rect 8430 24178 8486 24234
rect 8554 24178 8610 24234
rect 7562 24054 7618 24110
rect 7686 24054 7742 24110
rect 7810 24054 7866 24110
rect 7934 24054 7990 24110
rect 8058 24054 8114 24110
rect 8182 24054 8238 24110
rect 8306 24054 8362 24110
rect 8430 24054 8486 24110
rect 8554 24054 8610 24110
rect 7562 23930 7618 23986
rect 7686 23930 7742 23986
rect 7810 23930 7866 23986
rect 7934 23930 7990 23986
rect 8058 23930 8114 23986
rect 8182 23930 8238 23986
rect 8306 23930 8362 23986
rect 8430 23930 8486 23986
rect 8554 23930 8610 23986
rect 7562 23806 7618 23862
rect 7686 23806 7742 23862
rect 7810 23806 7866 23862
rect 7934 23806 7990 23862
rect 8058 23806 8114 23862
rect 8182 23806 8238 23862
rect 8306 23806 8362 23862
rect 8430 23806 8486 23862
rect 8554 23806 8610 23862
rect 7562 23682 7618 23738
rect 7686 23682 7742 23738
rect 7810 23682 7866 23738
rect 7934 23682 7990 23738
rect 8058 23682 8114 23738
rect 8182 23682 8238 23738
rect 8306 23682 8362 23738
rect 8430 23682 8486 23738
rect 8554 23682 8610 23738
rect 7562 23558 7618 23614
rect 7686 23558 7742 23614
rect 7810 23558 7866 23614
rect 7934 23558 7990 23614
rect 8058 23558 8114 23614
rect 8182 23558 8238 23614
rect 8306 23558 8362 23614
rect 8430 23558 8486 23614
rect 8554 23558 8610 23614
rect 7562 23434 7618 23490
rect 7686 23434 7742 23490
rect 7810 23434 7866 23490
rect 7934 23434 7990 23490
rect 8058 23434 8114 23490
rect 8182 23434 8238 23490
rect 8306 23434 8362 23490
rect 8430 23434 8486 23490
rect 8554 23434 8610 23490
rect 7562 23310 7618 23366
rect 7686 23310 7742 23366
rect 7810 23310 7866 23366
rect 7934 23310 7990 23366
rect 8058 23310 8114 23366
rect 8182 23310 8238 23366
rect 8306 23310 8362 23366
rect 8430 23310 8486 23366
rect 8554 23310 8610 23366
rect 7562 23186 7618 23242
rect 7686 23186 7742 23242
rect 7810 23186 7866 23242
rect 7934 23186 7990 23242
rect 8058 23186 8114 23242
rect 8182 23186 8238 23242
rect 8306 23186 8362 23242
rect 8430 23186 8486 23242
rect 8554 23186 8610 23242
rect 7562 23062 7618 23118
rect 7686 23062 7742 23118
rect 7810 23062 7866 23118
rect 7934 23062 7990 23118
rect 8058 23062 8114 23118
rect 8182 23062 8238 23118
rect 8306 23062 8362 23118
rect 8430 23062 8486 23118
rect 8554 23062 8610 23118
rect 7562 22938 7618 22994
rect 7686 22938 7742 22994
rect 7810 22938 7866 22994
rect 7934 22938 7990 22994
rect 8058 22938 8114 22994
rect 8182 22938 8238 22994
rect 8306 22938 8362 22994
rect 8430 22938 8486 22994
rect 8554 22938 8610 22994
rect 7562 22814 7618 22870
rect 7686 22814 7742 22870
rect 7810 22814 7866 22870
rect 7934 22814 7990 22870
rect 8058 22814 8114 22870
rect 8182 22814 8238 22870
rect 8306 22814 8362 22870
rect 8430 22814 8486 22870
rect 8554 22814 8610 22870
rect 7562 22690 7618 22746
rect 7686 22690 7742 22746
rect 7810 22690 7866 22746
rect 7934 22690 7990 22746
rect 8058 22690 8114 22746
rect 8182 22690 8238 22746
rect 8306 22690 8362 22746
rect 8430 22690 8486 22746
rect 8554 22690 8610 22746
rect 7562 22566 7618 22622
rect 7686 22566 7742 22622
rect 7810 22566 7866 22622
rect 7934 22566 7990 22622
rect 8058 22566 8114 22622
rect 8182 22566 8238 22622
rect 8306 22566 8362 22622
rect 8430 22566 8486 22622
rect 8554 22566 8610 22622
rect 7562 22442 7618 22498
rect 7686 22442 7742 22498
rect 7810 22442 7866 22498
rect 7934 22442 7990 22498
rect 8058 22442 8114 22498
rect 8182 22442 8238 22498
rect 8306 22442 8362 22498
rect 8430 22442 8486 22498
rect 8554 22442 8610 22498
rect 10679 25294 10735 25350
rect 10803 25294 10859 25350
rect 10927 25294 10983 25350
rect 11051 25294 11107 25350
rect 11175 25294 11231 25350
rect 11299 25294 11355 25350
rect 11423 25294 11479 25350
rect 11547 25294 11603 25350
rect 11671 25294 11727 25350
rect 11795 25294 11851 25350
rect 11919 25294 11975 25350
rect 12043 25294 12099 25350
rect 12167 25294 12223 25350
rect 12291 25294 12347 25350
rect 12415 25294 12471 25350
rect 10679 25170 10735 25226
rect 10803 25170 10859 25226
rect 10927 25170 10983 25226
rect 11051 25170 11107 25226
rect 11175 25170 11231 25226
rect 11299 25170 11355 25226
rect 11423 25170 11479 25226
rect 11547 25170 11603 25226
rect 11671 25170 11727 25226
rect 11795 25170 11851 25226
rect 11919 25170 11975 25226
rect 12043 25170 12099 25226
rect 12167 25170 12223 25226
rect 12291 25170 12347 25226
rect 12415 25170 12471 25226
rect 10679 25046 10735 25102
rect 10803 25046 10859 25102
rect 10927 25046 10983 25102
rect 11051 25046 11107 25102
rect 11175 25046 11231 25102
rect 11299 25046 11355 25102
rect 11423 25046 11479 25102
rect 11547 25046 11603 25102
rect 11671 25046 11727 25102
rect 11795 25046 11851 25102
rect 11919 25046 11975 25102
rect 12043 25046 12099 25102
rect 12167 25046 12223 25102
rect 12291 25046 12347 25102
rect 12415 25046 12471 25102
rect 10679 24922 10735 24978
rect 10803 24922 10859 24978
rect 10927 24922 10983 24978
rect 11051 24922 11107 24978
rect 11175 24922 11231 24978
rect 11299 24922 11355 24978
rect 11423 24922 11479 24978
rect 11547 24922 11603 24978
rect 11671 24922 11727 24978
rect 11795 24922 11851 24978
rect 11919 24922 11975 24978
rect 12043 24922 12099 24978
rect 12167 24922 12223 24978
rect 12291 24922 12347 24978
rect 12415 24922 12471 24978
rect 10679 24798 10735 24854
rect 10803 24798 10859 24854
rect 10927 24798 10983 24854
rect 11051 24798 11107 24854
rect 11175 24798 11231 24854
rect 11299 24798 11355 24854
rect 11423 24798 11479 24854
rect 11547 24798 11603 24854
rect 11671 24798 11727 24854
rect 11795 24798 11851 24854
rect 11919 24798 11975 24854
rect 12043 24798 12099 24854
rect 12167 24798 12223 24854
rect 12291 24798 12347 24854
rect 12415 24798 12471 24854
rect 10679 24674 10735 24730
rect 10803 24674 10859 24730
rect 10927 24674 10983 24730
rect 11051 24674 11107 24730
rect 11175 24674 11231 24730
rect 11299 24674 11355 24730
rect 11423 24674 11479 24730
rect 11547 24674 11603 24730
rect 11671 24674 11727 24730
rect 11795 24674 11851 24730
rect 11919 24674 11975 24730
rect 12043 24674 12099 24730
rect 12167 24674 12223 24730
rect 12291 24674 12347 24730
rect 12415 24674 12471 24730
rect 10679 24550 10735 24606
rect 10803 24550 10859 24606
rect 10927 24550 10983 24606
rect 11051 24550 11107 24606
rect 11175 24550 11231 24606
rect 11299 24550 11355 24606
rect 11423 24550 11479 24606
rect 11547 24550 11603 24606
rect 11671 24550 11727 24606
rect 11795 24550 11851 24606
rect 11919 24550 11975 24606
rect 12043 24550 12099 24606
rect 12167 24550 12223 24606
rect 12291 24550 12347 24606
rect 12415 24550 12471 24606
rect 10679 24426 10735 24482
rect 10803 24426 10859 24482
rect 10927 24426 10983 24482
rect 11051 24426 11107 24482
rect 11175 24426 11231 24482
rect 11299 24426 11355 24482
rect 11423 24426 11479 24482
rect 11547 24426 11603 24482
rect 11671 24426 11727 24482
rect 11795 24426 11851 24482
rect 11919 24426 11975 24482
rect 12043 24426 12099 24482
rect 12167 24426 12223 24482
rect 12291 24426 12347 24482
rect 12415 24426 12471 24482
rect 10679 24302 10735 24358
rect 10803 24302 10859 24358
rect 10927 24302 10983 24358
rect 11051 24302 11107 24358
rect 11175 24302 11231 24358
rect 11299 24302 11355 24358
rect 11423 24302 11479 24358
rect 11547 24302 11603 24358
rect 11671 24302 11727 24358
rect 11795 24302 11851 24358
rect 11919 24302 11975 24358
rect 12043 24302 12099 24358
rect 12167 24302 12223 24358
rect 12291 24302 12347 24358
rect 12415 24302 12471 24358
rect 10679 24178 10735 24234
rect 10803 24178 10859 24234
rect 10927 24178 10983 24234
rect 11051 24178 11107 24234
rect 11175 24178 11231 24234
rect 11299 24178 11355 24234
rect 11423 24178 11479 24234
rect 11547 24178 11603 24234
rect 11671 24178 11727 24234
rect 11795 24178 11851 24234
rect 11919 24178 11975 24234
rect 12043 24178 12099 24234
rect 12167 24178 12223 24234
rect 12291 24178 12347 24234
rect 12415 24178 12471 24234
rect 10679 24054 10735 24110
rect 10803 24054 10859 24110
rect 10927 24054 10983 24110
rect 11051 24054 11107 24110
rect 11175 24054 11231 24110
rect 11299 24054 11355 24110
rect 11423 24054 11479 24110
rect 11547 24054 11603 24110
rect 11671 24054 11727 24110
rect 11795 24054 11851 24110
rect 11919 24054 11975 24110
rect 12043 24054 12099 24110
rect 12167 24054 12223 24110
rect 12291 24054 12347 24110
rect 12415 24054 12471 24110
rect 10679 23930 10735 23986
rect 10803 23930 10859 23986
rect 10927 23930 10983 23986
rect 11051 23930 11107 23986
rect 11175 23930 11231 23986
rect 11299 23930 11355 23986
rect 11423 23930 11479 23986
rect 11547 23930 11603 23986
rect 11671 23930 11727 23986
rect 11795 23930 11851 23986
rect 11919 23930 11975 23986
rect 12043 23930 12099 23986
rect 12167 23930 12223 23986
rect 12291 23930 12347 23986
rect 12415 23930 12471 23986
rect 10679 23806 10735 23862
rect 10803 23806 10859 23862
rect 10927 23806 10983 23862
rect 11051 23806 11107 23862
rect 11175 23806 11231 23862
rect 11299 23806 11355 23862
rect 11423 23806 11479 23862
rect 11547 23806 11603 23862
rect 11671 23806 11727 23862
rect 11795 23806 11851 23862
rect 11919 23806 11975 23862
rect 12043 23806 12099 23862
rect 12167 23806 12223 23862
rect 12291 23806 12347 23862
rect 12415 23806 12471 23862
rect 10679 23682 10735 23738
rect 10803 23682 10859 23738
rect 10927 23682 10983 23738
rect 11051 23682 11107 23738
rect 11175 23682 11231 23738
rect 11299 23682 11355 23738
rect 11423 23682 11479 23738
rect 11547 23682 11603 23738
rect 11671 23682 11727 23738
rect 11795 23682 11851 23738
rect 11919 23682 11975 23738
rect 12043 23682 12099 23738
rect 12167 23682 12223 23738
rect 12291 23682 12347 23738
rect 12415 23682 12471 23738
rect 10679 23558 10735 23614
rect 10803 23558 10859 23614
rect 10927 23558 10983 23614
rect 11051 23558 11107 23614
rect 11175 23558 11231 23614
rect 11299 23558 11355 23614
rect 11423 23558 11479 23614
rect 11547 23558 11603 23614
rect 11671 23558 11727 23614
rect 11795 23558 11851 23614
rect 11919 23558 11975 23614
rect 12043 23558 12099 23614
rect 12167 23558 12223 23614
rect 12291 23558 12347 23614
rect 12415 23558 12471 23614
rect 10679 23434 10735 23490
rect 10803 23434 10859 23490
rect 10927 23434 10983 23490
rect 11051 23434 11107 23490
rect 11175 23434 11231 23490
rect 11299 23434 11355 23490
rect 11423 23434 11479 23490
rect 11547 23434 11603 23490
rect 11671 23434 11727 23490
rect 11795 23434 11851 23490
rect 11919 23434 11975 23490
rect 12043 23434 12099 23490
rect 12167 23434 12223 23490
rect 12291 23434 12347 23490
rect 12415 23434 12471 23490
rect 10679 23310 10735 23366
rect 10803 23310 10859 23366
rect 10927 23310 10983 23366
rect 11051 23310 11107 23366
rect 11175 23310 11231 23366
rect 11299 23310 11355 23366
rect 11423 23310 11479 23366
rect 11547 23310 11603 23366
rect 11671 23310 11727 23366
rect 11795 23310 11851 23366
rect 11919 23310 11975 23366
rect 12043 23310 12099 23366
rect 12167 23310 12223 23366
rect 12291 23310 12347 23366
rect 12415 23310 12471 23366
rect 10679 23186 10735 23242
rect 10803 23186 10859 23242
rect 10927 23186 10983 23242
rect 11051 23186 11107 23242
rect 11175 23186 11231 23242
rect 11299 23186 11355 23242
rect 11423 23186 11479 23242
rect 11547 23186 11603 23242
rect 11671 23186 11727 23242
rect 11795 23186 11851 23242
rect 11919 23186 11975 23242
rect 12043 23186 12099 23242
rect 12167 23186 12223 23242
rect 12291 23186 12347 23242
rect 12415 23186 12471 23242
rect 10679 23062 10735 23118
rect 10803 23062 10859 23118
rect 10927 23062 10983 23118
rect 11051 23062 11107 23118
rect 11175 23062 11231 23118
rect 11299 23062 11355 23118
rect 11423 23062 11479 23118
rect 11547 23062 11603 23118
rect 11671 23062 11727 23118
rect 11795 23062 11851 23118
rect 11919 23062 11975 23118
rect 12043 23062 12099 23118
rect 12167 23062 12223 23118
rect 12291 23062 12347 23118
rect 12415 23062 12471 23118
rect 10679 22938 10735 22994
rect 10803 22938 10859 22994
rect 10927 22938 10983 22994
rect 11051 22938 11107 22994
rect 11175 22938 11231 22994
rect 11299 22938 11355 22994
rect 11423 22938 11479 22994
rect 11547 22938 11603 22994
rect 11671 22938 11727 22994
rect 11795 22938 11851 22994
rect 11919 22938 11975 22994
rect 12043 22938 12099 22994
rect 12167 22938 12223 22994
rect 12291 22938 12347 22994
rect 12415 22938 12471 22994
rect 10679 22814 10735 22870
rect 10803 22814 10859 22870
rect 10927 22814 10983 22870
rect 11051 22814 11107 22870
rect 11175 22814 11231 22870
rect 11299 22814 11355 22870
rect 11423 22814 11479 22870
rect 11547 22814 11603 22870
rect 11671 22814 11727 22870
rect 11795 22814 11851 22870
rect 11919 22814 11975 22870
rect 12043 22814 12099 22870
rect 12167 22814 12223 22870
rect 12291 22814 12347 22870
rect 12415 22814 12471 22870
rect 10679 22690 10735 22746
rect 10803 22690 10859 22746
rect 10927 22690 10983 22746
rect 11051 22690 11107 22746
rect 11175 22690 11231 22746
rect 11299 22690 11355 22746
rect 11423 22690 11479 22746
rect 11547 22690 11603 22746
rect 11671 22690 11727 22746
rect 11795 22690 11851 22746
rect 11919 22690 11975 22746
rect 12043 22690 12099 22746
rect 12167 22690 12223 22746
rect 12291 22690 12347 22746
rect 12415 22690 12471 22746
rect 10679 22566 10735 22622
rect 10803 22566 10859 22622
rect 10927 22566 10983 22622
rect 11051 22566 11107 22622
rect 11175 22566 11231 22622
rect 11299 22566 11355 22622
rect 11423 22566 11479 22622
rect 11547 22566 11603 22622
rect 11671 22566 11727 22622
rect 11795 22566 11851 22622
rect 11919 22566 11975 22622
rect 12043 22566 12099 22622
rect 12167 22566 12223 22622
rect 12291 22566 12347 22622
rect 12415 22566 12471 22622
rect 10679 22442 10735 22498
rect 10803 22442 10859 22498
rect 10927 22442 10983 22498
rect 11051 22442 11107 22498
rect 11175 22442 11231 22498
rect 11299 22442 11355 22498
rect 11423 22442 11479 22498
rect 11547 22442 11603 22498
rect 11671 22442 11727 22498
rect 11795 22442 11851 22498
rect 11919 22442 11975 22498
rect 12043 22442 12099 22498
rect 12167 22442 12223 22498
rect 12291 22442 12347 22498
rect 12415 22442 12471 22498
rect 1078 22094 1134 22150
rect 1202 22094 1258 22150
rect 1326 22094 1382 22150
rect 1450 22094 1506 22150
rect 1574 22094 1630 22150
rect 1698 22094 1754 22150
rect 1822 22094 1878 22150
rect 1946 22094 2002 22150
rect 2070 22094 2126 22150
rect 1078 21970 1134 22026
rect 1202 21970 1258 22026
rect 1326 21970 1382 22026
rect 1450 21970 1506 22026
rect 1574 21970 1630 22026
rect 1698 21970 1754 22026
rect 1822 21970 1878 22026
rect 1946 21970 2002 22026
rect 2070 21970 2126 22026
rect 1078 21846 1134 21902
rect 1202 21846 1258 21902
rect 1326 21846 1382 21902
rect 1450 21846 1506 21902
rect 1574 21846 1630 21902
rect 1698 21846 1754 21902
rect 1822 21846 1878 21902
rect 1946 21846 2002 21902
rect 2070 21846 2126 21902
rect 1078 21722 1134 21778
rect 1202 21722 1258 21778
rect 1326 21722 1382 21778
rect 1450 21722 1506 21778
rect 1574 21722 1630 21778
rect 1698 21722 1754 21778
rect 1822 21722 1878 21778
rect 1946 21722 2002 21778
rect 2070 21722 2126 21778
rect 1078 21598 1134 21654
rect 1202 21598 1258 21654
rect 1326 21598 1382 21654
rect 1450 21598 1506 21654
rect 1574 21598 1630 21654
rect 1698 21598 1754 21654
rect 1822 21598 1878 21654
rect 1946 21598 2002 21654
rect 2070 21598 2126 21654
rect 1078 21474 1134 21530
rect 1202 21474 1258 21530
rect 1326 21474 1382 21530
rect 1450 21474 1506 21530
rect 1574 21474 1630 21530
rect 1698 21474 1754 21530
rect 1822 21474 1878 21530
rect 1946 21474 2002 21530
rect 2070 21474 2126 21530
rect 1078 21350 1134 21406
rect 1202 21350 1258 21406
rect 1326 21350 1382 21406
rect 1450 21350 1506 21406
rect 1574 21350 1630 21406
rect 1698 21350 1754 21406
rect 1822 21350 1878 21406
rect 1946 21350 2002 21406
rect 2070 21350 2126 21406
rect 1078 21226 1134 21282
rect 1202 21226 1258 21282
rect 1326 21226 1382 21282
rect 1450 21226 1506 21282
rect 1574 21226 1630 21282
rect 1698 21226 1754 21282
rect 1822 21226 1878 21282
rect 1946 21226 2002 21282
rect 2070 21226 2126 21282
rect 1078 21102 1134 21158
rect 1202 21102 1258 21158
rect 1326 21102 1382 21158
rect 1450 21102 1506 21158
rect 1574 21102 1630 21158
rect 1698 21102 1754 21158
rect 1822 21102 1878 21158
rect 1946 21102 2002 21158
rect 2070 21102 2126 21158
rect 1078 20978 1134 21034
rect 1202 20978 1258 21034
rect 1326 20978 1382 21034
rect 1450 20978 1506 21034
rect 1574 20978 1630 21034
rect 1698 20978 1754 21034
rect 1822 20978 1878 21034
rect 1946 20978 2002 21034
rect 2070 20978 2126 21034
rect 1078 20854 1134 20910
rect 1202 20854 1258 20910
rect 1326 20854 1382 20910
rect 1450 20854 1506 20910
rect 1574 20854 1630 20910
rect 1698 20854 1754 20910
rect 1822 20854 1878 20910
rect 1946 20854 2002 20910
rect 2070 20854 2126 20910
rect 1078 20730 1134 20786
rect 1202 20730 1258 20786
rect 1326 20730 1382 20786
rect 1450 20730 1506 20786
rect 1574 20730 1630 20786
rect 1698 20730 1754 20786
rect 1822 20730 1878 20786
rect 1946 20730 2002 20786
rect 2070 20730 2126 20786
rect 1078 20606 1134 20662
rect 1202 20606 1258 20662
rect 1326 20606 1382 20662
rect 1450 20606 1506 20662
rect 1574 20606 1630 20662
rect 1698 20606 1754 20662
rect 1822 20606 1878 20662
rect 1946 20606 2002 20662
rect 2070 20606 2126 20662
rect 1078 20482 1134 20538
rect 1202 20482 1258 20538
rect 1326 20482 1382 20538
rect 1450 20482 1506 20538
rect 1574 20482 1630 20538
rect 1698 20482 1754 20538
rect 1822 20482 1878 20538
rect 1946 20482 2002 20538
rect 2070 20482 2126 20538
rect 1078 20358 1134 20414
rect 1202 20358 1258 20414
rect 1326 20358 1382 20414
rect 1450 20358 1506 20414
rect 1574 20358 1630 20414
rect 1698 20358 1754 20414
rect 1822 20358 1878 20414
rect 1946 20358 2002 20414
rect 2070 20358 2126 20414
rect 1078 20234 1134 20290
rect 1202 20234 1258 20290
rect 1326 20234 1382 20290
rect 1450 20234 1506 20290
rect 1574 20234 1630 20290
rect 1698 20234 1754 20290
rect 1822 20234 1878 20290
rect 1946 20234 2002 20290
rect 2070 20234 2126 20290
rect 1078 20110 1134 20166
rect 1202 20110 1258 20166
rect 1326 20110 1382 20166
rect 1450 20110 1506 20166
rect 1574 20110 1630 20166
rect 1698 20110 1754 20166
rect 1822 20110 1878 20166
rect 1946 20110 2002 20166
rect 2070 20110 2126 20166
rect 1078 19986 1134 20042
rect 1202 19986 1258 20042
rect 1326 19986 1382 20042
rect 1450 19986 1506 20042
rect 1574 19986 1630 20042
rect 1698 19986 1754 20042
rect 1822 19986 1878 20042
rect 1946 19986 2002 20042
rect 2070 19986 2126 20042
rect 1078 19862 1134 19918
rect 1202 19862 1258 19918
rect 1326 19862 1382 19918
rect 1450 19862 1506 19918
rect 1574 19862 1630 19918
rect 1698 19862 1754 19918
rect 1822 19862 1878 19918
rect 1946 19862 2002 19918
rect 2070 19862 2126 19918
rect 1078 19738 1134 19794
rect 1202 19738 1258 19794
rect 1326 19738 1382 19794
rect 1450 19738 1506 19794
rect 1574 19738 1630 19794
rect 1698 19738 1754 19794
rect 1822 19738 1878 19794
rect 1946 19738 2002 19794
rect 2070 19738 2126 19794
rect 1078 19614 1134 19670
rect 1202 19614 1258 19670
rect 1326 19614 1382 19670
rect 1450 19614 1506 19670
rect 1574 19614 1630 19670
rect 1698 19614 1754 19670
rect 1822 19614 1878 19670
rect 1946 19614 2002 19670
rect 2070 19614 2126 19670
rect 1078 19490 1134 19546
rect 1202 19490 1258 19546
rect 1326 19490 1382 19546
rect 1450 19490 1506 19546
rect 1574 19490 1630 19546
rect 1698 19490 1754 19546
rect 1822 19490 1878 19546
rect 1946 19490 2002 19546
rect 2070 19490 2126 19546
rect 1078 19366 1134 19422
rect 1202 19366 1258 19422
rect 1326 19366 1382 19422
rect 1450 19366 1506 19422
rect 1574 19366 1630 19422
rect 1698 19366 1754 19422
rect 1822 19366 1878 19422
rect 1946 19366 2002 19422
rect 2070 19366 2126 19422
rect 1078 19242 1134 19298
rect 1202 19242 1258 19298
rect 1326 19242 1382 19298
rect 1450 19242 1506 19298
rect 1574 19242 1630 19298
rect 1698 19242 1754 19298
rect 1822 19242 1878 19298
rect 1946 19242 2002 19298
rect 2070 19242 2126 19298
rect 4435 22094 4491 22150
rect 4559 22094 4615 22150
rect 4683 22094 4739 22150
rect 4807 22094 4863 22150
rect 4931 22094 4987 22150
rect 5055 22094 5111 22150
rect 5179 22094 5235 22150
rect 5303 22094 5359 22150
rect 5427 22094 5483 22150
rect 5551 22094 5607 22150
rect 5675 22094 5731 22150
rect 5799 22094 5855 22150
rect 5923 22094 5979 22150
rect 6047 22094 6103 22150
rect 6171 22094 6227 22150
rect 4435 21970 4491 22026
rect 4559 21970 4615 22026
rect 4683 21970 4739 22026
rect 4807 21970 4863 22026
rect 4931 21970 4987 22026
rect 5055 21970 5111 22026
rect 5179 21970 5235 22026
rect 5303 21970 5359 22026
rect 5427 21970 5483 22026
rect 5551 21970 5607 22026
rect 5675 21970 5731 22026
rect 5799 21970 5855 22026
rect 5923 21970 5979 22026
rect 6047 21970 6103 22026
rect 6171 21970 6227 22026
rect 4435 21846 4491 21902
rect 4559 21846 4615 21902
rect 4683 21846 4739 21902
rect 4807 21846 4863 21902
rect 4931 21846 4987 21902
rect 5055 21846 5111 21902
rect 5179 21846 5235 21902
rect 5303 21846 5359 21902
rect 5427 21846 5483 21902
rect 5551 21846 5607 21902
rect 5675 21846 5731 21902
rect 5799 21846 5855 21902
rect 5923 21846 5979 21902
rect 6047 21846 6103 21902
rect 6171 21846 6227 21902
rect 4435 21722 4491 21778
rect 4559 21722 4615 21778
rect 4683 21722 4739 21778
rect 4807 21722 4863 21778
rect 4931 21722 4987 21778
rect 5055 21722 5111 21778
rect 5179 21722 5235 21778
rect 5303 21722 5359 21778
rect 5427 21722 5483 21778
rect 5551 21722 5607 21778
rect 5675 21722 5731 21778
rect 5799 21722 5855 21778
rect 5923 21722 5979 21778
rect 6047 21722 6103 21778
rect 6171 21722 6227 21778
rect 4435 21598 4491 21654
rect 4559 21598 4615 21654
rect 4683 21598 4739 21654
rect 4807 21598 4863 21654
rect 4931 21598 4987 21654
rect 5055 21598 5111 21654
rect 5179 21598 5235 21654
rect 5303 21598 5359 21654
rect 5427 21598 5483 21654
rect 5551 21598 5607 21654
rect 5675 21598 5731 21654
rect 5799 21598 5855 21654
rect 5923 21598 5979 21654
rect 6047 21598 6103 21654
rect 6171 21598 6227 21654
rect 4435 21474 4491 21530
rect 4559 21474 4615 21530
rect 4683 21474 4739 21530
rect 4807 21474 4863 21530
rect 4931 21474 4987 21530
rect 5055 21474 5111 21530
rect 5179 21474 5235 21530
rect 5303 21474 5359 21530
rect 5427 21474 5483 21530
rect 5551 21474 5607 21530
rect 5675 21474 5731 21530
rect 5799 21474 5855 21530
rect 5923 21474 5979 21530
rect 6047 21474 6103 21530
rect 6171 21474 6227 21530
rect 4435 21350 4491 21406
rect 4559 21350 4615 21406
rect 4683 21350 4739 21406
rect 4807 21350 4863 21406
rect 4931 21350 4987 21406
rect 5055 21350 5111 21406
rect 5179 21350 5235 21406
rect 5303 21350 5359 21406
rect 5427 21350 5483 21406
rect 5551 21350 5607 21406
rect 5675 21350 5731 21406
rect 5799 21350 5855 21406
rect 5923 21350 5979 21406
rect 6047 21350 6103 21406
rect 6171 21350 6227 21406
rect 4435 21226 4491 21282
rect 4559 21226 4615 21282
rect 4683 21226 4739 21282
rect 4807 21226 4863 21282
rect 4931 21226 4987 21282
rect 5055 21226 5111 21282
rect 5179 21226 5235 21282
rect 5303 21226 5359 21282
rect 5427 21226 5483 21282
rect 5551 21226 5607 21282
rect 5675 21226 5731 21282
rect 5799 21226 5855 21282
rect 5923 21226 5979 21282
rect 6047 21226 6103 21282
rect 6171 21226 6227 21282
rect 4435 21102 4491 21158
rect 4559 21102 4615 21158
rect 4683 21102 4739 21158
rect 4807 21102 4863 21158
rect 4931 21102 4987 21158
rect 5055 21102 5111 21158
rect 5179 21102 5235 21158
rect 5303 21102 5359 21158
rect 5427 21102 5483 21158
rect 5551 21102 5607 21158
rect 5675 21102 5731 21158
rect 5799 21102 5855 21158
rect 5923 21102 5979 21158
rect 6047 21102 6103 21158
rect 6171 21102 6227 21158
rect 4435 20978 4491 21034
rect 4559 20978 4615 21034
rect 4683 20978 4739 21034
rect 4807 20978 4863 21034
rect 4931 20978 4987 21034
rect 5055 20978 5111 21034
rect 5179 20978 5235 21034
rect 5303 20978 5359 21034
rect 5427 20978 5483 21034
rect 5551 20978 5607 21034
rect 5675 20978 5731 21034
rect 5799 20978 5855 21034
rect 5923 20978 5979 21034
rect 6047 20978 6103 21034
rect 6171 20978 6227 21034
rect 4435 20854 4491 20910
rect 4559 20854 4615 20910
rect 4683 20854 4739 20910
rect 4807 20854 4863 20910
rect 4931 20854 4987 20910
rect 5055 20854 5111 20910
rect 5179 20854 5235 20910
rect 5303 20854 5359 20910
rect 5427 20854 5483 20910
rect 5551 20854 5607 20910
rect 5675 20854 5731 20910
rect 5799 20854 5855 20910
rect 5923 20854 5979 20910
rect 6047 20854 6103 20910
rect 6171 20854 6227 20910
rect 4435 20730 4491 20786
rect 4559 20730 4615 20786
rect 4683 20730 4739 20786
rect 4807 20730 4863 20786
rect 4931 20730 4987 20786
rect 5055 20730 5111 20786
rect 5179 20730 5235 20786
rect 5303 20730 5359 20786
rect 5427 20730 5483 20786
rect 5551 20730 5607 20786
rect 5675 20730 5731 20786
rect 5799 20730 5855 20786
rect 5923 20730 5979 20786
rect 6047 20730 6103 20786
rect 6171 20730 6227 20786
rect 4435 20606 4491 20662
rect 4559 20606 4615 20662
rect 4683 20606 4739 20662
rect 4807 20606 4863 20662
rect 4931 20606 4987 20662
rect 5055 20606 5111 20662
rect 5179 20606 5235 20662
rect 5303 20606 5359 20662
rect 5427 20606 5483 20662
rect 5551 20606 5607 20662
rect 5675 20606 5731 20662
rect 5799 20606 5855 20662
rect 5923 20606 5979 20662
rect 6047 20606 6103 20662
rect 6171 20606 6227 20662
rect 4435 20482 4491 20538
rect 4559 20482 4615 20538
rect 4683 20482 4739 20538
rect 4807 20482 4863 20538
rect 4931 20482 4987 20538
rect 5055 20482 5111 20538
rect 5179 20482 5235 20538
rect 5303 20482 5359 20538
rect 5427 20482 5483 20538
rect 5551 20482 5607 20538
rect 5675 20482 5731 20538
rect 5799 20482 5855 20538
rect 5923 20482 5979 20538
rect 6047 20482 6103 20538
rect 6171 20482 6227 20538
rect 4435 20358 4491 20414
rect 4559 20358 4615 20414
rect 4683 20358 4739 20414
rect 4807 20358 4863 20414
rect 4931 20358 4987 20414
rect 5055 20358 5111 20414
rect 5179 20358 5235 20414
rect 5303 20358 5359 20414
rect 5427 20358 5483 20414
rect 5551 20358 5607 20414
rect 5675 20358 5731 20414
rect 5799 20358 5855 20414
rect 5923 20358 5979 20414
rect 6047 20358 6103 20414
rect 6171 20358 6227 20414
rect 4435 20234 4491 20290
rect 4559 20234 4615 20290
rect 4683 20234 4739 20290
rect 4807 20234 4863 20290
rect 4931 20234 4987 20290
rect 5055 20234 5111 20290
rect 5179 20234 5235 20290
rect 5303 20234 5359 20290
rect 5427 20234 5483 20290
rect 5551 20234 5607 20290
rect 5675 20234 5731 20290
rect 5799 20234 5855 20290
rect 5923 20234 5979 20290
rect 6047 20234 6103 20290
rect 6171 20234 6227 20290
rect 4435 20110 4491 20166
rect 4559 20110 4615 20166
rect 4683 20110 4739 20166
rect 4807 20110 4863 20166
rect 4931 20110 4987 20166
rect 5055 20110 5111 20166
rect 5179 20110 5235 20166
rect 5303 20110 5359 20166
rect 5427 20110 5483 20166
rect 5551 20110 5607 20166
rect 5675 20110 5731 20166
rect 5799 20110 5855 20166
rect 5923 20110 5979 20166
rect 6047 20110 6103 20166
rect 6171 20110 6227 20166
rect 4435 19986 4491 20042
rect 4559 19986 4615 20042
rect 4683 19986 4739 20042
rect 4807 19986 4863 20042
rect 4931 19986 4987 20042
rect 5055 19986 5111 20042
rect 5179 19986 5235 20042
rect 5303 19986 5359 20042
rect 5427 19986 5483 20042
rect 5551 19986 5607 20042
rect 5675 19986 5731 20042
rect 5799 19986 5855 20042
rect 5923 19986 5979 20042
rect 6047 19986 6103 20042
rect 6171 19986 6227 20042
rect 4435 19862 4491 19918
rect 4559 19862 4615 19918
rect 4683 19862 4739 19918
rect 4807 19862 4863 19918
rect 4931 19862 4987 19918
rect 5055 19862 5111 19918
rect 5179 19862 5235 19918
rect 5303 19862 5359 19918
rect 5427 19862 5483 19918
rect 5551 19862 5607 19918
rect 5675 19862 5731 19918
rect 5799 19862 5855 19918
rect 5923 19862 5979 19918
rect 6047 19862 6103 19918
rect 6171 19862 6227 19918
rect 4435 19738 4491 19794
rect 4559 19738 4615 19794
rect 4683 19738 4739 19794
rect 4807 19738 4863 19794
rect 4931 19738 4987 19794
rect 5055 19738 5111 19794
rect 5179 19738 5235 19794
rect 5303 19738 5359 19794
rect 5427 19738 5483 19794
rect 5551 19738 5607 19794
rect 5675 19738 5731 19794
rect 5799 19738 5855 19794
rect 5923 19738 5979 19794
rect 6047 19738 6103 19794
rect 6171 19738 6227 19794
rect 4435 19614 4491 19670
rect 4559 19614 4615 19670
rect 4683 19614 4739 19670
rect 4807 19614 4863 19670
rect 4931 19614 4987 19670
rect 5055 19614 5111 19670
rect 5179 19614 5235 19670
rect 5303 19614 5359 19670
rect 5427 19614 5483 19670
rect 5551 19614 5607 19670
rect 5675 19614 5731 19670
rect 5799 19614 5855 19670
rect 5923 19614 5979 19670
rect 6047 19614 6103 19670
rect 6171 19614 6227 19670
rect 4435 19490 4491 19546
rect 4559 19490 4615 19546
rect 4683 19490 4739 19546
rect 4807 19490 4863 19546
rect 4931 19490 4987 19546
rect 5055 19490 5111 19546
rect 5179 19490 5235 19546
rect 5303 19490 5359 19546
rect 5427 19490 5483 19546
rect 5551 19490 5607 19546
rect 5675 19490 5731 19546
rect 5799 19490 5855 19546
rect 5923 19490 5979 19546
rect 6047 19490 6103 19546
rect 6171 19490 6227 19546
rect 4435 19366 4491 19422
rect 4559 19366 4615 19422
rect 4683 19366 4739 19422
rect 4807 19366 4863 19422
rect 4931 19366 4987 19422
rect 5055 19366 5111 19422
rect 5179 19366 5235 19422
rect 5303 19366 5359 19422
rect 5427 19366 5483 19422
rect 5551 19366 5607 19422
rect 5675 19366 5731 19422
rect 5799 19366 5855 19422
rect 5923 19366 5979 19422
rect 6047 19366 6103 19422
rect 6171 19366 6227 19422
rect 4435 19242 4491 19298
rect 4559 19242 4615 19298
rect 4683 19242 4739 19298
rect 4807 19242 4863 19298
rect 4931 19242 4987 19298
rect 5055 19242 5111 19298
rect 5179 19242 5235 19298
rect 5303 19242 5359 19298
rect 5427 19242 5483 19298
rect 5551 19242 5607 19298
rect 5675 19242 5731 19298
rect 5799 19242 5855 19298
rect 5923 19242 5979 19298
rect 6047 19242 6103 19298
rect 6171 19242 6227 19298
rect 7562 22094 7618 22150
rect 7686 22094 7742 22150
rect 7810 22094 7866 22150
rect 7934 22094 7990 22150
rect 8058 22094 8114 22150
rect 8182 22094 8238 22150
rect 8306 22094 8362 22150
rect 8430 22094 8486 22150
rect 8554 22094 8610 22150
rect 7562 21970 7618 22026
rect 7686 21970 7742 22026
rect 7810 21970 7866 22026
rect 7934 21970 7990 22026
rect 8058 21970 8114 22026
rect 8182 21970 8238 22026
rect 8306 21970 8362 22026
rect 8430 21970 8486 22026
rect 8554 21970 8610 22026
rect 7562 21846 7618 21902
rect 7686 21846 7742 21902
rect 7810 21846 7866 21902
rect 7934 21846 7990 21902
rect 8058 21846 8114 21902
rect 8182 21846 8238 21902
rect 8306 21846 8362 21902
rect 8430 21846 8486 21902
rect 8554 21846 8610 21902
rect 7562 21722 7618 21778
rect 7686 21722 7742 21778
rect 7810 21722 7866 21778
rect 7934 21722 7990 21778
rect 8058 21722 8114 21778
rect 8182 21722 8238 21778
rect 8306 21722 8362 21778
rect 8430 21722 8486 21778
rect 8554 21722 8610 21778
rect 7562 21598 7618 21654
rect 7686 21598 7742 21654
rect 7810 21598 7866 21654
rect 7934 21598 7990 21654
rect 8058 21598 8114 21654
rect 8182 21598 8238 21654
rect 8306 21598 8362 21654
rect 8430 21598 8486 21654
rect 8554 21598 8610 21654
rect 7562 21474 7618 21530
rect 7686 21474 7742 21530
rect 7810 21474 7866 21530
rect 7934 21474 7990 21530
rect 8058 21474 8114 21530
rect 8182 21474 8238 21530
rect 8306 21474 8362 21530
rect 8430 21474 8486 21530
rect 8554 21474 8610 21530
rect 7562 21350 7618 21406
rect 7686 21350 7742 21406
rect 7810 21350 7866 21406
rect 7934 21350 7990 21406
rect 8058 21350 8114 21406
rect 8182 21350 8238 21406
rect 8306 21350 8362 21406
rect 8430 21350 8486 21406
rect 8554 21350 8610 21406
rect 7562 21226 7618 21282
rect 7686 21226 7742 21282
rect 7810 21226 7866 21282
rect 7934 21226 7990 21282
rect 8058 21226 8114 21282
rect 8182 21226 8238 21282
rect 8306 21226 8362 21282
rect 8430 21226 8486 21282
rect 8554 21226 8610 21282
rect 7562 21102 7618 21158
rect 7686 21102 7742 21158
rect 7810 21102 7866 21158
rect 7934 21102 7990 21158
rect 8058 21102 8114 21158
rect 8182 21102 8238 21158
rect 8306 21102 8362 21158
rect 8430 21102 8486 21158
rect 8554 21102 8610 21158
rect 7562 20978 7618 21034
rect 7686 20978 7742 21034
rect 7810 20978 7866 21034
rect 7934 20978 7990 21034
rect 8058 20978 8114 21034
rect 8182 20978 8238 21034
rect 8306 20978 8362 21034
rect 8430 20978 8486 21034
rect 8554 20978 8610 21034
rect 7562 20854 7618 20910
rect 7686 20854 7742 20910
rect 7810 20854 7866 20910
rect 7934 20854 7990 20910
rect 8058 20854 8114 20910
rect 8182 20854 8238 20910
rect 8306 20854 8362 20910
rect 8430 20854 8486 20910
rect 8554 20854 8610 20910
rect 7562 20730 7618 20786
rect 7686 20730 7742 20786
rect 7810 20730 7866 20786
rect 7934 20730 7990 20786
rect 8058 20730 8114 20786
rect 8182 20730 8238 20786
rect 8306 20730 8362 20786
rect 8430 20730 8486 20786
rect 8554 20730 8610 20786
rect 7562 20606 7618 20662
rect 7686 20606 7742 20662
rect 7810 20606 7866 20662
rect 7934 20606 7990 20662
rect 8058 20606 8114 20662
rect 8182 20606 8238 20662
rect 8306 20606 8362 20662
rect 8430 20606 8486 20662
rect 8554 20606 8610 20662
rect 7562 20482 7618 20538
rect 7686 20482 7742 20538
rect 7810 20482 7866 20538
rect 7934 20482 7990 20538
rect 8058 20482 8114 20538
rect 8182 20482 8238 20538
rect 8306 20482 8362 20538
rect 8430 20482 8486 20538
rect 8554 20482 8610 20538
rect 7562 20358 7618 20414
rect 7686 20358 7742 20414
rect 7810 20358 7866 20414
rect 7934 20358 7990 20414
rect 8058 20358 8114 20414
rect 8182 20358 8238 20414
rect 8306 20358 8362 20414
rect 8430 20358 8486 20414
rect 8554 20358 8610 20414
rect 7562 20234 7618 20290
rect 7686 20234 7742 20290
rect 7810 20234 7866 20290
rect 7934 20234 7990 20290
rect 8058 20234 8114 20290
rect 8182 20234 8238 20290
rect 8306 20234 8362 20290
rect 8430 20234 8486 20290
rect 8554 20234 8610 20290
rect 7562 20110 7618 20166
rect 7686 20110 7742 20166
rect 7810 20110 7866 20166
rect 7934 20110 7990 20166
rect 8058 20110 8114 20166
rect 8182 20110 8238 20166
rect 8306 20110 8362 20166
rect 8430 20110 8486 20166
rect 8554 20110 8610 20166
rect 7562 19986 7618 20042
rect 7686 19986 7742 20042
rect 7810 19986 7866 20042
rect 7934 19986 7990 20042
rect 8058 19986 8114 20042
rect 8182 19986 8238 20042
rect 8306 19986 8362 20042
rect 8430 19986 8486 20042
rect 8554 19986 8610 20042
rect 7562 19862 7618 19918
rect 7686 19862 7742 19918
rect 7810 19862 7866 19918
rect 7934 19862 7990 19918
rect 8058 19862 8114 19918
rect 8182 19862 8238 19918
rect 8306 19862 8362 19918
rect 8430 19862 8486 19918
rect 8554 19862 8610 19918
rect 7562 19738 7618 19794
rect 7686 19738 7742 19794
rect 7810 19738 7866 19794
rect 7934 19738 7990 19794
rect 8058 19738 8114 19794
rect 8182 19738 8238 19794
rect 8306 19738 8362 19794
rect 8430 19738 8486 19794
rect 8554 19738 8610 19794
rect 7562 19614 7618 19670
rect 7686 19614 7742 19670
rect 7810 19614 7866 19670
rect 7934 19614 7990 19670
rect 8058 19614 8114 19670
rect 8182 19614 8238 19670
rect 8306 19614 8362 19670
rect 8430 19614 8486 19670
rect 8554 19614 8610 19670
rect 7562 19490 7618 19546
rect 7686 19490 7742 19546
rect 7810 19490 7866 19546
rect 7934 19490 7990 19546
rect 8058 19490 8114 19546
rect 8182 19490 8238 19546
rect 8306 19490 8362 19546
rect 8430 19490 8486 19546
rect 8554 19490 8610 19546
rect 7562 19366 7618 19422
rect 7686 19366 7742 19422
rect 7810 19366 7866 19422
rect 7934 19366 7990 19422
rect 8058 19366 8114 19422
rect 8182 19366 8238 19422
rect 8306 19366 8362 19422
rect 8430 19366 8486 19422
rect 8554 19366 8610 19422
rect 7562 19242 7618 19298
rect 7686 19242 7742 19298
rect 7810 19242 7866 19298
rect 7934 19242 7990 19298
rect 8058 19242 8114 19298
rect 8182 19242 8238 19298
rect 8306 19242 8362 19298
rect 8430 19242 8486 19298
rect 8554 19242 8610 19298
rect 10679 22094 10735 22150
rect 10803 22094 10859 22150
rect 10927 22094 10983 22150
rect 11051 22094 11107 22150
rect 11175 22094 11231 22150
rect 11299 22094 11355 22150
rect 11423 22094 11479 22150
rect 11547 22094 11603 22150
rect 11671 22094 11727 22150
rect 11795 22094 11851 22150
rect 11919 22094 11975 22150
rect 12043 22094 12099 22150
rect 12167 22094 12223 22150
rect 12291 22094 12347 22150
rect 12415 22094 12471 22150
rect 10679 21970 10735 22026
rect 10803 21970 10859 22026
rect 10927 21970 10983 22026
rect 11051 21970 11107 22026
rect 11175 21970 11231 22026
rect 11299 21970 11355 22026
rect 11423 21970 11479 22026
rect 11547 21970 11603 22026
rect 11671 21970 11727 22026
rect 11795 21970 11851 22026
rect 11919 21970 11975 22026
rect 12043 21970 12099 22026
rect 12167 21970 12223 22026
rect 12291 21970 12347 22026
rect 12415 21970 12471 22026
rect 10679 21846 10735 21902
rect 10803 21846 10859 21902
rect 10927 21846 10983 21902
rect 11051 21846 11107 21902
rect 11175 21846 11231 21902
rect 11299 21846 11355 21902
rect 11423 21846 11479 21902
rect 11547 21846 11603 21902
rect 11671 21846 11727 21902
rect 11795 21846 11851 21902
rect 11919 21846 11975 21902
rect 12043 21846 12099 21902
rect 12167 21846 12223 21902
rect 12291 21846 12347 21902
rect 12415 21846 12471 21902
rect 10679 21722 10735 21778
rect 10803 21722 10859 21778
rect 10927 21722 10983 21778
rect 11051 21722 11107 21778
rect 11175 21722 11231 21778
rect 11299 21722 11355 21778
rect 11423 21722 11479 21778
rect 11547 21722 11603 21778
rect 11671 21722 11727 21778
rect 11795 21722 11851 21778
rect 11919 21722 11975 21778
rect 12043 21722 12099 21778
rect 12167 21722 12223 21778
rect 12291 21722 12347 21778
rect 12415 21722 12471 21778
rect 10679 21598 10735 21654
rect 10803 21598 10859 21654
rect 10927 21598 10983 21654
rect 11051 21598 11107 21654
rect 11175 21598 11231 21654
rect 11299 21598 11355 21654
rect 11423 21598 11479 21654
rect 11547 21598 11603 21654
rect 11671 21598 11727 21654
rect 11795 21598 11851 21654
rect 11919 21598 11975 21654
rect 12043 21598 12099 21654
rect 12167 21598 12223 21654
rect 12291 21598 12347 21654
rect 12415 21598 12471 21654
rect 10679 21474 10735 21530
rect 10803 21474 10859 21530
rect 10927 21474 10983 21530
rect 11051 21474 11107 21530
rect 11175 21474 11231 21530
rect 11299 21474 11355 21530
rect 11423 21474 11479 21530
rect 11547 21474 11603 21530
rect 11671 21474 11727 21530
rect 11795 21474 11851 21530
rect 11919 21474 11975 21530
rect 12043 21474 12099 21530
rect 12167 21474 12223 21530
rect 12291 21474 12347 21530
rect 12415 21474 12471 21530
rect 10679 21350 10735 21406
rect 10803 21350 10859 21406
rect 10927 21350 10983 21406
rect 11051 21350 11107 21406
rect 11175 21350 11231 21406
rect 11299 21350 11355 21406
rect 11423 21350 11479 21406
rect 11547 21350 11603 21406
rect 11671 21350 11727 21406
rect 11795 21350 11851 21406
rect 11919 21350 11975 21406
rect 12043 21350 12099 21406
rect 12167 21350 12223 21406
rect 12291 21350 12347 21406
rect 12415 21350 12471 21406
rect 10679 21226 10735 21282
rect 10803 21226 10859 21282
rect 10927 21226 10983 21282
rect 11051 21226 11107 21282
rect 11175 21226 11231 21282
rect 11299 21226 11355 21282
rect 11423 21226 11479 21282
rect 11547 21226 11603 21282
rect 11671 21226 11727 21282
rect 11795 21226 11851 21282
rect 11919 21226 11975 21282
rect 12043 21226 12099 21282
rect 12167 21226 12223 21282
rect 12291 21226 12347 21282
rect 12415 21226 12471 21282
rect 10679 21102 10735 21158
rect 10803 21102 10859 21158
rect 10927 21102 10983 21158
rect 11051 21102 11107 21158
rect 11175 21102 11231 21158
rect 11299 21102 11355 21158
rect 11423 21102 11479 21158
rect 11547 21102 11603 21158
rect 11671 21102 11727 21158
rect 11795 21102 11851 21158
rect 11919 21102 11975 21158
rect 12043 21102 12099 21158
rect 12167 21102 12223 21158
rect 12291 21102 12347 21158
rect 12415 21102 12471 21158
rect 10679 20978 10735 21034
rect 10803 20978 10859 21034
rect 10927 20978 10983 21034
rect 11051 20978 11107 21034
rect 11175 20978 11231 21034
rect 11299 20978 11355 21034
rect 11423 20978 11479 21034
rect 11547 20978 11603 21034
rect 11671 20978 11727 21034
rect 11795 20978 11851 21034
rect 11919 20978 11975 21034
rect 12043 20978 12099 21034
rect 12167 20978 12223 21034
rect 12291 20978 12347 21034
rect 12415 20978 12471 21034
rect 10679 20854 10735 20910
rect 10803 20854 10859 20910
rect 10927 20854 10983 20910
rect 11051 20854 11107 20910
rect 11175 20854 11231 20910
rect 11299 20854 11355 20910
rect 11423 20854 11479 20910
rect 11547 20854 11603 20910
rect 11671 20854 11727 20910
rect 11795 20854 11851 20910
rect 11919 20854 11975 20910
rect 12043 20854 12099 20910
rect 12167 20854 12223 20910
rect 12291 20854 12347 20910
rect 12415 20854 12471 20910
rect 10679 20730 10735 20786
rect 10803 20730 10859 20786
rect 10927 20730 10983 20786
rect 11051 20730 11107 20786
rect 11175 20730 11231 20786
rect 11299 20730 11355 20786
rect 11423 20730 11479 20786
rect 11547 20730 11603 20786
rect 11671 20730 11727 20786
rect 11795 20730 11851 20786
rect 11919 20730 11975 20786
rect 12043 20730 12099 20786
rect 12167 20730 12223 20786
rect 12291 20730 12347 20786
rect 12415 20730 12471 20786
rect 10679 20606 10735 20662
rect 10803 20606 10859 20662
rect 10927 20606 10983 20662
rect 11051 20606 11107 20662
rect 11175 20606 11231 20662
rect 11299 20606 11355 20662
rect 11423 20606 11479 20662
rect 11547 20606 11603 20662
rect 11671 20606 11727 20662
rect 11795 20606 11851 20662
rect 11919 20606 11975 20662
rect 12043 20606 12099 20662
rect 12167 20606 12223 20662
rect 12291 20606 12347 20662
rect 12415 20606 12471 20662
rect 10679 20482 10735 20538
rect 10803 20482 10859 20538
rect 10927 20482 10983 20538
rect 11051 20482 11107 20538
rect 11175 20482 11231 20538
rect 11299 20482 11355 20538
rect 11423 20482 11479 20538
rect 11547 20482 11603 20538
rect 11671 20482 11727 20538
rect 11795 20482 11851 20538
rect 11919 20482 11975 20538
rect 12043 20482 12099 20538
rect 12167 20482 12223 20538
rect 12291 20482 12347 20538
rect 12415 20482 12471 20538
rect 10679 20358 10735 20414
rect 10803 20358 10859 20414
rect 10927 20358 10983 20414
rect 11051 20358 11107 20414
rect 11175 20358 11231 20414
rect 11299 20358 11355 20414
rect 11423 20358 11479 20414
rect 11547 20358 11603 20414
rect 11671 20358 11727 20414
rect 11795 20358 11851 20414
rect 11919 20358 11975 20414
rect 12043 20358 12099 20414
rect 12167 20358 12223 20414
rect 12291 20358 12347 20414
rect 12415 20358 12471 20414
rect 10679 20234 10735 20290
rect 10803 20234 10859 20290
rect 10927 20234 10983 20290
rect 11051 20234 11107 20290
rect 11175 20234 11231 20290
rect 11299 20234 11355 20290
rect 11423 20234 11479 20290
rect 11547 20234 11603 20290
rect 11671 20234 11727 20290
rect 11795 20234 11851 20290
rect 11919 20234 11975 20290
rect 12043 20234 12099 20290
rect 12167 20234 12223 20290
rect 12291 20234 12347 20290
rect 12415 20234 12471 20290
rect 10679 20110 10735 20166
rect 10803 20110 10859 20166
rect 10927 20110 10983 20166
rect 11051 20110 11107 20166
rect 11175 20110 11231 20166
rect 11299 20110 11355 20166
rect 11423 20110 11479 20166
rect 11547 20110 11603 20166
rect 11671 20110 11727 20166
rect 11795 20110 11851 20166
rect 11919 20110 11975 20166
rect 12043 20110 12099 20166
rect 12167 20110 12223 20166
rect 12291 20110 12347 20166
rect 12415 20110 12471 20166
rect 10679 19986 10735 20042
rect 10803 19986 10859 20042
rect 10927 19986 10983 20042
rect 11051 19986 11107 20042
rect 11175 19986 11231 20042
rect 11299 19986 11355 20042
rect 11423 19986 11479 20042
rect 11547 19986 11603 20042
rect 11671 19986 11727 20042
rect 11795 19986 11851 20042
rect 11919 19986 11975 20042
rect 12043 19986 12099 20042
rect 12167 19986 12223 20042
rect 12291 19986 12347 20042
rect 12415 19986 12471 20042
rect 10679 19862 10735 19918
rect 10803 19862 10859 19918
rect 10927 19862 10983 19918
rect 11051 19862 11107 19918
rect 11175 19862 11231 19918
rect 11299 19862 11355 19918
rect 11423 19862 11479 19918
rect 11547 19862 11603 19918
rect 11671 19862 11727 19918
rect 11795 19862 11851 19918
rect 11919 19862 11975 19918
rect 12043 19862 12099 19918
rect 12167 19862 12223 19918
rect 12291 19862 12347 19918
rect 12415 19862 12471 19918
rect 10679 19738 10735 19794
rect 10803 19738 10859 19794
rect 10927 19738 10983 19794
rect 11051 19738 11107 19794
rect 11175 19738 11231 19794
rect 11299 19738 11355 19794
rect 11423 19738 11479 19794
rect 11547 19738 11603 19794
rect 11671 19738 11727 19794
rect 11795 19738 11851 19794
rect 11919 19738 11975 19794
rect 12043 19738 12099 19794
rect 12167 19738 12223 19794
rect 12291 19738 12347 19794
rect 12415 19738 12471 19794
rect 10679 19614 10735 19670
rect 10803 19614 10859 19670
rect 10927 19614 10983 19670
rect 11051 19614 11107 19670
rect 11175 19614 11231 19670
rect 11299 19614 11355 19670
rect 11423 19614 11479 19670
rect 11547 19614 11603 19670
rect 11671 19614 11727 19670
rect 11795 19614 11851 19670
rect 11919 19614 11975 19670
rect 12043 19614 12099 19670
rect 12167 19614 12223 19670
rect 12291 19614 12347 19670
rect 12415 19614 12471 19670
rect 10679 19490 10735 19546
rect 10803 19490 10859 19546
rect 10927 19490 10983 19546
rect 11051 19490 11107 19546
rect 11175 19490 11231 19546
rect 11299 19490 11355 19546
rect 11423 19490 11479 19546
rect 11547 19490 11603 19546
rect 11671 19490 11727 19546
rect 11795 19490 11851 19546
rect 11919 19490 11975 19546
rect 12043 19490 12099 19546
rect 12167 19490 12223 19546
rect 12291 19490 12347 19546
rect 12415 19490 12471 19546
rect 10679 19366 10735 19422
rect 10803 19366 10859 19422
rect 10927 19366 10983 19422
rect 11051 19366 11107 19422
rect 11175 19366 11231 19422
rect 11299 19366 11355 19422
rect 11423 19366 11479 19422
rect 11547 19366 11603 19422
rect 11671 19366 11727 19422
rect 11795 19366 11851 19422
rect 11919 19366 11975 19422
rect 12043 19366 12099 19422
rect 12167 19366 12223 19422
rect 12291 19366 12347 19422
rect 12415 19366 12471 19422
rect 10679 19242 10735 19298
rect 10803 19242 10859 19298
rect 10927 19242 10983 19298
rect 11051 19242 11107 19298
rect 11175 19242 11231 19298
rect 11299 19242 11355 19298
rect 11423 19242 11479 19298
rect 11547 19242 11603 19298
rect 11671 19242 11727 19298
rect 11795 19242 11851 19298
rect 11919 19242 11975 19298
rect 12043 19242 12099 19298
rect 12167 19242 12223 19298
rect 12291 19242 12347 19298
rect 12415 19242 12471 19298
rect 1078 18894 1134 18950
rect 1202 18894 1258 18950
rect 1326 18894 1382 18950
rect 1450 18894 1506 18950
rect 1574 18894 1630 18950
rect 1698 18894 1754 18950
rect 1822 18894 1878 18950
rect 1946 18894 2002 18950
rect 2070 18894 2126 18950
rect 1078 18770 1134 18826
rect 1202 18770 1258 18826
rect 1326 18770 1382 18826
rect 1450 18770 1506 18826
rect 1574 18770 1630 18826
rect 1698 18770 1754 18826
rect 1822 18770 1878 18826
rect 1946 18770 2002 18826
rect 2070 18770 2126 18826
rect 1078 18646 1134 18702
rect 1202 18646 1258 18702
rect 1326 18646 1382 18702
rect 1450 18646 1506 18702
rect 1574 18646 1630 18702
rect 1698 18646 1754 18702
rect 1822 18646 1878 18702
rect 1946 18646 2002 18702
rect 2070 18646 2126 18702
rect 1078 18522 1134 18578
rect 1202 18522 1258 18578
rect 1326 18522 1382 18578
rect 1450 18522 1506 18578
rect 1574 18522 1630 18578
rect 1698 18522 1754 18578
rect 1822 18522 1878 18578
rect 1946 18522 2002 18578
rect 2070 18522 2126 18578
rect 1078 18398 1134 18454
rect 1202 18398 1258 18454
rect 1326 18398 1382 18454
rect 1450 18398 1506 18454
rect 1574 18398 1630 18454
rect 1698 18398 1754 18454
rect 1822 18398 1878 18454
rect 1946 18398 2002 18454
rect 2070 18398 2126 18454
rect 1078 18274 1134 18330
rect 1202 18274 1258 18330
rect 1326 18274 1382 18330
rect 1450 18274 1506 18330
rect 1574 18274 1630 18330
rect 1698 18274 1754 18330
rect 1822 18274 1878 18330
rect 1946 18274 2002 18330
rect 2070 18274 2126 18330
rect 1078 18150 1134 18206
rect 1202 18150 1258 18206
rect 1326 18150 1382 18206
rect 1450 18150 1506 18206
rect 1574 18150 1630 18206
rect 1698 18150 1754 18206
rect 1822 18150 1878 18206
rect 1946 18150 2002 18206
rect 2070 18150 2126 18206
rect 1078 18026 1134 18082
rect 1202 18026 1258 18082
rect 1326 18026 1382 18082
rect 1450 18026 1506 18082
rect 1574 18026 1630 18082
rect 1698 18026 1754 18082
rect 1822 18026 1878 18082
rect 1946 18026 2002 18082
rect 2070 18026 2126 18082
rect 1078 17902 1134 17958
rect 1202 17902 1258 17958
rect 1326 17902 1382 17958
rect 1450 17902 1506 17958
rect 1574 17902 1630 17958
rect 1698 17902 1754 17958
rect 1822 17902 1878 17958
rect 1946 17902 2002 17958
rect 2070 17902 2126 17958
rect 1078 17778 1134 17834
rect 1202 17778 1258 17834
rect 1326 17778 1382 17834
rect 1450 17778 1506 17834
rect 1574 17778 1630 17834
rect 1698 17778 1754 17834
rect 1822 17778 1878 17834
rect 1946 17778 2002 17834
rect 2070 17778 2126 17834
rect 1078 17654 1134 17710
rect 1202 17654 1258 17710
rect 1326 17654 1382 17710
rect 1450 17654 1506 17710
rect 1574 17654 1630 17710
rect 1698 17654 1754 17710
rect 1822 17654 1878 17710
rect 1946 17654 2002 17710
rect 2070 17654 2126 17710
rect 1078 17530 1134 17586
rect 1202 17530 1258 17586
rect 1326 17530 1382 17586
rect 1450 17530 1506 17586
rect 1574 17530 1630 17586
rect 1698 17530 1754 17586
rect 1822 17530 1878 17586
rect 1946 17530 2002 17586
rect 2070 17530 2126 17586
rect 1078 17406 1134 17462
rect 1202 17406 1258 17462
rect 1326 17406 1382 17462
rect 1450 17406 1506 17462
rect 1574 17406 1630 17462
rect 1698 17406 1754 17462
rect 1822 17406 1878 17462
rect 1946 17406 2002 17462
rect 2070 17406 2126 17462
rect 1078 17282 1134 17338
rect 1202 17282 1258 17338
rect 1326 17282 1382 17338
rect 1450 17282 1506 17338
rect 1574 17282 1630 17338
rect 1698 17282 1754 17338
rect 1822 17282 1878 17338
rect 1946 17282 2002 17338
rect 2070 17282 2126 17338
rect 1078 17158 1134 17214
rect 1202 17158 1258 17214
rect 1326 17158 1382 17214
rect 1450 17158 1506 17214
rect 1574 17158 1630 17214
rect 1698 17158 1754 17214
rect 1822 17158 1878 17214
rect 1946 17158 2002 17214
rect 2070 17158 2126 17214
rect 1078 17034 1134 17090
rect 1202 17034 1258 17090
rect 1326 17034 1382 17090
rect 1450 17034 1506 17090
rect 1574 17034 1630 17090
rect 1698 17034 1754 17090
rect 1822 17034 1878 17090
rect 1946 17034 2002 17090
rect 2070 17034 2126 17090
rect 1078 16910 1134 16966
rect 1202 16910 1258 16966
rect 1326 16910 1382 16966
rect 1450 16910 1506 16966
rect 1574 16910 1630 16966
rect 1698 16910 1754 16966
rect 1822 16910 1878 16966
rect 1946 16910 2002 16966
rect 2070 16910 2126 16966
rect 1078 16786 1134 16842
rect 1202 16786 1258 16842
rect 1326 16786 1382 16842
rect 1450 16786 1506 16842
rect 1574 16786 1630 16842
rect 1698 16786 1754 16842
rect 1822 16786 1878 16842
rect 1946 16786 2002 16842
rect 2070 16786 2126 16842
rect 1078 16662 1134 16718
rect 1202 16662 1258 16718
rect 1326 16662 1382 16718
rect 1450 16662 1506 16718
rect 1574 16662 1630 16718
rect 1698 16662 1754 16718
rect 1822 16662 1878 16718
rect 1946 16662 2002 16718
rect 2070 16662 2126 16718
rect 1078 16538 1134 16594
rect 1202 16538 1258 16594
rect 1326 16538 1382 16594
rect 1450 16538 1506 16594
rect 1574 16538 1630 16594
rect 1698 16538 1754 16594
rect 1822 16538 1878 16594
rect 1946 16538 2002 16594
rect 2070 16538 2126 16594
rect 1078 16414 1134 16470
rect 1202 16414 1258 16470
rect 1326 16414 1382 16470
rect 1450 16414 1506 16470
rect 1574 16414 1630 16470
rect 1698 16414 1754 16470
rect 1822 16414 1878 16470
rect 1946 16414 2002 16470
rect 2070 16414 2126 16470
rect 1078 16290 1134 16346
rect 1202 16290 1258 16346
rect 1326 16290 1382 16346
rect 1450 16290 1506 16346
rect 1574 16290 1630 16346
rect 1698 16290 1754 16346
rect 1822 16290 1878 16346
rect 1946 16290 2002 16346
rect 2070 16290 2126 16346
rect 1078 16166 1134 16222
rect 1202 16166 1258 16222
rect 1326 16166 1382 16222
rect 1450 16166 1506 16222
rect 1574 16166 1630 16222
rect 1698 16166 1754 16222
rect 1822 16166 1878 16222
rect 1946 16166 2002 16222
rect 2070 16166 2126 16222
rect 1078 16042 1134 16098
rect 1202 16042 1258 16098
rect 1326 16042 1382 16098
rect 1450 16042 1506 16098
rect 1574 16042 1630 16098
rect 1698 16042 1754 16098
rect 1822 16042 1878 16098
rect 1946 16042 2002 16098
rect 2070 16042 2126 16098
rect 4435 18894 4491 18950
rect 4559 18894 4615 18950
rect 4683 18894 4739 18950
rect 4807 18894 4863 18950
rect 4931 18894 4987 18950
rect 5055 18894 5111 18950
rect 5179 18894 5235 18950
rect 5303 18894 5359 18950
rect 5427 18894 5483 18950
rect 5551 18894 5607 18950
rect 5675 18894 5731 18950
rect 5799 18894 5855 18950
rect 5923 18894 5979 18950
rect 6047 18894 6103 18950
rect 6171 18894 6227 18950
rect 4435 18770 4491 18826
rect 4559 18770 4615 18826
rect 4683 18770 4739 18826
rect 4807 18770 4863 18826
rect 4931 18770 4987 18826
rect 5055 18770 5111 18826
rect 5179 18770 5235 18826
rect 5303 18770 5359 18826
rect 5427 18770 5483 18826
rect 5551 18770 5607 18826
rect 5675 18770 5731 18826
rect 5799 18770 5855 18826
rect 5923 18770 5979 18826
rect 6047 18770 6103 18826
rect 6171 18770 6227 18826
rect 4435 18646 4491 18702
rect 4559 18646 4615 18702
rect 4683 18646 4739 18702
rect 4807 18646 4863 18702
rect 4931 18646 4987 18702
rect 5055 18646 5111 18702
rect 5179 18646 5235 18702
rect 5303 18646 5359 18702
rect 5427 18646 5483 18702
rect 5551 18646 5607 18702
rect 5675 18646 5731 18702
rect 5799 18646 5855 18702
rect 5923 18646 5979 18702
rect 6047 18646 6103 18702
rect 6171 18646 6227 18702
rect 4435 18522 4491 18578
rect 4559 18522 4615 18578
rect 4683 18522 4739 18578
rect 4807 18522 4863 18578
rect 4931 18522 4987 18578
rect 5055 18522 5111 18578
rect 5179 18522 5235 18578
rect 5303 18522 5359 18578
rect 5427 18522 5483 18578
rect 5551 18522 5607 18578
rect 5675 18522 5731 18578
rect 5799 18522 5855 18578
rect 5923 18522 5979 18578
rect 6047 18522 6103 18578
rect 6171 18522 6227 18578
rect 4435 18398 4491 18454
rect 4559 18398 4615 18454
rect 4683 18398 4739 18454
rect 4807 18398 4863 18454
rect 4931 18398 4987 18454
rect 5055 18398 5111 18454
rect 5179 18398 5235 18454
rect 5303 18398 5359 18454
rect 5427 18398 5483 18454
rect 5551 18398 5607 18454
rect 5675 18398 5731 18454
rect 5799 18398 5855 18454
rect 5923 18398 5979 18454
rect 6047 18398 6103 18454
rect 6171 18398 6227 18454
rect 4435 18274 4491 18330
rect 4559 18274 4615 18330
rect 4683 18274 4739 18330
rect 4807 18274 4863 18330
rect 4931 18274 4987 18330
rect 5055 18274 5111 18330
rect 5179 18274 5235 18330
rect 5303 18274 5359 18330
rect 5427 18274 5483 18330
rect 5551 18274 5607 18330
rect 5675 18274 5731 18330
rect 5799 18274 5855 18330
rect 5923 18274 5979 18330
rect 6047 18274 6103 18330
rect 6171 18274 6227 18330
rect 4435 18150 4491 18206
rect 4559 18150 4615 18206
rect 4683 18150 4739 18206
rect 4807 18150 4863 18206
rect 4931 18150 4987 18206
rect 5055 18150 5111 18206
rect 5179 18150 5235 18206
rect 5303 18150 5359 18206
rect 5427 18150 5483 18206
rect 5551 18150 5607 18206
rect 5675 18150 5731 18206
rect 5799 18150 5855 18206
rect 5923 18150 5979 18206
rect 6047 18150 6103 18206
rect 6171 18150 6227 18206
rect 4435 18026 4491 18082
rect 4559 18026 4615 18082
rect 4683 18026 4739 18082
rect 4807 18026 4863 18082
rect 4931 18026 4987 18082
rect 5055 18026 5111 18082
rect 5179 18026 5235 18082
rect 5303 18026 5359 18082
rect 5427 18026 5483 18082
rect 5551 18026 5607 18082
rect 5675 18026 5731 18082
rect 5799 18026 5855 18082
rect 5923 18026 5979 18082
rect 6047 18026 6103 18082
rect 6171 18026 6227 18082
rect 4435 17902 4491 17958
rect 4559 17902 4615 17958
rect 4683 17902 4739 17958
rect 4807 17902 4863 17958
rect 4931 17902 4987 17958
rect 5055 17902 5111 17958
rect 5179 17902 5235 17958
rect 5303 17902 5359 17958
rect 5427 17902 5483 17958
rect 5551 17902 5607 17958
rect 5675 17902 5731 17958
rect 5799 17902 5855 17958
rect 5923 17902 5979 17958
rect 6047 17902 6103 17958
rect 6171 17902 6227 17958
rect 4435 17778 4491 17834
rect 4559 17778 4615 17834
rect 4683 17778 4739 17834
rect 4807 17778 4863 17834
rect 4931 17778 4987 17834
rect 5055 17778 5111 17834
rect 5179 17778 5235 17834
rect 5303 17778 5359 17834
rect 5427 17778 5483 17834
rect 5551 17778 5607 17834
rect 5675 17778 5731 17834
rect 5799 17778 5855 17834
rect 5923 17778 5979 17834
rect 6047 17778 6103 17834
rect 6171 17778 6227 17834
rect 4435 17654 4491 17710
rect 4559 17654 4615 17710
rect 4683 17654 4739 17710
rect 4807 17654 4863 17710
rect 4931 17654 4987 17710
rect 5055 17654 5111 17710
rect 5179 17654 5235 17710
rect 5303 17654 5359 17710
rect 5427 17654 5483 17710
rect 5551 17654 5607 17710
rect 5675 17654 5731 17710
rect 5799 17654 5855 17710
rect 5923 17654 5979 17710
rect 6047 17654 6103 17710
rect 6171 17654 6227 17710
rect 4435 17530 4491 17586
rect 4559 17530 4615 17586
rect 4683 17530 4739 17586
rect 4807 17530 4863 17586
rect 4931 17530 4987 17586
rect 5055 17530 5111 17586
rect 5179 17530 5235 17586
rect 5303 17530 5359 17586
rect 5427 17530 5483 17586
rect 5551 17530 5607 17586
rect 5675 17530 5731 17586
rect 5799 17530 5855 17586
rect 5923 17530 5979 17586
rect 6047 17530 6103 17586
rect 6171 17530 6227 17586
rect 4435 17406 4491 17462
rect 4559 17406 4615 17462
rect 4683 17406 4739 17462
rect 4807 17406 4863 17462
rect 4931 17406 4987 17462
rect 5055 17406 5111 17462
rect 5179 17406 5235 17462
rect 5303 17406 5359 17462
rect 5427 17406 5483 17462
rect 5551 17406 5607 17462
rect 5675 17406 5731 17462
rect 5799 17406 5855 17462
rect 5923 17406 5979 17462
rect 6047 17406 6103 17462
rect 6171 17406 6227 17462
rect 4435 17282 4491 17338
rect 4559 17282 4615 17338
rect 4683 17282 4739 17338
rect 4807 17282 4863 17338
rect 4931 17282 4987 17338
rect 5055 17282 5111 17338
rect 5179 17282 5235 17338
rect 5303 17282 5359 17338
rect 5427 17282 5483 17338
rect 5551 17282 5607 17338
rect 5675 17282 5731 17338
rect 5799 17282 5855 17338
rect 5923 17282 5979 17338
rect 6047 17282 6103 17338
rect 6171 17282 6227 17338
rect 4435 17158 4491 17214
rect 4559 17158 4615 17214
rect 4683 17158 4739 17214
rect 4807 17158 4863 17214
rect 4931 17158 4987 17214
rect 5055 17158 5111 17214
rect 5179 17158 5235 17214
rect 5303 17158 5359 17214
rect 5427 17158 5483 17214
rect 5551 17158 5607 17214
rect 5675 17158 5731 17214
rect 5799 17158 5855 17214
rect 5923 17158 5979 17214
rect 6047 17158 6103 17214
rect 6171 17158 6227 17214
rect 4435 17034 4491 17090
rect 4559 17034 4615 17090
rect 4683 17034 4739 17090
rect 4807 17034 4863 17090
rect 4931 17034 4987 17090
rect 5055 17034 5111 17090
rect 5179 17034 5235 17090
rect 5303 17034 5359 17090
rect 5427 17034 5483 17090
rect 5551 17034 5607 17090
rect 5675 17034 5731 17090
rect 5799 17034 5855 17090
rect 5923 17034 5979 17090
rect 6047 17034 6103 17090
rect 6171 17034 6227 17090
rect 4435 16910 4491 16966
rect 4559 16910 4615 16966
rect 4683 16910 4739 16966
rect 4807 16910 4863 16966
rect 4931 16910 4987 16966
rect 5055 16910 5111 16966
rect 5179 16910 5235 16966
rect 5303 16910 5359 16966
rect 5427 16910 5483 16966
rect 5551 16910 5607 16966
rect 5675 16910 5731 16966
rect 5799 16910 5855 16966
rect 5923 16910 5979 16966
rect 6047 16910 6103 16966
rect 6171 16910 6227 16966
rect 4435 16786 4491 16842
rect 4559 16786 4615 16842
rect 4683 16786 4739 16842
rect 4807 16786 4863 16842
rect 4931 16786 4987 16842
rect 5055 16786 5111 16842
rect 5179 16786 5235 16842
rect 5303 16786 5359 16842
rect 5427 16786 5483 16842
rect 5551 16786 5607 16842
rect 5675 16786 5731 16842
rect 5799 16786 5855 16842
rect 5923 16786 5979 16842
rect 6047 16786 6103 16842
rect 6171 16786 6227 16842
rect 4435 16662 4491 16718
rect 4559 16662 4615 16718
rect 4683 16662 4739 16718
rect 4807 16662 4863 16718
rect 4931 16662 4987 16718
rect 5055 16662 5111 16718
rect 5179 16662 5235 16718
rect 5303 16662 5359 16718
rect 5427 16662 5483 16718
rect 5551 16662 5607 16718
rect 5675 16662 5731 16718
rect 5799 16662 5855 16718
rect 5923 16662 5979 16718
rect 6047 16662 6103 16718
rect 6171 16662 6227 16718
rect 4435 16538 4491 16594
rect 4559 16538 4615 16594
rect 4683 16538 4739 16594
rect 4807 16538 4863 16594
rect 4931 16538 4987 16594
rect 5055 16538 5111 16594
rect 5179 16538 5235 16594
rect 5303 16538 5359 16594
rect 5427 16538 5483 16594
rect 5551 16538 5607 16594
rect 5675 16538 5731 16594
rect 5799 16538 5855 16594
rect 5923 16538 5979 16594
rect 6047 16538 6103 16594
rect 6171 16538 6227 16594
rect 4435 16414 4491 16470
rect 4559 16414 4615 16470
rect 4683 16414 4739 16470
rect 4807 16414 4863 16470
rect 4931 16414 4987 16470
rect 5055 16414 5111 16470
rect 5179 16414 5235 16470
rect 5303 16414 5359 16470
rect 5427 16414 5483 16470
rect 5551 16414 5607 16470
rect 5675 16414 5731 16470
rect 5799 16414 5855 16470
rect 5923 16414 5979 16470
rect 6047 16414 6103 16470
rect 6171 16414 6227 16470
rect 4435 16290 4491 16346
rect 4559 16290 4615 16346
rect 4683 16290 4739 16346
rect 4807 16290 4863 16346
rect 4931 16290 4987 16346
rect 5055 16290 5111 16346
rect 5179 16290 5235 16346
rect 5303 16290 5359 16346
rect 5427 16290 5483 16346
rect 5551 16290 5607 16346
rect 5675 16290 5731 16346
rect 5799 16290 5855 16346
rect 5923 16290 5979 16346
rect 6047 16290 6103 16346
rect 6171 16290 6227 16346
rect 4435 16166 4491 16222
rect 4559 16166 4615 16222
rect 4683 16166 4739 16222
rect 4807 16166 4863 16222
rect 4931 16166 4987 16222
rect 5055 16166 5111 16222
rect 5179 16166 5235 16222
rect 5303 16166 5359 16222
rect 5427 16166 5483 16222
rect 5551 16166 5607 16222
rect 5675 16166 5731 16222
rect 5799 16166 5855 16222
rect 5923 16166 5979 16222
rect 6047 16166 6103 16222
rect 6171 16166 6227 16222
rect 4435 16042 4491 16098
rect 4559 16042 4615 16098
rect 4683 16042 4739 16098
rect 4807 16042 4863 16098
rect 4931 16042 4987 16098
rect 5055 16042 5111 16098
rect 5179 16042 5235 16098
rect 5303 16042 5359 16098
rect 5427 16042 5483 16098
rect 5551 16042 5607 16098
rect 5675 16042 5731 16098
rect 5799 16042 5855 16098
rect 5923 16042 5979 16098
rect 6047 16042 6103 16098
rect 6171 16042 6227 16098
rect 7562 18894 7618 18950
rect 7686 18894 7742 18950
rect 7810 18894 7866 18950
rect 7934 18894 7990 18950
rect 8058 18894 8114 18950
rect 8182 18894 8238 18950
rect 8306 18894 8362 18950
rect 8430 18894 8486 18950
rect 8554 18894 8610 18950
rect 7562 18770 7618 18826
rect 7686 18770 7742 18826
rect 7810 18770 7866 18826
rect 7934 18770 7990 18826
rect 8058 18770 8114 18826
rect 8182 18770 8238 18826
rect 8306 18770 8362 18826
rect 8430 18770 8486 18826
rect 8554 18770 8610 18826
rect 7562 18646 7618 18702
rect 7686 18646 7742 18702
rect 7810 18646 7866 18702
rect 7934 18646 7990 18702
rect 8058 18646 8114 18702
rect 8182 18646 8238 18702
rect 8306 18646 8362 18702
rect 8430 18646 8486 18702
rect 8554 18646 8610 18702
rect 7562 18522 7618 18578
rect 7686 18522 7742 18578
rect 7810 18522 7866 18578
rect 7934 18522 7990 18578
rect 8058 18522 8114 18578
rect 8182 18522 8238 18578
rect 8306 18522 8362 18578
rect 8430 18522 8486 18578
rect 8554 18522 8610 18578
rect 7562 18398 7618 18454
rect 7686 18398 7742 18454
rect 7810 18398 7866 18454
rect 7934 18398 7990 18454
rect 8058 18398 8114 18454
rect 8182 18398 8238 18454
rect 8306 18398 8362 18454
rect 8430 18398 8486 18454
rect 8554 18398 8610 18454
rect 7562 18274 7618 18330
rect 7686 18274 7742 18330
rect 7810 18274 7866 18330
rect 7934 18274 7990 18330
rect 8058 18274 8114 18330
rect 8182 18274 8238 18330
rect 8306 18274 8362 18330
rect 8430 18274 8486 18330
rect 8554 18274 8610 18330
rect 7562 18150 7618 18206
rect 7686 18150 7742 18206
rect 7810 18150 7866 18206
rect 7934 18150 7990 18206
rect 8058 18150 8114 18206
rect 8182 18150 8238 18206
rect 8306 18150 8362 18206
rect 8430 18150 8486 18206
rect 8554 18150 8610 18206
rect 7562 18026 7618 18082
rect 7686 18026 7742 18082
rect 7810 18026 7866 18082
rect 7934 18026 7990 18082
rect 8058 18026 8114 18082
rect 8182 18026 8238 18082
rect 8306 18026 8362 18082
rect 8430 18026 8486 18082
rect 8554 18026 8610 18082
rect 7562 17902 7618 17958
rect 7686 17902 7742 17958
rect 7810 17902 7866 17958
rect 7934 17902 7990 17958
rect 8058 17902 8114 17958
rect 8182 17902 8238 17958
rect 8306 17902 8362 17958
rect 8430 17902 8486 17958
rect 8554 17902 8610 17958
rect 7562 17778 7618 17834
rect 7686 17778 7742 17834
rect 7810 17778 7866 17834
rect 7934 17778 7990 17834
rect 8058 17778 8114 17834
rect 8182 17778 8238 17834
rect 8306 17778 8362 17834
rect 8430 17778 8486 17834
rect 8554 17778 8610 17834
rect 7562 17654 7618 17710
rect 7686 17654 7742 17710
rect 7810 17654 7866 17710
rect 7934 17654 7990 17710
rect 8058 17654 8114 17710
rect 8182 17654 8238 17710
rect 8306 17654 8362 17710
rect 8430 17654 8486 17710
rect 8554 17654 8610 17710
rect 7562 17530 7618 17586
rect 7686 17530 7742 17586
rect 7810 17530 7866 17586
rect 7934 17530 7990 17586
rect 8058 17530 8114 17586
rect 8182 17530 8238 17586
rect 8306 17530 8362 17586
rect 8430 17530 8486 17586
rect 8554 17530 8610 17586
rect 7562 17406 7618 17462
rect 7686 17406 7742 17462
rect 7810 17406 7866 17462
rect 7934 17406 7990 17462
rect 8058 17406 8114 17462
rect 8182 17406 8238 17462
rect 8306 17406 8362 17462
rect 8430 17406 8486 17462
rect 8554 17406 8610 17462
rect 7562 17282 7618 17338
rect 7686 17282 7742 17338
rect 7810 17282 7866 17338
rect 7934 17282 7990 17338
rect 8058 17282 8114 17338
rect 8182 17282 8238 17338
rect 8306 17282 8362 17338
rect 8430 17282 8486 17338
rect 8554 17282 8610 17338
rect 7562 17158 7618 17214
rect 7686 17158 7742 17214
rect 7810 17158 7866 17214
rect 7934 17158 7990 17214
rect 8058 17158 8114 17214
rect 8182 17158 8238 17214
rect 8306 17158 8362 17214
rect 8430 17158 8486 17214
rect 8554 17158 8610 17214
rect 7562 17034 7618 17090
rect 7686 17034 7742 17090
rect 7810 17034 7866 17090
rect 7934 17034 7990 17090
rect 8058 17034 8114 17090
rect 8182 17034 8238 17090
rect 8306 17034 8362 17090
rect 8430 17034 8486 17090
rect 8554 17034 8610 17090
rect 7562 16910 7618 16966
rect 7686 16910 7742 16966
rect 7810 16910 7866 16966
rect 7934 16910 7990 16966
rect 8058 16910 8114 16966
rect 8182 16910 8238 16966
rect 8306 16910 8362 16966
rect 8430 16910 8486 16966
rect 8554 16910 8610 16966
rect 7562 16786 7618 16842
rect 7686 16786 7742 16842
rect 7810 16786 7866 16842
rect 7934 16786 7990 16842
rect 8058 16786 8114 16842
rect 8182 16786 8238 16842
rect 8306 16786 8362 16842
rect 8430 16786 8486 16842
rect 8554 16786 8610 16842
rect 7562 16662 7618 16718
rect 7686 16662 7742 16718
rect 7810 16662 7866 16718
rect 7934 16662 7990 16718
rect 8058 16662 8114 16718
rect 8182 16662 8238 16718
rect 8306 16662 8362 16718
rect 8430 16662 8486 16718
rect 8554 16662 8610 16718
rect 7562 16538 7618 16594
rect 7686 16538 7742 16594
rect 7810 16538 7866 16594
rect 7934 16538 7990 16594
rect 8058 16538 8114 16594
rect 8182 16538 8238 16594
rect 8306 16538 8362 16594
rect 8430 16538 8486 16594
rect 8554 16538 8610 16594
rect 7562 16414 7618 16470
rect 7686 16414 7742 16470
rect 7810 16414 7866 16470
rect 7934 16414 7990 16470
rect 8058 16414 8114 16470
rect 8182 16414 8238 16470
rect 8306 16414 8362 16470
rect 8430 16414 8486 16470
rect 8554 16414 8610 16470
rect 7562 16290 7618 16346
rect 7686 16290 7742 16346
rect 7810 16290 7866 16346
rect 7934 16290 7990 16346
rect 8058 16290 8114 16346
rect 8182 16290 8238 16346
rect 8306 16290 8362 16346
rect 8430 16290 8486 16346
rect 8554 16290 8610 16346
rect 7562 16166 7618 16222
rect 7686 16166 7742 16222
rect 7810 16166 7866 16222
rect 7934 16166 7990 16222
rect 8058 16166 8114 16222
rect 8182 16166 8238 16222
rect 8306 16166 8362 16222
rect 8430 16166 8486 16222
rect 8554 16166 8610 16222
rect 7562 16042 7618 16098
rect 7686 16042 7742 16098
rect 7810 16042 7866 16098
rect 7934 16042 7990 16098
rect 8058 16042 8114 16098
rect 8182 16042 8238 16098
rect 8306 16042 8362 16098
rect 8430 16042 8486 16098
rect 8554 16042 8610 16098
rect 10679 18894 10735 18950
rect 10803 18894 10859 18950
rect 10927 18894 10983 18950
rect 11051 18894 11107 18950
rect 11175 18894 11231 18950
rect 11299 18894 11355 18950
rect 11423 18894 11479 18950
rect 11547 18894 11603 18950
rect 11671 18894 11727 18950
rect 11795 18894 11851 18950
rect 11919 18894 11975 18950
rect 12043 18894 12099 18950
rect 12167 18894 12223 18950
rect 12291 18894 12347 18950
rect 12415 18894 12471 18950
rect 10679 18770 10735 18826
rect 10803 18770 10859 18826
rect 10927 18770 10983 18826
rect 11051 18770 11107 18826
rect 11175 18770 11231 18826
rect 11299 18770 11355 18826
rect 11423 18770 11479 18826
rect 11547 18770 11603 18826
rect 11671 18770 11727 18826
rect 11795 18770 11851 18826
rect 11919 18770 11975 18826
rect 12043 18770 12099 18826
rect 12167 18770 12223 18826
rect 12291 18770 12347 18826
rect 12415 18770 12471 18826
rect 10679 18646 10735 18702
rect 10803 18646 10859 18702
rect 10927 18646 10983 18702
rect 11051 18646 11107 18702
rect 11175 18646 11231 18702
rect 11299 18646 11355 18702
rect 11423 18646 11479 18702
rect 11547 18646 11603 18702
rect 11671 18646 11727 18702
rect 11795 18646 11851 18702
rect 11919 18646 11975 18702
rect 12043 18646 12099 18702
rect 12167 18646 12223 18702
rect 12291 18646 12347 18702
rect 12415 18646 12471 18702
rect 10679 18522 10735 18578
rect 10803 18522 10859 18578
rect 10927 18522 10983 18578
rect 11051 18522 11107 18578
rect 11175 18522 11231 18578
rect 11299 18522 11355 18578
rect 11423 18522 11479 18578
rect 11547 18522 11603 18578
rect 11671 18522 11727 18578
rect 11795 18522 11851 18578
rect 11919 18522 11975 18578
rect 12043 18522 12099 18578
rect 12167 18522 12223 18578
rect 12291 18522 12347 18578
rect 12415 18522 12471 18578
rect 10679 18398 10735 18454
rect 10803 18398 10859 18454
rect 10927 18398 10983 18454
rect 11051 18398 11107 18454
rect 11175 18398 11231 18454
rect 11299 18398 11355 18454
rect 11423 18398 11479 18454
rect 11547 18398 11603 18454
rect 11671 18398 11727 18454
rect 11795 18398 11851 18454
rect 11919 18398 11975 18454
rect 12043 18398 12099 18454
rect 12167 18398 12223 18454
rect 12291 18398 12347 18454
rect 12415 18398 12471 18454
rect 10679 18274 10735 18330
rect 10803 18274 10859 18330
rect 10927 18274 10983 18330
rect 11051 18274 11107 18330
rect 11175 18274 11231 18330
rect 11299 18274 11355 18330
rect 11423 18274 11479 18330
rect 11547 18274 11603 18330
rect 11671 18274 11727 18330
rect 11795 18274 11851 18330
rect 11919 18274 11975 18330
rect 12043 18274 12099 18330
rect 12167 18274 12223 18330
rect 12291 18274 12347 18330
rect 12415 18274 12471 18330
rect 10679 18150 10735 18206
rect 10803 18150 10859 18206
rect 10927 18150 10983 18206
rect 11051 18150 11107 18206
rect 11175 18150 11231 18206
rect 11299 18150 11355 18206
rect 11423 18150 11479 18206
rect 11547 18150 11603 18206
rect 11671 18150 11727 18206
rect 11795 18150 11851 18206
rect 11919 18150 11975 18206
rect 12043 18150 12099 18206
rect 12167 18150 12223 18206
rect 12291 18150 12347 18206
rect 12415 18150 12471 18206
rect 10679 18026 10735 18082
rect 10803 18026 10859 18082
rect 10927 18026 10983 18082
rect 11051 18026 11107 18082
rect 11175 18026 11231 18082
rect 11299 18026 11355 18082
rect 11423 18026 11479 18082
rect 11547 18026 11603 18082
rect 11671 18026 11727 18082
rect 11795 18026 11851 18082
rect 11919 18026 11975 18082
rect 12043 18026 12099 18082
rect 12167 18026 12223 18082
rect 12291 18026 12347 18082
rect 12415 18026 12471 18082
rect 10679 17902 10735 17958
rect 10803 17902 10859 17958
rect 10927 17902 10983 17958
rect 11051 17902 11107 17958
rect 11175 17902 11231 17958
rect 11299 17902 11355 17958
rect 11423 17902 11479 17958
rect 11547 17902 11603 17958
rect 11671 17902 11727 17958
rect 11795 17902 11851 17958
rect 11919 17902 11975 17958
rect 12043 17902 12099 17958
rect 12167 17902 12223 17958
rect 12291 17902 12347 17958
rect 12415 17902 12471 17958
rect 10679 17778 10735 17834
rect 10803 17778 10859 17834
rect 10927 17778 10983 17834
rect 11051 17778 11107 17834
rect 11175 17778 11231 17834
rect 11299 17778 11355 17834
rect 11423 17778 11479 17834
rect 11547 17778 11603 17834
rect 11671 17778 11727 17834
rect 11795 17778 11851 17834
rect 11919 17778 11975 17834
rect 12043 17778 12099 17834
rect 12167 17778 12223 17834
rect 12291 17778 12347 17834
rect 12415 17778 12471 17834
rect 10679 17654 10735 17710
rect 10803 17654 10859 17710
rect 10927 17654 10983 17710
rect 11051 17654 11107 17710
rect 11175 17654 11231 17710
rect 11299 17654 11355 17710
rect 11423 17654 11479 17710
rect 11547 17654 11603 17710
rect 11671 17654 11727 17710
rect 11795 17654 11851 17710
rect 11919 17654 11975 17710
rect 12043 17654 12099 17710
rect 12167 17654 12223 17710
rect 12291 17654 12347 17710
rect 12415 17654 12471 17710
rect 10679 17530 10735 17586
rect 10803 17530 10859 17586
rect 10927 17530 10983 17586
rect 11051 17530 11107 17586
rect 11175 17530 11231 17586
rect 11299 17530 11355 17586
rect 11423 17530 11479 17586
rect 11547 17530 11603 17586
rect 11671 17530 11727 17586
rect 11795 17530 11851 17586
rect 11919 17530 11975 17586
rect 12043 17530 12099 17586
rect 12167 17530 12223 17586
rect 12291 17530 12347 17586
rect 12415 17530 12471 17586
rect 10679 17406 10735 17462
rect 10803 17406 10859 17462
rect 10927 17406 10983 17462
rect 11051 17406 11107 17462
rect 11175 17406 11231 17462
rect 11299 17406 11355 17462
rect 11423 17406 11479 17462
rect 11547 17406 11603 17462
rect 11671 17406 11727 17462
rect 11795 17406 11851 17462
rect 11919 17406 11975 17462
rect 12043 17406 12099 17462
rect 12167 17406 12223 17462
rect 12291 17406 12347 17462
rect 12415 17406 12471 17462
rect 10679 17282 10735 17338
rect 10803 17282 10859 17338
rect 10927 17282 10983 17338
rect 11051 17282 11107 17338
rect 11175 17282 11231 17338
rect 11299 17282 11355 17338
rect 11423 17282 11479 17338
rect 11547 17282 11603 17338
rect 11671 17282 11727 17338
rect 11795 17282 11851 17338
rect 11919 17282 11975 17338
rect 12043 17282 12099 17338
rect 12167 17282 12223 17338
rect 12291 17282 12347 17338
rect 12415 17282 12471 17338
rect 10679 17158 10735 17214
rect 10803 17158 10859 17214
rect 10927 17158 10983 17214
rect 11051 17158 11107 17214
rect 11175 17158 11231 17214
rect 11299 17158 11355 17214
rect 11423 17158 11479 17214
rect 11547 17158 11603 17214
rect 11671 17158 11727 17214
rect 11795 17158 11851 17214
rect 11919 17158 11975 17214
rect 12043 17158 12099 17214
rect 12167 17158 12223 17214
rect 12291 17158 12347 17214
rect 12415 17158 12471 17214
rect 10679 17034 10735 17090
rect 10803 17034 10859 17090
rect 10927 17034 10983 17090
rect 11051 17034 11107 17090
rect 11175 17034 11231 17090
rect 11299 17034 11355 17090
rect 11423 17034 11479 17090
rect 11547 17034 11603 17090
rect 11671 17034 11727 17090
rect 11795 17034 11851 17090
rect 11919 17034 11975 17090
rect 12043 17034 12099 17090
rect 12167 17034 12223 17090
rect 12291 17034 12347 17090
rect 12415 17034 12471 17090
rect 10679 16910 10735 16966
rect 10803 16910 10859 16966
rect 10927 16910 10983 16966
rect 11051 16910 11107 16966
rect 11175 16910 11231 16966
rect 11299 16910 11355 16966
rect 11423 16910 11479 16966
rect 11547 16910 11603 16966
rect 11671 16910 11727 16966
rect 11795 16910 11851 16966
rect 11919 16910 11975 16966
rect 12043 16910 12099 16966
rect 12167 16910 12223 16966
rect 12291 16910 12347 16966
rect 12415 16910 12471 16966
rect 10679 16786 10735 16842
rect 10803 16786 10859 16842
rect 10927 16786 10983 16842
rect 11051 16786 11107 16842
rect 11175 16786 11231 16842
rect 11299 16786 11355 16842
rect 11423 16786 11479 16842
rect 11547 16786 11603 16842
rect 11671 16786 11727 16842
rect 11795 16786 11851 16842
rect 11919 16786 11975 16842
rect 12043 16786 12099 16842
rect 12167 16786 12223 16842
rect 12291 16786 12347 16842
rect 12415 16786 12471 16842
rect 10679 16662 10735 16718
rect 10803 16662 10859 16718
rect 10927 16662 10983 16718
rect 11051 16662 11107 16718
rect 11175 16662 11231 16718
rect 11299 16662 11355 16718
rect 11423 16662 11479 16718
rect 11547 16662 11603 16718
rect 11671 16662 11727 16718
rect 11795 16662 11851 16718
rect 11919 16662 11975 16718
rect 12043 16662 12099 16718
rect 12167 16662 12223 16718
rect 12291 16662 12347 16718
rect 12415 16662 12471 16718
rect 10679 16538 10735 16594
rect 10803 16538 10859 16594
rect 10927 16538 10983 16594
rect 11051 16538 11107 16594
rect 11175 16538 11231 16594
rect 11299 16538 11355 16594
rect 11423 16538 11479 16594
rect 11547 16538 11603 16594
rect 11671 16538 11727 16594
rect 11795 16538 11851 16594
rect 11919 16538 11975 16594
rect 12043 16538 12099 16594
rect 12167 16538 12223 16594
rect 12291 16538 12347 16594
rect 12415 16538 12471 16594
rect 10679 16414 10735 16470
rect 10803 16414 10859 16470
rect 10927 16414 10983 16470
rect 11051 16414 11107 16470
rect 11175 16414 11231 16470
rect 11299 16414 11355 16470
rect 11423 16414 11479 16470
rect 11547 16414 11603 16470
rect 11671 16414 11727 16470
rect 11795 16414 11851 16470
rect 11919 16414 11975 16470
rect 12043 16414 12099 16470
rect 12167 16414 12223 16470
rect 12291 16414 12347 16470
rect 12415 16414 12471 16470
rect 10679 16290 10735 16346
rect 10803 16290 10859 16346
rect 10927 16290 10983 16346
rect 11051 16290 11107 16346
rect 11175 16290 11231 16346
rect 11299 16290 11355 16346
rect 11423 16290 11479 16346
rect 11547 16290 11603 16346
rect 11671 16290 11727 16346
rect 11795 16290 11851 16346
rect 11919 16290 11975 16346
rect 12043 16290 12099 16346
rect 12167 16290 12223 16346
rect 12291 16290 12347 16346
rect 12415 16290 12471 16346
rect 10679 16166 10735 16222
rect 10803 16166 10859 16222
rect 10927 16166 10983 16222
rect 11051 16166 11107 16222
rect 11175 16166 11231 16222
rect 11299 16166 11355 16222
rect 11423 16166 11479 16222
rect 11547 16166 11603 16222
rect 11671 16166 11727 16222
rect 11795 16166 11851 16222
rect 11919 16166 11975 16222
rect 12043 16166 12099 16222
rect 12167 16166 12223 16222
rect 12291 16166 12347 16222
rect 12415 16166 12471 16222
rect 10679 16042 10735 16098
rect 10803 16042 10859 16098
rect 10927 16042 10983 16098
rect 11051 16042 11107 16098
rect 11175 16042 11231 16098
rect 11299 16042 11355 16098
rect 11423 16042 11479 16098
rect 11547 16042 11603 16098
rect 11671 16042 11727 16098
rect 11795 16042 11851 16098
rect 11919 16042 11975 16098
rect 12043 16042 12099 16098
rect 12167 16042 12223 16098
rect 12291 16042 12347 16098
rect 12415 16042 12471 16098
rect 1078 15694 1134 15750
rect 1202 15694 1258 15750
rect 1326 15694 1382 15750
rect 1450 15694 1506 15750
rect 1574 15694 1630 15750
rect 1698 15694 1754 15750
rect 1822 15694 1878 15750
rect 1946 15694 2002 15750
rect 2070 15694 2126 15750
rect 1078 15570 1134 15626
rect 1202 15570 1258 15626
rect 1326 15570 1382 15626
rect 1450 15570 1506 15626
rect 1574 15570 1630 15626
rect 1698 15570 1754 15626
rect 1822 15570 1878 15626
rect 1946 15570 2002 15626
rect 2070 15570 2126 15626
rect 1078 15446 1134 15502
rect 1202 15446 1258 15502
rect 1326 15446 1382 15502
rect 1450 15446 1506 15502
rect 1574 15446 1630 15502
rect 1698 15446 1754 15502
rect 1822 15446 1878 15502
rect 1946 15446 2002 15502
rect 2070 15446 2126 15502
rect 1078 15322 1134 15378
rect 1202 15322 1258 15378
rect 1326 15322 1382 15378
rect 1450 15322 1506 15378
rect 1574 15322 1630 15378
rect 1698 15322 1754 15378
rect 1822 15322 1878 15378
rect 1946 15322 2002 15378
rect 2070 15322 2126 15378
rect 1078 15198 1134 15254
rect 1202 15198 1258 15254
rect 1326 15198 1382 15254
rect 1450 15198 1506 15254
rect 1574 15198 1630 15254
rect 1698 15198 1754 15254
rect 1822 15198 1878 15254
rect 1946 15198 2002 15254
rect 2070 15198 2126 15254
rect 1078 15074 1134 15130
rect 1202 15074 1258 15130
rect 1326 15074 1382 15130
rect 1450 15074 1506 15130
rect 1574 15074 1630 15130
rect 1698 15074 1754 15130
rect 1822 15074 1878 15130
rect 1946 15074 2002 15130
rect 2070 15074 2126 15130
rect 1078 14950 1134 15006
rect 1202 14950 1258 15006
rect 1326 14950 1382 15006
rect 1450 14950 1506 15006
rect 1574 14950 1630 15006
rect 1698 14950 1754 15006
rect 1822 14950 1878 15006
rect 1946 14950 2002 15006
rect 2070 14950 2126 15006
rect 1078 14826 1134 14882
rect 1202 14826 1258 14882
rect 1326 14826 1382 14882
rect 1450 14826 1506 14882
rect 1574 14826 1630 14882
rect 1698 14826 1754 14882
rect 1822 14826 1878 14882
rect 1946 14826 2002 14882
rect 2070 14826 2126 14882
rect 1078 14702 1134 14758
rect 1202 14702 1258 14758
rect 1326 14702 1382 14758
rect 1450 14702 1506 14758
rect 1574 14702 1630 14758
rect 1698 14702 1754 14758
rect 1822 14702 1878 14758
rect 1946 14702 2002 14758
rect 2070 14702 2126 14758
rect 1078 14578 1134 14634
rect 1202 14578 1258 14634
rect 1326 14578 1382 14634
rect 1450 14578 1506 14634
rect 1574 14578 1630 14634
rect 1698 14578 1754 14634
rect 1822 14578 1878 14634
rect 1946 14578 2002 14634
rect 2070 14578 2126 14634
rect 1078 14454 1134 14510
rect 1202 14454 1258 14510
rect 1326 14454 1382 14510
rect 1450 14454 1506 14510
rect 1574 14454 1630 14510
rect 1698 14454 1754 14510
rect 1822 14454 1878 14510
rect 1946 14454 2002 14510
rect 2070 14454 2126 14510
rect 1078 14330 1134 14386
rect 1202 14330 1258 14386
rect 1326 14330 1382 14386
rect 1450 14330 1506 14386
rect 1574 14330 1630 14386
rect 1698 14330 1754 14386
rect 1822 14330 1878 14386
rect 1946 14330 2002 14386
rect 2070 14330 2126 14386
rect 1078 14206 1134 14262
rect 1202 14206 1258 14262
rect 1326 14206 1382 14262
rect 1450 14206 1506 14262
rect 1574 14206 1630 14262
rect 1698 14206 1754 14262
rect 1822 14206 1878 14262
rect 1946 14206 2002 14262
rect 2070 14206 2126 14262
rect 1078 14082 1134 14138
rect 1202 14082 1258 14138
rect 1326 14082 1382 14138
rect 1450 14082 1506 14138
rect 1574 14082 1630 14138
rect 1698 14082 1754 14138
rect 1822 14082 1878 14138
rect 1946 14082 2002 14138
rect 2070 14082 2126 14138
rect 1078 13958 1134 14014
rect 1202 13958 1258 14014
rect 1326 13958 1382 14014
rect 1450 13958 1506 14014
rect 1574 13958 1630 14014
rect 1698 13958 1754 14014
rect 1822 13958 1878 14014
rect 1946 13958 2002 14014
rect 2070 13958 2126 14014
rect 1078 13834 1134 13890
rect 1202 13834 1258 13890
rect 1326 13834 1382 13890
rect 1450 13834 1506 13890
rect 1574 13834 1630 13890
rect 1698 13834 1754 13890
rect 1822 13834 1878 13890
rect 1946 13834 2002 13890
rect 2070 13834 2126 13890
rect 1078 13710 1134 13766
rect 1202 13710 1258 13766
rect 1326 13710 1382 13766
rect 1450 13710 1506 13766
rect 1574 13710 1630 13766
rect 1698 13710 1754 13766
rect 1822 13710 1878 13766
rect 1946 13710 2002 13766
rect 2070 13710 2126 13766
rect 1078 13586 1134 13642
rect 1202 13586 1258 13642
rect 1326 13586 1382 13642
rect 1450 13586 1506 13642
rect 1574 13586 1630 13642
rect 1698 13586 1754 13642
rect 1822 13586 1878 13642
rect 1946 13586 2002 13642
rect 2070 13586 2126 13642
rect 1078 13462 1134 13518
rect 1202 13462 1258 13518
rect 1326 13462 1382 13518
rect 1450 13462 1506 13518
rect 1574 13462 1630 13518
rect 1698 13462 1754 13518
rect 1822 13462 1878 13518
rect 1946 13462 2002 13518
rect 2070 13462 2126 13518
rect 1078 13338 1134 13394
rect 1202 13338 1258 13394
rect 1326 13338 1382 13394
rect 1450 13338 1506 13394
rect 1574 13338 1630 13394
rect 1698 13338 1754 13394
rect 1822 13338 1878 13394
rect 1946 13338 2002 13394
rect 2070 13338 2126 13394
rect 1078 13214 1134 13270
rect 1202 13214 1258 13270
rect 1326 13214 1382 13270
rect 1450 13214 1506 13270
rect 1574 13214 1630 13270
rect 1698 13214 1754 13270
rect 1822 13214 1878 13270
rect 1946 13214 2002 13270
rect 2070 13214 2126 13270
rect 1078 13090 1134 13146
rect 1202 13090 1258 13146
rect 1326 13090 1382 13146
rect 1450 13090 1506 13146
rect 1574 13090 1630 13146
rect 1698 13090 1754 13146
rect 1822 13090 1878 13146
rect 1946 13090 2002 13146
rect 2070 13090 2126 13146
rect 1078 12966 1134 13022
rect 1202 12966 1258 13022
rect 1326 12966 1382 13022
rect 1450 12966 1506 13022
rect 1574 12966 1630 13022
rect 1698 12966 1754 13022
rect 1822 12966 1878 13022
rect 1946 12966 2002 13022
rect 2070 12966 2126 13022
rect 1078 12842 1134 12898
rect 1202 12842 1258 12898
rect 1326 12842 1382 12898
rect 1450 12842 1506 12898
rect 1574 12842 1630 12898
rect 1698 12842 1754 12898
rect 1822 12842 1878 12898
rect 1946 12842 2002 12898
rect 2070 12842 2126 12898
rect 4435 15694 4491 15750
rect 4559 15694 4615 15750
rect 4683 15694 4739 15750
rect 4807 15694 4863 15750
rect 4931 15694 4987 15750
rect 5055 15694 5111 15750
rect 5179 15694 5235 15750
rect 5303 15694 5359 15750
rect 5427 15694 5483 15750
rect 5551 15694 5607 15750
rect 5675 15694 5731 15750
rect 5799 15694 5855 15750
rect 5923 15694 5979 15750
rect 6047 15694 6103 15750
rect 6171 15694 6227 15750
rect 4435 15570 4491 15626
rect 4559 15570 4615 15626
rect 4683 15570 4739 15626
rect 4807 15570 4863 15626
rect 4931 15570 4987 15626
rect 5055 15570 5111 15626
rect 5179 15570 5235 15626
rect 5303 15570 5359 15626
rect 5427 15570 5483 15626
rect 5551 15570 5607 15626
rect 5675 15570 5731 15626
rect 5799 15570 5855 15626
rect 5923 15570 5979 15626
rect 6047 15570 6103 15626
rect 6171 15570 6227 15626
rect 4435 15446 4491 15502
rect 4559 15446 4615 15502
rect 4683 15446 4739 15502
rect 4807 15446 4863 15502
rect 4931 15446 4987 15502
rect 5055 15446 5111 15502
rect 5179 15446 5235 15502
rect 5303 15446 5359 15502
rect 5427 15446 5483 15502
rect 5551 15446 5607 15502
rect 5675 15446 5731 15502
rect 5799 15446 5855 15502
rect 5923 15446 5979 15502
rect 6047 15446 6103 15502
rect 6171 15446 6227 15502
rect 4435 15322 4491 15378
rect 4559 15322 4615 15378
rect 4683 15322 4739 15378
rect 4807 15322 4863 15378
rect 4931 15322 4987 15378
rect 5055 15322 5111 15378
rect 5179 15322 5235 15378
rect 5303 15322 5359 15378
rect 5427 15322 5483 15378
rect 5551 15322 5607 15378
rect 5675 15322 5731 15378
rect 5799 15322 5855 15378
rect 5923 15322 5979 15378
rect 6047 15322 6103 15378
rect 6171 15322 6227 15378
rect 4435 15198 4491 15254
rect 4559 15198 4615 15254
rect 4683 15198 4739 15254
rect 4807 15198 4863 15254
rect 4931 15198 4987 15254
rect 5055 15198 5111 15254
rect 5179 15198 5235 15254
rect 5303 15198 5359 15254
rect 5427 15198 5483 15254
rect 5551 15198 5607 15254
rect 5675 15198 5731 15254
rect 5799 15198 5855 15254
rect 5923 15198 5979 15254
rect 6047 15198 6103 15254
rect 6171 15198 6227 15254
rect 4435 15074 4491 15130
rect 4559 15074 4615 15130
rect 4683 15074 4739 15130
rect 4807 15074 4863 15130
rect 4931 15074 4987 15130
rect 5055 15074 5111 15130
rect 5179 15074 5235 15130
rect 5303 15074 5359 15130
rect 5427 15074 5483 15130
rect 5551 15074 5607 15130
rect 5675 15074 5731 15130
rect 5799 15074 5855 15130
rect 5923 15074 5979 15130
rect 6047 15074 6103 15130
rect 6171 15074 6227 15130
rect 4435 14950 4491 15006
rect 4559 14950 4615 15006
rect 4683 14950 4739 15006
rect 4807 14950 4863 15006
rect 4931 14950 4987 15006
rect 5055 14950 5111 15006
rect 5179 14950 5235 15006
rect 5303 14950 5359 15006
rect 5427 14950 5483 15006
rect 5551 14950 5607 15006
rect 5675 14950 5731 15006
rect 5799 14950 5855 15006
rect 5923 14950 5979 15006
rect 6047 14950 6103 15006
rect 6171 14950 6227 15006
rect 4435 14826 4491 14882
rect 4559 14826 4615 14882
rect 4683 14826 4739 14882
rect 4807 14826 4863 14882
rect 4931 14826 4987 14882
rect 5055 14826 5111 14882
rect 5179 14826 5235 14882
rect 5303 14826 5359 14882
rect 5427 14826 5483 14882
rect 5551 14826 5607 14882
rect 5675 14826 5731 14882
rect 5799 14826 5855 14882
rect 5923 14826 5979 14882
rect 6047 14826 6103 14882
rect 6171 14826 6227 14882
rect 4435 14702 4491 14758
rect 4559 14702 4615 14758
rect 4683 14702 4739 14758
rect 4807 14702 4863 14758
rect 4931 14702 4987 14758
rect 5055 14702 5111 14758
rect 5179 14702 5235 14758
rect 5303 14702 5359 14758
rect 5427 14702 5483 14758
rect 5551 14702 5607 14758
rect 5675 14702 5731 14758
rect 5799 14702 5855 14758
rect 5923 14702 5979 14758
rect 6047 14702 6103 14758
rect 6171 14702 6227 14758
rect 4435 14578 4491 14634
rect 4559 14578 4615 14634
rect 4683 14578 4739 14634
rect 4807 14578 4863 14634
rect 4931 14578 4987 14634
rect 5055 14578 5111 14634
rect 5179 14578 5235 14634
rect 5303 14578 5359 14634
rect 5427 14578 5483 14634
rect 5551 14578 5607 14634
rect 5675 14578 5731 14634
rect 5799 14578 5855 14634
rect 5923 14578 5979 14634
rect 6047 14578 6103 14634
rect 6171 14578 6227 14634
rect 4435 14454 4491 14510
rect 4559 14454 4615 14510
rect 4683 14454 4739 14510
rect 4807 14454 4863 14510
rect 4931 14454 4987 14510
rect 5055 14454 5111 14510
rect 5179 14454 5235 14510
rect 5303 14454 5359 14510
rect 5427 14454 5483 14510
rect 5551 14454 5607 14510
rect 5675 14454 5731 14510
rect 5799 14454 5855 14510
rect 5923 14454 5979 14510
rect 6047 14454 6103 14510
rect 6171 14454 6227 14510
rect 4435 14330 4491 14386
rect 4559 14330 4615 14386
rect 4683 14330 4739 14386
rect 4807 14330 4863 14386
rect 4931 14330 4987 14386
rect 5055 14330 5111 14386
rect 5179 14330 5235 14386
rect 5303 14330 5359 14386
rect 5427 14330 5483 14386
rect 5551 14330 5607 14386
rect 5675 14330 5731 14386
rect 5799 14330 5855 14386
rect 5923 14330 5979 14386
rect 6047 14330 6103 14386
rect 6171 14330 6227 14386
rect 4435 14206 4491 14262
rect 4559 14206 4615 14262
rect 4683 14206 4739 14262
rect 4807 14206 4863 14262
rect 4931 14206 4987 14262
rect 5055 14206 5111 14262
rect 5179 14206 5235 14262
rect 5303 14206 5359 14262
rect 5427 14206 5483 14262
rect 5551 14206 5607 14262
rect 5675 14206 5731 14262
rect 5799 14206 5855 14262
rect 5923 14206 5979 14262
rect 6047 14206 6103 14262
rect 6171 14206 6227 14262
rect 4435 14082 4491 14138
rect 4559 14082 4615 14138
rect 4683 14082 4739 14138
rect 4807 14082 4863 14138
rect 4931 14082 4987 14138
rect 5055 14082 5111 14138
rect 5179 14082 5235 14138
rect 5303 14082 5359 14138
rect 5427 14082 5483 14138
rect 5551 14082 5607 14138
rect 5675 14082 5731 14138
rect 5799 14082 5855 14138
rect 5923 14082 5979 14138
rect 6047 14082 6103 14138
rect 6171 14082 6227 14138
rect 4435 13958 4491 14014
rect 4559 13958 4615 14014
rect 4683 13958 4739 14014
rect 4807 13958 4863 14014
rect 4931 13958 4987 14014
rect 5055 13958 5111 14014
rect 5179 13958 5235 14014
rect 5303 13958 5359 14014
rect 5427 13958 5483 14014
rect 5551 13958 5607 14014
rect 5675 13958 5731 14014
rect 5799 13958 5855 14014
rect 5923 13958 5979 14014
rect 6047 13958 6103 14014
rect 6171 13958 6227 14014
rect 4435 13834 4491 13890
rect 4559 13834 4615 13890
rect 4683 13834 4739 13890
rect 4807 13834 4863 13890
rect 4931 13834 4987 13890
rect 5055 13834 5111 13890
rect 5179 13834 5235 13890
rect 5303 13834 5359 13890
rect 5427 13834 5483 13890
rect 5551 13834 5607 13890
rect 5675 13834 5731 13890
rect 5799 13834 5855 13890
rect 5923 13834 5979 13890
rect 6047 13834 6103 13890
rect 6171 13834 6227 13890
rect 4435 13710 4491 13766
rect 4559 13710 4615 13766
rect 4683 13710 4739 13766
rect 4807 13710 4863 13766
rect 4931 13710 4987 13766
rect 5055 13710 5111 13766
rect 5179 13710 5235 13766
rect 5303 13710 5359 13766
rect 5427 13710 5483 13766
rect 5551 13710 5607 13766
rect 5675 13710 5731 13766
rect 5799 13710 5855 13766
rect 5923 13710 5979 13766
rect 6047 13710 6103 13766
rect 6171 13710 6227 13766
rect 4435 13586 4491 13642
rect 4559 13586 4615 13642
rect 4683 13586 4739 13642
rect 4807 13586 4863 13642
rect 4931 13586 4987 13642
rect 5055 13586 5111 13642
rect 5179 13586 5235 13642
rect 5303 13586 5359 13642
rect 5427 13586 5483 13642
rect 5551 13586 5607 13642
rect 5675 13586 5731 13642
rect 5799 13586 5855 13642
rect 5923 13586 5979 13642
rect 6047 13586 6103 13642
rect 6171 13586 6227 13642
rect 4435 13462 4491 13518
rect 4559 13462 4615 13518
rect 4683 13462 4739 13518
rect 4807 13462 4863 13518
rect 4931 13462 4987 13518
rect 5055 13462 5111 13518
rect 5179 13462 5235 13518
rect 5303 13462 5359 13518
rect 5427 13462 5483 13518
rect 5551 13462 5607 13518
rect 5675 13462 5731 13518
rect 5799 13462 5855 13518
rect 5923 13462 5979 13518
rect 6047 13462 6103 13518
rect 6171 13462 6227 13518
rect 4435 13338 4491 13394
rect 4559 13338 4615 13394
rect 4683 13338 4739 13394
rect 4807 13338 4863 13394
rect 4931 13338 4987 13394
rect 5055 13338 5111 13394
rect 5179 13338 5235 13394
rect 5303 13338 5359 13394
rect 5427 13338 5483 13394
rect 5551 13338 5607 13394
rect 5675 13338 5731 13394
rect 5799 13338 5855 13394
rect 5923 13338 5979 13394
rect 6047 13338 6103 13394
rect 6171 13338 6227 13394
rect 4435 13214 4491 13270
rect 4559 13214 4615 13270
rect 4683 13214 4739 13270
rect 4807 13214 4863 13270
rect 4931 13214 4987 13270
rect 5055 13214 5111 13270
rect 5179 13214 5235 13270
rect 5303 13214 5359 13270
rect 5427 13214 5483 13270
rect 5551 13214 5607 13270
rect 5675 13214 5731 13270
rect 5799 13214 5855 13270
rect 5923 13214 5979 13270
rect 6047 13214 6103 13270
rect 6171 13214 6227 13270
rect 4435 13090 4491 13146
rect 4559 13090 4615 13146
rect 4683 13090 4739 13146
rect 4807 13090 4863 13146
rect 4931 13090 4987 13146
rect 5055 13090 5111 13146
rect 5179 13090 5235 13146
rect 5303 13090 5359 13146
rect 5427 13090 5483 13146
rect 5551 13090 5607 13146
rect 5675 13090 5731 13146
rect 5799 13090 5855 13146
rect 5923 13090 5979 13146
rect 6047 13090 6103 13146
rect 6171 13090 6227 13146
rect 4435 12966 4491 13022
rect 4559 12966 4615 13022
rect 4683 12966 4739 13022
rect 4807 12966 4863 13022
rect 4931 12966 4987 13022
rect 5055 12966 5111 13022
rect 5179 12966 5235 13022
rect 5303 12966 5359 13022
rect 5427 12966 5483 13022
rect 5551 12966 5607 13022
rect 5675 12966 5731 13022
rect 5799 12966 5855 13022
rect 5923 12966 5979 13022
rect 6047 12966 6103 13022
rect 6171 12966 6227 13022
rect 4435 12842 4491 12898
rect 4559 12842 4615 12898
rect 4683 12842 4739 12898
rect 4807 12842 4863 12898
rect 4931 12842 4987 12898
rect 5055 12842 5111 12898
rect 5179 12842 5235 12898
rect 5303 12842 5359 12898
rect 5427 12842 5483 12898
rect 5551 12842 5607 12898
rect 5675 12842 5731 12898
rect 5799 12842 5855 12898
rect 5923 12842 5979 12898
rect 6047 12842 6103 12898
rect 6171 12842 6227 12898
rect 7562 15694 7618 15750
rect 7686 15694 7742 15750
rect 7810 15694 7866 15750
rect 7934 15694 7990 15750
rect 8058 15694 8114 15750
rect 8182 15694 8238 15750
rect 8306 15694 8362 15750
rect 8430 15694 8486 15750
rect 8554 15694 8610 15750
rect 7562 15570 7618 15626
rect 7686 15570 7742 15626
rect 7810 15570 7866 15626
rect 7934 15570 7990 15626
rect 8058 15570 8114 15626
rect 8182 15570 8238 15626
rect 8306 15570 8362 15626
rect 8430 15570 8486 15626
rect 8554 15570 8610 15626
rect 7562 15446 7618 15502
rect 7686 15446 7742 15502
rect 7810 15446 7866 15502
rect 7934 15446 7990 15502
rect 8058 15446 8114 15502
rect 8182 15446 8238 15502
rect 8306 15446 8362 15502
rect 8430 15446 8486 15502
rect 8554 15446 8610 15502
rect 7562 15322 7618 15378
rect 7686 15322 7742 15378
rect 7810 15322 7866 15378
rect 7934 15322 7990 15378
rect 8058 15322 8114 15378
rect 8182 15322 8238 15378
rect 8306 15322 8362 15378
rect 8430 15322 8486 15378
rect 8554 15322 8610 15378
rect 7562 15198 7618 15254
rect 7686 15198 7742 15254
rect 7810 15198 7866 15254
rect 7934 15198 7990 15254
rect 8058 15198 8114 15254
rect 8182 15198 8238 15254
rect 8306 15198 8362 15254
rect 8430 15198 8486 15254
rect 8554 15198 8610 15254
rect 7562 15074 7618 15130
rect 7686 15074 7742 15130
rect 7810 15074 7866 15130
rect 7934 15074 7990 15130
rect 8058 15074 8114 15130
rect 8182 15074 8238 15130
rect 8306 15074 8362 15130
rect 8430 15074 8486 15130
rect 8554 15074 8610 15130
rect 7562 14950 7618 15006
rect 7686 14950 7742 15006
rect 7810 14950 7866 15006
rect 7934 14950 7990 15006
rect 8058 14950 8114 15006
rect 8182 14950 8238 15006
rect 8306 14950 8362 15006
rect 8430 14950 8486 15006
rect 8554 14950 8610 15006
rect 7562 14826 7618 14882
rect 7686 14826 7742 14882
rect 7810 14826 7866 14882
rect 7934 14826 7990 14882
rect 8058 14826 8114 14882
rect 8182 14826 8238 14882
rect 8306 14826 8362 14882
rect 8430 14826 8486 14882
rect 8554 14826 8610 14882
rect 7562 14702 7618 14758
rect 7686 14702 7742 14758
rect 7810 14702 7866 14758
rect 7934 14702 7990 14758
rect 8058 14702 8114 14758
rect 8182 14702 8238 14758
rect 8306 14702 8362 14758
rect 8430 14702 8486 14758
rect 8554 14702 8610 14758
rect 7562 14578 7618 14634
rect 7686 14578 7742 14634
rect 7810 14578 7866 14634
rect 7934 14578 7990 14634
rect 8058 14578 8114 14634
rect 8182 14578 8238 14634
rect 8306 14578 8362 14634
rect 8430 14578 8486 14634
rect 8554 14578 8610 14634
rect 7562 14454 7618 14510
rect 7686 14454 7742 14510
rect 7810 14454 7866 14510
rect 7934 14454 7990 14510
rect 8058 14454 8114 14510
rect 8182 14454 8238 14510
rect 8306 14454 8362 14510
rect 8430 14454 8486 14510
rect 8554 14454 8610 14510
rect 7562 14330 7618 14386
rect 7686 14330 7742 14386
rect 7810 14330 7866 14386
rect 7934 14330 7990 14386
rect 8058 14330 8114 14386
rect 8182 14330 8238 14386
rect 8306 14330 8362 14386
rect 8430 14330 8486 14386
rect 8554 14330 8610 14386
rect 7562 14206 7618 14262
rect 7686 14206 7742 14262
rect 7810 14206 7866 14262
rect 7934 14206 7990 14262
rect 8058 14206 8114 14262
rect 8182 14206 8238 14262
rect 8306 14206 8362 14262
rect 8430 14206 8486 14262
rect 8554 14206 8610 14262
rect 7562 14082 7618 14138
rect 7686 14082 7742 14138
rect 7810 14082 7866 14138
rect 7934 14082 7990 14138
rect 8058 14082 8114 14138
rect 8182 14082 8238 14138
rect 8306 14082 8362 14138
rect 8430 14082 8486 14138
rect 8554 14082 8610 14138
rect 7562 13958 7618 14014
rect 7686 13958 7742 14014
rect 7810 13958 7866 14014
rect 7934 13958 7990 14014
rect 8058 13958 8114 14014
rect 8182 13958 8238 14014
rect 8306 13958 8362 14014
rect 8430 13958 8486 14014
rect 8554 13958 8610 14014
rect 7562 13834 7618 13890
rect 7686 13834 7742 13890
rect 7810 13834 7866 13890
rect 7934 13834 7990 13890
rect 8058 13834 8114 13890
rect 8182 13834 8238 13890
rect 8306 13834 8362 13890
rect 8430 13834 8486 13890
rect 8554 13834 8610 13890
rect 7562 13710 7618 13766
rect 7686 13710 7742 13766
rect 7810 13710 7866 13766
rect 7934 13710 7990 13766
rect 8058 13710 8114 13766
rect 8182 13710 8238 13766
rect 8306 13710 8362 13766
rect 8430 13710 8486 13766
rect 8554 13710 8610 13766
rect 7562 13586 7618 13642
rect 7686 13586 7742 13642
rect 7810 13586 7866 13642
rect 7934 13586 7990 13642
rect 8058 13586 8114 13642
rect 8182 13586 8238 13642
rect 8306 13586 8362 13642
rect 8430 13586 8486 13642
rect 8554 13586 8610 13642
rect 7562 13462 7618 13518
rect 7686 13462 7742 13518
rect 7810 13462 7866 13518
rect 7934 13462 7990 13518
rect 8058 13462 8114 13518
rect 8182 13462 8238 13518
rect 8306 13462 8362 13518
rect 8430 13462 8486 13518
rect 8554 13462 8610 13518
rect 7562 13338 7618 13394
rect 7686 13338 7742 13394
rect 7810 13338 7866 13394
rect 7934 13338 7990 13394
rect 8058 13338 8114 13394
rect 8182 13338 8238 13394
rect 8306 13338 8362 13394
rect 8430 13338 8486 13394
rect 8554 13338 8610 13394
rect 7562 13214 7618 13270
rect 7686 13214 7742 13270
rect 7810 13214 7866 13270
rect 7934 13214 7990 13270
rect 8058 13214 8114 13270
rect 8182 13214 8238 13270
rect 8306 13214 8362 13270
rect 8430 13214 8486 13270
rect 8554 13214 8610 13270
rect 7562 13090 7618 13146
rect 7686 13090 7742 13146
rect 7810 13090 7866 13146
rect 7934 13090 7990 13146
rect 8058 13090 8114 13146
rect 8182 13090 8238 13146
rect 8306 13090 8362 13146
rect 8430 13090 8486 13146
rect 8554 13090 8610 13146
rect 7562 12966 7618 13022
rect 7686 12966 7742 13022
rect 7810 12966 7866 13022
rect 7934 12966 7990 13022
rect 8058 12966 8114 13022
rect 8182 12966 8238 13022
rect 8306 12966 8362 13022
rect 8430 12966 8486 13022
rect 8554 12966 8610 13022
rect 7562 12842 7618 12898
rect 7686 12842 7742 12898
rect 7810 12842 7866 12898
rect 7934 12842 7990 12898
rect 8058 12842 8114 12898
rect 8182 12842 8238 12898
rect 8306 12842 8362 12898
rect 8430 12842 8486 12898
rect 8554 12842 8610 12898
rect 10679 15694 10735 15750
rect 10803 15694 10859 15750
rect 10927 15694 10983 15750
rect 11051 15694 11107 15750
rect 11175 15694 11231 15750
rect 11299 15694 11355 15750
rect 11423 15694 11479 15750
rect 11547 15694 11603 15750
rect 11671 15694 11727 15750
rect 11795 15694 11851 15750
rect 11919 15694 11975 15750
rect 12043 15694 12099 15750
rect 12167 15694 12223 15750
rect 12291 15694 12347 15750
rect 12415 15694 12471 15750
rect 10679 15570 10735 15626
rect 10803 15570 10859 15626
rect 10927 15570 10983 15626
rect 11051 15570 11107 15626
rect 11175 15570 11231 15626
rect 11299 15570 11355 15626
rect 11423 15570 11479 15626
rect 11547 15570 11603 15626
rect 11671 15570 11727 15626
rect 11795 15570 11851 15626
rect 11919 15570 11975 15626
rect 12043 15570 12099 15626
rect 12167 15570 12223 15626
rect 12291 15570 12347 15626
rect 12415 15570 12471 15626
rect 10679 15446 10735 15502
rect 10803 15446 10859 15502
rect 10927 15446 10983 15502
rect 11051 15446 11107 15502
rect 11175 15446 11231 15502
rect 11299 15446 11355 15502
rect 11423 15446 11479 15502
rect 11547 15446 11603 15502
rect 11671 15446 11727 15502
rect 11795 15446 11851 15502
rect 11919 15446 11975 15502
rect 12043 15446 12099 15502
rect 12167 15446 12223 15502
rect 12291 15446 12347 15502
rect 12415 15446 12471 15502
rect 10679 15322 10735 15378
rect 10803 15322 10859 15378
rect 10927 15322 10983 15378
rect 11051 15322 11107 15378
rect 11175 15322 11231 15378
rect 11299 15322 11355 15378
rect 11423 15322 11479 15378
rect 11547 15322 11603 15378
rect 11671 15322 11727 15378
rect 11795 15322 11851 15378
rect 11919 15322 11975 15378
rect 12043 15322 12099 15378
rect 12167 15322 12223 15378
rect 12291 15322 12347 15378
rect 12415 15322 12471 15378
rect 10679 15198 10735 15254
rect 10803 15198 10859 15254
rect 10927 15198 10983 15254
rect 11051 15198 11107 15254
rect 11175 15198 11231 15254
rect 11299 15198 11355 15254
rect 11423 15198 11479 15254
rect 11547 15198 11603 15254
rect 11671 15198 11727 15254
rect 11795 15198 11851 15254
rect 11919 15198 11975 15254
rect 12043 15198 12099 15254
rect 12167 15198 12223 15254
rect 12291 15198 12347 15254
rect 12415 15198 12471 15254
rect 10679 15074 10735 15130
rect 10803 15074 10859 15130
rect 10927 15074 10983 15130
rect 11051 15074 11107 15130
rect 11175 15074 11231 15130
rect 11299 15074 11355 15130
rect 11423 15074 11479 15130
rect 11547 15074 11603 15130
rect 11671 15074 11727 15130
rect 11795 15074 11851 15130
rect 11919 15074 11975 15130
rect 12043 15074 12099 15130
rect 12167 15074 12223 15130
rect 12291 15074 12347 15130
rect 12415 15074 12471 15130
rect 10679 14950 10735 15006
rect 10803 14950 10859 15006
rect 10927 14950 10983 15006
rect 11051 14950 11107 15006
rect 11175 14950 11231 15006
rect 11299 14950 11355 15006
rect 11423 14950 11479 15006
rect 11547 14950 11603 15006
rect 11671 14950 11727 15006
rect 11795 14950 11851 15006
rect 11919 14950 11975 15006
rect 12043 14950 12099 15006
rect 12167 14950 12223 15006
rect 12291 14950 12347 15006
rect 12415 14950 12471 15006
rect 10679 14826 10735 14882
rect 10803 14826 10859 14882
rect 10927 14826 10983 14882
rect 11051 14826 11107 14882
rect 11175 14826 11231 14882
rect 11299 14826 11355 14882
rect 11423 14826 11479 14882
rect 11547 14826 11603 14882
rect 11671 14826 11727 14882
rect 11795 14826 11851 14882
rect 11919 14826 11975 14882
rect 12043 14826 12099 14882
rect 12167 14826 12223 14882
rect 12291 14826 12347 14882
rect 12415 14826 12471 14882
rect 10679 14702 10735 14758
rect 10803 14702 10859 14758
rect 10927 14702 10983 14758
rect 11051 14702 11107 14758
rect 11175 14702 11231 14758
rect 11299 14702 11355 14758
rect 11423 14702 11479 14758
rect 11547 14702 11603 14758
rect 11671 14702 11727 14758
rect 11795 14702 11851 14758
rect 11919 14702 11975 14758
rect 12043 14702 12099 14758
rect 12167 14702 12223 14758
rect 12291 14702 12347 14758
rect 12415 14702 12471 14758
rect 10679 14578 10735 14634
rect 10803 14578 10859 14634
rect 10927 14578 10983 14634
rect 11051 14578 11107 14634
rect 11175 14578 11231 14634
rect 11299 14578 11355 14634
rect 11423 14578 11479 14634
rect 11547 14578 11603 14634
rect 11671 14578 11727 14634
rect 11795 14578 11851 14634
rect 11919 14578 11975 14634
rect 12043 14578 12099 14634
rect 12167 14578 12223 14634
rect 12291 14578 12347 14634
rect 12415 14578 12471 14634
rect 10679 14454 10735 14510
rect 10803 14454 10859 14510
rect 10927 14454 10983 14510
rect 11051 14454 11107 14510
rect 11175 14454 11231 14510
rect 11299 14454 11355 14510
rect 11423 14454 11479 14510
rect 11547 14454 11603 14510
rect 11671 14454 11727 14510
rect 11795 14454 11851 14510
rect 11919 14454 11975 14510
rect 12043 14454 12099 14510
rect 12167 14454 12223 14510
rect 12291 14454 12347 14510
rect 12415 14454 12471 14510
rect 10679 14330 10735 14386
rect 10803 14330 10859 14386
rect 10927 14330 10983 14386
rect 11051 14330 11107 14386
rect 11175 14330 11231 14386
rect 11299 14330 11355 14386
rect 11423 14330 11479 14386
rect 11547 14330 11603 14386
rect 11671 14330 11727 14386
rect 11795 14330 11851 14386
rect 11919 14330 11975 14386
rect 12043 14330 12099 14386
rect 12167 14330 12223 14386
rect 12291 14330 12347 14386
rect 12415 14330 12471 14386
rect 10679 14206 10735 14262
rect 10803 14206 10859 14262
rect 10927 14206 10983 14262
rect 11051 14206 11107 14262
rect 11175 14206 11231 14262
rect 11299 14206 11355 14262
rect 11423 14206 11479 14262
rect 11547 14206 11603 14262
rect 11671 14206 11727 14262
rect 11795 14206 11851 14262
rect 11919 14206 11975 14262
rect 12043 14206 12099 14262
rect 12167 14206 12223 14262
rect 12291 14206 12347 14262
rect 12415 14206 12471 14262
rect 10679 14082 10735 14138
rect 10803 14082 10859 14138
rect 10927 14082 10983 14138
rect 11051 14082 11107 14138
rect 11175 14082 11231 14138
rect 11299 14082 11355 14138
rect 11423 14082 11479 14138
rect 11547 14082 11603 14138
rect 11671 14082 11727 14138
rect 11795 14082 11851 14138
rect 11919 14082 11975 14138
rect 12043 14082 12099 14138
rect 12167 14082 12223 14138
rect 12291 14082 12347 14138
rect 12415 14082 12471 14138
rect 10679 13958 10735 14014
rect 10803 13958 10859 14014
rect 10927 13958 10983 14014
rect 11051 13958 11107 14014
rect 11175 13958 11231 14014
rect 11299 13958 11355 14014
rect 11423 13958 11479 14014
rect 11547 13958 11603 14014
rect 11671 13958 11727 14014
rect 11795 13958 11851 14014
rect 11919 13958 11975 14014
rect 12043 13958 12099 14014
rect 12167 13958 12223 14014
rect 12291 13958 12347 14014
rect 12415 13958 12471 14014
rect 10679 13834 10735 13890
rect 10803 13834 10859 13890
rect 10927 13834 10983 13890
rect 11051 13834 11107 13890
rect 11175 13834 11231 13890
rect 11299 13834 11355 13890
rect 11423 13834 11479 13890
rect 11547 13834 11603 13890
rect 11671 13834 11727 13890
rect 11795 13834 11851 13890
rect 11919 13834 11975 13890
rect 12043 13834 12099 13890
rect 12167 13834 12223 13890
rect 12291 13834 12347 13890
rect 12415 13834 12471 13890
rect 10679 13710 10735 13766
rect 10803 13710 10859 13766
rect 10927 13710 10983 13766
rect 11051 13710 11107 13766
rect 11175 13710 11231 13766
rect 11299 13710 11355 13766
rect 11423 13710 11479 13766
rect 11547 13710 11603 13766
rect 11671 13710 11727 13766
rect 11795 13710 11851 13766
rect 11919 13710 11975 13766
rect 12043 13710 12099 13766
rect 12167 13710 12223 13766
rect 12291 13710 12347 13766
rect 12415 13710 12471 13766
rect 10679 13586 10735 13642
rect 10803 13586 10859 13642
rect 10927 13586 10983 13642
rect 11051 13586 11107 13642
rect 11175 13586 11231 13642
rect 11299 13586 11355 13642
rect 11423 13586 11479 13642
rect 11547 13586 11603 13642
rect 11671 13586 11727 13642
rect 11795 13586 11851 13642
rect 11919 13586 11975 13642
rect 12043 13586 12099 13642
rect 12167 13586 12223 13642
rect 12291 13586 12347 13642
rect 12415 13586 12471 13642
rect 10679 13462 10735 13518
rect 10803 13462 10859 13518
rect 10927 13462 10983 13518
rect 11051 13462 11107 13518
rect 11175 13462 11231 13518
rect 11299 13462 11355 13518
rect 11423 13462 11479 13518
rect 11547 13462 11603 13518
rect 11671 13462 11727 13518
rect 11795 13462 11851 13518
rect 11919 13462 11975 13518
rect 12043 13462 12099 13518
rect 12167 13462 12223 13518
rect 12291 13462 12347 13518
rect 12415 13462 12471 13518
rect 10679 13338 10735 13394
rect 10803 13338 10859 13394
rect 10927 13338 10983 13394
rect 11051 13338 11107 13394
rect 11175 13338 11231 13394
rect 11299 13338 11355 13394
rect 11423 13338 11479 13394
rect 11547 13338 11603 13394
rect 11671 13338 11727 13394
rect 11795 13338 11851 13394
rect 11919 13338 11975 13394
rect 12043 13338 12099 13394
rect 12167 13338 12223 13394
rect 12291 13338 12347 13394
rect 12415 13338 12471 13394
rect 10679 13214 10735 13270
rect 10803 13214 10859 13270
rect 10927 13214 10983 13270
rect 11051 13214 11107 13270
rect 11175 13214 11231 13270
rect 11299 13214 11355 13270
rect 11423 13214 11479 13270
rect 11547 13214 11603 13270
rect 11671 13214 11727 13270
rect 11795 13214 11851 13270
rect 11919 13214 11975 13270
rect 12043 13214 12099 13270
rect 12167 13214 12223 13270
rect 12291 13214 12347 13270
rect 12415 13214 12471 13270
rect 10679 13090 10735 13146
rect 10803 13090 10859 13146
rect 10927 13090 10983 13146
rect 11051 13090 11107 13146
rect 11175 13090 11231 13146
rect 11299 13090 11355 13146
rect 11423 13090 11479 13146
rect 11547 13090 11603 13146
rect 11671 13090 11727 13146
rect 11795 13090 11851 13146
rect 11919 13090 11975 13146
rect 12043 13090 12099 13146
rect 12167 13090 12223 13146
rect 12291 13090 12347 13146
rect 12415 13090 12471 13146
rect 10679 12966 10735 13022
rect 10803 12966 10859 13022
rect 10927 12966 10983 13022
rect 11051 12966 11107 13022
rect 11175 12966 11231 13022
rect 11299 12966 11355 13022
rect 11423 12966 11479 13022
rect 11547 12966 11603 13022
rect 11671 12966 11727 13022
rect 11795 12966 11851 13022
rect 11919 12966 11975 13022
rect 12043 12966 12099 13022
rect 12167 12966 12223 13022
rect 12291 12966 12347 13022
rect 12415 12966 12471 13022
rect 10679 12842 10735 12898
rect 10803 12842 10859 12898
rect 10927 12842 10983 12898
rect 11051 12842 11107 12898
rect 11175 12842 11231 12898
rect 11299 12842 11355 12898
rect 11423 12842 11479 12898
rect 11547 12842 11603 12898
rect 11671 12842 11727 12898
rect 11795 12842 11851 12898
rect 11919 12842 11975 12898
rect 12043 12842 12099 12898
rect 12167 12842 12223 12898
rect 12291 12842 12347 12898
rect 12415 12842 12471 12898
rect 2507 12488 2563 12544
rect 2631 12488 2687 12544
rect 2755 12488 2811 12544
rect 2879 12488 2935 12544
rect 3003 12488 3059 12544
rect 3127 12488 3183 12544
rect 3251 12488 3307 12544
rect 3375 12488 3431 12544
rect 3499 12488 3555 12544
rect 3623 12488 3679 12544
rect 3747 12488 3803 12544
rect 3871 12488 3927 12544
rect 3995 12488 4051 12544
rect 4119 12488 4175 12544
rect 4243 12488 4299 12544
rect 2507 12364 2563 12420
rect 2631 12364 2687 12420
rect 2755 12364 2811 12420
rect 2879 12364 2935 12420
rect 3003 12364 3059 12420
rect 3127 12364 3183 12420
rect 3251 12364 3307 12420
rect 3375 12364 3431 12420
rect 3499 12364 3555 12420
rect 3623 12364 3679 12420
rect 3747 12364 3803 12420
rect 3871 12364 3927 12420
rect 3995 12364 4051 12420
rect 4119 12364 4175 12420
rect 4243 12364 4299 12420
rect 2507 12240 2563 12296
rect 2631 12240 2687 12296
rect 2755 12240 2811 12296
rect 2879 12240 2935 12296
rect 3003 12240 3059 12296
rect 3127 12240 3183 12296
rect 3251 12240 3307 12296
rect 3375 12240 3431 12296
rect 3499 12240 3555 12296
rect 3623 12240 3679 12296
rect 3747 12240 3803 12296
rect 3871 12240 3927 12296
rect 3995 12240 4051 12296
rect 4119 12240 4175 12296
rect 4243 12240 4299 12296
rect 2507 12116 2563 12172
rect 2631 12116 2687 12172
rect 2755 12116 2811 12172
rect 2879 12116 2935 12172
rect 3003 12116 3059 12172
rect 3127 12116 3183 12172
rect 3251 12116 3307 12172
rect 3375 12116 3431 12172
rect 3499 12116 3555 12172
rect 3623 12116 3679 12172
rect 3747 12116 3803 12172
rect 3871 12116 3927 12172
rect 3995 12116 4051 12172
rect 4119 12116 4175 12172
rect 4243 12116 4299 12172
rect 2507 11992 2563 12048
rect 2631 11992 2687 12048
rect 2755 11992 2811 12048
rect 2879 11992 2935 12048
rect 3003 11992 3059 12048
rect 3127 11992 3183 12048
rect 3251 11992 3307 12048
rect 3375 11992 3431 12048
rect 3499 11992 3555 12048
rect 3623 11992 3679 12048
rect 3747 11992 3803 12048
rect 3871 11992 3927 12048
rect 3995 11992 4051 12048
rect 4119 11992 4175 12048
rect 4243 11992 4299 12048
rect 2507 11868 2563 11924
rect 2631 11868 2687 11924
rect 2755 11868 2811 11924
rect 2879 11868 2935 11924
rect 3003 11868 3059 11924
rect 3127 11868 3183 11924
rect 3251 11868 3307 11924
rect 3375 11868 3431 11924
rect 3499 11868 3555 11924
rect 3623 11868 3679 11924
rect 3747 11868 3803 11924
rect 3871 11868 3927 11924
rect 3995 11868 4051 11924
rect 4119 11868 4175 11924
rect 4243 11868 4299 11924
rect 2507 11744 2563 11800
rect 2631 11744 2687 11800
rect 2755 11744 2811 11800
rect 2879 11744 2935 11800
rect 3003 11744 3059 11800
rect 3127 11744 3183 11800
rect 3251 11744 3307 11800
rect 3375 11744 3431 11800
rect 3499 11744 3555 11800
rect 3623 11744 3679 11800
rect 3747 11744 3803 11800
rect 3871 11744 3927 11800
rect 3995 11744 4051 11800
rect 4119 11744 4175 11800
rect 4243 11744 4299 11800
rect 2507 11620 2563 11676
rect 2631 11620 2687 11676
rect 2755 11620 2811 11676
rect 2879 11620 2935 11676
rect 3003 11620 3059 11676
rect 3127 11620 3183 11676
rect 3251 11620 3307 11676
rect 3375 11620 3431 11676
rect 3499 11620 3555 11676
rect 3623 11620 3679 11676
rect 3747 11620 3803 11676
rect 3871 11620 3927 11676
rect 3995 11620 4051 11676
rect 4119 11620 4175 11676
rect 4243 11620 4299 11676
rect 2507 11496 2563 11552
rect 2631 11496 2687 11552
rect 2755 11496 2811 11552
rect 2879 11496 2935 11552
rect 3003 11496 3059 11552
rect 3127 11496 3183 11552
rect 3251 11496 3307 11552
rect 3375 11496 3431 11552
rect 3499 11496 3555 11552
rect 3623 11496 3679 11552
rect 3747 11496 3803 11552
rect 3871 11496 3927 11552
rect 3995 11496 4051 11552
rect 4119 11496 4175 11552
rect 4243 11496 4299 11552
rect 2507 11372 2563 11428
rect 2631 11372 2687 11428
rect 2755 11372 2811 11428
rect 2879 11372 2935 11428
rect 3003 11372 3059 11428
rect 3127 11372 3183 11428
rect 3251 11372 3307 11428
rect 3375 11372 3431 11428
rect 3499 11372 3555 11428
rect 3623 11372 3679 11428
rect 3747 11372 3803 11428
rect 3871 11372 3927 11428
rect 3995 11372 4051 11428
rect 4119 11372 4175 11428
rect 4243 11372 4299 11428
rect 2507 11248 2563 11304
rect 2631 11248 2687 11304
rect 2755 11248 2811 11304
rect 2879 11248 2935 11304
rect 3003 11248 3059 11304
rect 3127 11248 3183 11304
rect 3251 11248 3307 11304
rect 3375 11248 3431 11304
rect 3499 11248 3555 11304
rect 3623 11248 3679 11304
rect 3747 11248 3803 11304
rect 3871 11248 3927 11304
rect 3995 11248 4051 11304
rect 4119 11248 4175 11304
rect 4243 11248 4299 11304
rect 6368 12488 6424 12544
rect 6492 12488 6548 12544
rect 6616 12488 6672 12544
rect 6740 12488 6796 12544
rect 6864 12488 6920 12544
rect 6988 12488 7044 12544
rect 7112 12488 7168 12544
rect 7236 12488 7292 12544
rect 7360 12488 7416 12544
rect 6368 12364 6424 12420
rect 6492 12364 6548 12420
rect 6616 12364 6672 12420
rect 6740 12364 6796 12420
rect 6864 12364 6920 12420
rect 6988 12364 7044 12420
rect 7112 12364 7168 12420
rect 7236 12364 7292 12420
rect 7360 12364 7416 12420
rect 6368 12240 6424 12296
rect 6492 12240 6548 12296
rect 6616 12240 6672 12296
rect 6740 12240 6796 12296
rect 6864 12240 6920 12296
rect 6988 12240 7044 12296
rect 7112 12240 7168 12296
rect 7236 12240 7292 12296
rect 7360 12240 7416 12296
rect 6368 12116 6424 12172
rect 6492 12116 6548 12172
rect 6616 12116 6672 12172
rect 6740 12116 6796 12172
rect 6864 12116 6920 12172
rect 6988 12116 7044 12172
rect 7112 12116 7168 12172
rect 7236 12116 7292 12172
rect 7360 12116 7416 12172
rect 6368 11992 6424 12048
rect 6492 11992 6548 12048
rect 6616 11992 6672 12048
rect 6740 11992 6796 12048
rect 6864 11992 6920 12048
rect 6988 11992 7044 12048
rect 7112 11992 7168 12048
rect 7236 11992 7292 12048
rect 7360 11992 7416 12048
rect 6368 11868 6424 11924
rect 6492 11868 6548 11924
rect 6616 11868 6672 11924
rect 6740 11868 6796 11924
rect 6864 11868 6920 11924
rect 6988 11868 7044 11924
rect 7112 11868 7168 11924
rect 7236 11868 7292 11924
rect 7360 11868 7416 11924
rect 6368 11744 6424 11800
rect 6492 11744 6548 11800
rect 6616 11744 6672 11800
rect 6740 11744 6796 11800
rect 6864 11744 6920 11800
rect 6988 11744 7044 11800
rect 7112 11744 7168 11800
rect 7236 11744 7292 11800
rect 7360 11744 7416 11800
rect 6368 11620 6424 11676
rect 6492 11620 6548 11676
rect 6616 11620 6672 11676
rect 6740 11620 6796 11676
rect 6864 11620 6920 11676
rect 6988 11620 7044 11676
rect 7112 11620 7168 11676
rect 7236 11620 7292 11676
rect 7360 11620 7416 11676
rect 6368 11496 6424 11552
rect 6492 11496 6548 11552
rect 6616 11496 6672 11552
rect 6740 11496 6796 11552
rect 6864 11496 6920 11552
rect 6988 11496 7044 11552
rect 7112 11496 7168 11552
rect 7236 11496 7292 11552
rect 7360 11496 7416 11552
rect 6368 11372 6424 11428
rect 6492 11372 6548 11428
rect 6616 11372 6672 11428
rect 6740 11372 6796 11428
rect 6864 11372 6920 11428
rect 6988 11372 7044 11428
rect 7112 11372 7168 11428
rect 7236 11372 7292 11428
rect 7360 11372 7416 11428
rect 6368 11248 6424 11304
rect 6492 11248 6548 11304
rect 6616 11248 6672 11304
rect 6740 11248 6796 11304
rect 6864 11248 6920 11304
rect 6988 11248 7044 11304
rect 7112 11248 7168 11304
rect 7236 11248 7292 11304
rect 7360 11248 7416 11304
rect 8751 12488 8807 12544
rect 8875 12488 8931 12544
rect 8999 12488 9055 12544
rect 9123 12488 9179 12544
rect 9247 12488 9303 12544
rect 9371 12488 9427 12544
rect 9495 12488 9551 12544
rect 9619 12488 9675 12544
rect 9743 12488 9799 12544
rect 9867 12488 9923 12544
rect 9991 12488 10047 12544
rect 10115 12488 10171 12544
rect 10239 12488 10295 12544
rect 10363 12488 10419 12544
rect 10487 12488 10543 12544
rect 8751 12364 8807 12420
rect 8875 12364 8931 12420
rect 8999 12364 9055 12420
rect 9123 12364 9179 12420
rect 9247 12364 9303 12420
rect 9371 12364 9427 12420
rect 9495 12364 9551 12420
rect 9619 12364 9675 12420
rect 9743 12364 9799 12420
rect 9867 12364 9923 12420
rect 9991 12364 10047 12420
rect 10115 12364 10171 12420
rect 10239 12364 10295 12420
rect 10363 12364 10419 12420
rect 10487 12364 10543 12420
rect 8751 12240 8807 12296
rect 8875 12240 8931 12296
rect 8999 12240 9055 12296
rect 9123 12240 9179 12296
rect 9247 12240 9303 12296
rect 9371 12240 9427 12296
rect 9495 12240 9551 12296
rect 9619 12240 9675 12296
rect 9743 12240 9799 12296
rect 9867 12240 9923 12296
rect 9991 12240 10047 12296
rect 10115 12240 10171 12296
rect 10239 12240 10295 12296
rect 10363 12240 10419 12296
rect 10487 12240 10543 12296
rect 8751 12116 8807 12172
rect 8875 12116 8931 12172
rect 8999 12116 9055 12172
rect 9123 12116 9179 12172
rect 9247 12116 9303 12172
rect 9371 12116 9427 12172
rect 9495 12116 9551 12172
rect 9619 12116 9675 12172
rect 9743 12116 9799 12172
rect 9867 12116 9923 12172
rect 9991 12116 10047 12172
rect 10115 12116 10171 12172
rect 10239 12116 10295 12172
rect 10363 12116 10419 12172
rect 10487 12116 10543 12172
rect 8751 11992 8807 12048
rect 8875 11992 8931 12048
rect 8999 11992 9055 12048
rect 9123 11992 9179 12048
rect 9247 11992 9303 12048
rect 9371 11992 9427 12048
rect 9495 11992 9551 12048
rect 9619 11992 9675 12048
rect 9743 11992 9799 12048
rect 9867 11992 9923 12048
rect 9991 11992 10047 12048
rect 10115 11992 10171 12048
rect 10239 11992 10295 12048
rect 10363 11992 10419 12048
rect 10487 11992 10543 12048
rect 8751 11868 8807 11924
rect 8875 11868 8931 11924
rect 8999 11868 9055 11924
rect 9123 11868 9179 11924
rect 9247 11868 9303 11924
rect 9371 11868 9427 11924
rect 9495 11868 9551 11924
rect 9619 11868 9675 11924
rect 9743 11868 9799 11924
rect 9867 11868 9923 11924
rect 9991 11868 10047 11924
rect 10115 11868 10171 11924
rect 10239 11868 10295 11924
rect 10363 11868 10419 11924
rect 10487 11868 10543 11924
rect 8751 11744 8807 11800
rect 8875 11744 8931 11800
rect 8999 11744 9055 11800
rect 9123 11744 9179 11800
rect 9247 11744 9303 11800
rect 9371 11744 9427 11800
rect 9495 11744 9551 11800
rect 9619 11744 9675 11800
rect 9743 11744 9799 11800
rect 9867 11744 9923 11800
rect 9991 11744 10047 11800
rect 10115 11744 10171 11800
rect 10239 11744 10295 11800
rect 10363 11744 10419 11800
rect 10487 11744 10543 11800
rect 8751 11620 8807 11676
rect 8875 11620 8931 11676
rect 8999 11620 9055 11676
rect 9123 11620 9179 11676
rect 9247 11620 9303 11676
rect 9371 11620 9427 11676
rect 9495 11620 9551 11676
rect 9619 11620 9675 11676
rect 9743 11620 9799 11676
rect 9867 11620 9923 11676
rect 9991 11620 10047 11676
rect 10115 11620 10171 11676
rect 10239 11620 10295 11676
rect 10363 11620 10419 11676
rect 10487 11620 10543 11676
rect 8751 11496 8807 11552
rect 8875 11496 8931 11552
rect 8999 11496 9055 11552
rect 9123 11496 9179 11552
rect 9247 11496 9303 11552
rect 9371 11496 9427 11552
rect 9495 11496 9551 11552
rect 9619 11496 9675 11552
rect 9743 11496 9799 11552
rect 9867 11496 9923 11552
rect 9991 11496 10047 11552
rect 10115 11496 10171 11552
rect 10239 11496 10295 11552
rect 10363 11496 10419 11552
rect 10487 11496 10543 11552
rect 8751 11372 8807 11428
rect 8875 11372 8931 11428
rect 8999 11372 9055 11428
rect 9123 11372 9179 11428
rect 9247 11372 9303 11428
rect 9371 11372 9427 11428
rect 9495 11372 9551 11428
rect 9619 11372 9675 11428
rect 9743 11372 9799 11428
rect 9867 11372 9923 11428
rect 9991 11372 10047 11428
rect 10115 11372 10171 11428
rect 10239 11372 10295 11428
rect 10363 11372 10419 11428
rect 10487 11372 10543 11428
rect 8751 11248 8807 11304
rect 8875 11248 8931 11304
rect 8999 11248 9055 11304
rect 9123 11248 9179 11304
rect 9247 11248 9303 11304
rect 9371 11248 9427 11304
rect 9495 11248 9551 11304
rect 9619 11248 9675 11304
rect 9743 11248 9799 11304
rect 9867 11248 9923 11304
rect 9991 11248 10047 11304
rect 10115 11248 10171 11304
rect 10239 11248 10295 11304
rect 10363 11248 10419 11304
rect 10487 11248 10543 11304
rect 12852 12488 12908 12544
rect 12976 12488 13032 12544
rect 13100 12488 13156 12544
rect 13224 12488 13280 12544
rect 13348 12488 13404 12544
rect 13472 12488 13528 12544
rect 13596 12488 13652 12544
rect 13720 12488 13776 12544
rect 13844 12488 13900 12544
rect 12852 12364 12908 12420
rect 12976 12364 13032 12420
rect 13100 12364 13156 12420
rect 13224 12364 13280 12420
rect 13348 12364 13404 12420
rect 13472 12364 13528 12420
rect 13596 12364 13652 12420
rect 13720 12364 13776 12420
rect 13844 12364 13900 12420
rect 12852 12240 12908 12296
rect 12976 12240 13032 12296
rect 13100 12240 13156 12296
rect 13224 12240 13280 12296
rect 13348 12240 13404 12296
rect 13472 12240 13528 12296
rect 13596 12240 13652 12296
rect 13720 12240 13776 12296
rect 13844 12240 13900 12296
rect 12852 12116 12908 12172
rect 12976 12116 13032 12172
rect 13100 12116 13156 12172
rect 13224 12116 13280 12172
rect 13348 12116 13404 12172
rect 13472 12116 13528 12172
rect 13596 12116 13652 12172
rect 13720 12116 13776 12172
rect 13844 12116 13900 12172
rect 12852 11992 12908 12048
rect 12976 11992 13032 12048
rect 13100 11992 13156 12048
rect 13224 11992 13280 12048
rect 13348 11992 13404 12048
rect 13472 11992 13528 12048
rect 13596 11992 13652 12048
rect 13720 11992 13776 12048
rect 13844 11992 13900 12048
rect 12852 11868 12908 11924
rect 12976 11868 13032 11924
rect 13100 11868 13156 11924
rect 13224 11868 13280 11924
rect 13348 11868 13404 11924
rect 13472 11868 13528 11924
rect 13596 11868 13652 11924
rect 13720 11868 13776 11924
rect 13844 11868 13900 11924
rect 12852 11744 12908 11800
rect 12976 11744 13032 11800
rect 13100 11744 13156 11800
rect 13224 11744 13280 11800
rect 13348 11744 13404 11800
rect 13472 11744 13528 11800
rect 13596 11744 13652 11800
rect 13720 11744 13776 11800
rect 13844 11744 13900 11800
rect 12852 11620 12908 11676
rect 12976 11620 13032 11676
rect 13100 11620 13156 11676
rect 13224 11620 13280 11676
rect 13348 11620 13404 11676
rect 13472 11620 13528 11676
rect 13596 11620 13652 11676
rect 13720 11620 13776 11676
rect 13844 11620 13900 11676
rect 12852 11496 12908 11552
rect 12976 11496 13032 11552
rect 13100 11496 13156 11552
rect 13224 11496 13280 11552
rect 13348 11496 13404 11552
rect 13472 11496 13528 11552
rect 13596 11496 13652 11552
rect 13720 11496 13776 11552
rect 13844 11496 13900 11552
rect 12852 11372 12908 11428
rect 12976 11372 13032 11428
rect 13100 11372 13156 11428
rect 13224 11372 13280 11428
rect 13348 11372 13404 11428
rect 13472 11372 13528 11428
rect 13596 11372 13652 11428
rect 13720 11372 13776 11428
rect 13844 11372 13900 11428
rect 12852 11248 12908 11304
rect 12976 11248 13032 11304
rect 13100 11248 13156 11304
rect 13224 11248 13280 11304
rect 13348 11248 13404 11304
rect 13472 11248 13528 11304
rect 13596 11248 13652 11304
rect 13720 11248 13776 11304
rect 13844 11248 13900 11304
rect 1078 10888 1134 10944
rect 1202 10888 1258 10944
rect 1326 10888 1382 10944
rect 1450 10888 1506 10944
rect 1574 10888 1630 10944
rect 1698 10888 1754 10944
rect 1822 10888 1878 10944
rect 1946 10888 2002 10944
rect 2070 10888 2126 10944
rect 1078 10764 1134 10820
rect 1202 10764 1258 10820
rect 1326 10764 1382 10820
rect 1450 10764 1506 10820
rect 1574 10764 1630 10820
rect 1698 10764 1754 10820
rect 1822 10764 1878 10820
rect 1946 10764 2002 10820
rect 2070 10764 2126 10820
rect 1078 10640 1134 10696
rect 1202 10640 1258 10696
rect 1326 10640 1382 10696
rect 1450 10640 1506 10696
rect 1574 10640 1630 10696
rect 1698 10640 1754 10696
rect 1822 10640 1878 10696
rect 1946 10640 2002 10696
rect 2070 10640 2126 10696
rect 1078 10516 1134 10572
rect 1202 10516 1258 10572
rect 1326 10516 1382 10572
rect 1450 10516 1506 10572
rect 1574 10516 1630 10572
rect 1698 10516 1754 10572
rect 1822 10516 1878 10572
rect 1946 10516 2002 10572
rect 2070 10516 2126 10572
rect 1078 10392 1134 10448
rect 1202 10392 1258 10448
rect 1326 10392 1382 10448
rect 1450 10392 1506 10448
rect 1574 10392 1630 10448
rect 1698 10392 1754 10448
rect 1822 10392 1878 10448
rect 1946 10392 2002 10448
rect 2070 10392 2126 10448
rect 1078 10268 1134 10324
rect 1202 10268 1258 10324
rect 1326 10268 1382 10324
rect 1450 10268 1506 10324
rect 1574 10268 1630 10324
rect 1698 10268 1754 10324
rect 1822 10268 1878 10324
rect 1946 10268 2002 10324
rect 2070 10268 2126 10324
rect 1078 10144 1134 10200
rect 1202 10144 1258 10200
rect 1326 10144 1382 10200
rect 1450 10144 1506 10200
rect 1574 10144 1630 10200
rect 1698 10144 1754 10200
rect 1822 10144 1878 10200
rect 1946 10144 2002 10200
rect 2070 10144 2126 10200
rect 1078 10020 1134 10076
rect 1202 10020 1258 10076
rect 1326 10020 1382 10076
rect 1450 10020 1506 10076
rect 1574 10020 1630 10076
rect 1698 10020 1754 10076
rect 1822 10020 1878 10076
rect 1946 10020 2002 10076
rect 2070 10020 2126 10076
rect 1078 9896 1134 9952
rect 1202 9896 1258 9952
rect 1326 9896 1382 9952
rect 1450 9896 1506 9952
rect 1574 9896 1630 9952
rect 1698 9896 1754 9952
rect 1822 9896 1878 9952
rect 1946 9896 2002 9952
rect 2070 9896 2126 9952
rect 1078 9772 1134 9828
rect 1202 9772 1258 9828
rect 1326 9772 1382 9828
rect 1450 9772 1506 9828
rect 1574 9772 1630 9828
rect 1698 9772 1754 9828
rect 1822 9772 1878 9828
rect 1946 9772 2002 9828
rect 2070 9772 2126 9828
rect 1078 9648 1134 9704
rect 1202 9648 1258 9704
rect 1326 9648 1382 9704
rect 1450 9648 1506 9704
rect 1574 9648 1630 9704
rect 1698 9648 1754 9704
rect 1822 9648 1878 9704
rect 1946 9648 2002 9704
rect 2070 9648 2126 9704
rect 4435 10888 4491 10944
rect 4559 10888 4615 10944
rect 4683 10888 4739 10944
rect 4807 10888 4863 10944
rect 4931 10888 4987 10944
rect 5055 10888 5111 10944
rect 5179 10888 5235 10944
rect 5303 10888 5359 10944
rect 5427 10888 5483 10944
rect 5551 10888 5607 10944
rect 5675 10888 5731 10944
rect 5799 10888 5855 10944
rect 5923 10888 5979 10944
rect 6047 10888 6103 10944
rect 6171 10888 6227 10944
rect 4435 10764 4491 10820
rect 4559 10764 4615 10820
rect 4683 10764 4739 10820
rect 4807 10764 4863 10820
rect 4931 10764 4987 10820
rect 5055 10764 5111 10820
rect 5179 10764 5235 10820
rect 5303 10764 5359 10820
rect 5427 10764 5483 10820
rect 5551 10764 5607 10820
rect 5675 10764 5731 10820
rect 5799 10764 5855 10820
rect 5923 10764 5979 10820
rect 6047 10764 6103 10820
rect 6171 10764 6227 10820
rect 4435 10640 4491 10696
rect 4559 10640 4615 10696
rect 4683 10640 4739 10696
rect 4807 10640 4863 10696
rect 4931 10640 4987 10696
rect 5055 10640 5111 10696
rect 5179 10640 5235 10696
rect 5303 10640 5359 10696
rect 5427 10640 5483 10696
rect 5551 10640 5607 10696
rect 5675 10640 5731 10696
rect 5799 10640 5855 10696
rect 5923 10640 5979 10696
rect 6047 10640 6103 10696
rect 6171 10640 6227 10696
rect 4435 10516 4491 10572
rect 4559 10516 4615 10572
rect 4683 10516 4739 10572
rect 4807 10516 4863 10572
rect 4931 10516 4987 10572
rect 5055 10516 5111 10572
rect 5179 10516 5235 10572
rect 5303 10516 5359 10572
rect 5427 10516 5483 10572
rect 5551 10516 5607 10572
rect 5675 10516 5731 10572
rect 5799 10516 5855 10572
rect 5923 10516 5979 10572
rect 6047 10516 6103 10572
rect 6171 10516 6227 10572
rect 4435 10392 4491 10448
rect 4559 10392 4615 10448
rect 4683 10392 4739 10448
rect 4807 10392 4863 10448
rect 4931 10392 4987 10448
rect 5055 10392 5111 10448
rect 5179 10392 5235 10448
rect 5303 10392 5359 10448
rect 5427 10392 5483 10448
rect 5551 10392 5607 10448
rect 5675 10392 5731 10448
rect 5799 10392 5855 10448
rect 5923 10392 5979 10448
rect 6047 10392 6103 10448
rect 6171 10392 6227 10448
rect 4435 10268 4491 10324
rect 4559 10268 4615 10324
rect 4683 10268 4739 10324
rect 4807 10268 4863 10324
rect 4931 10268 4987 10324
rect 5055 10268 5111 10324
rect 5179 10268 5235 10324
rect 5303 10268 5359 10324
rect 5427 10268 5483 10324
rect 5551 10268 5607 10324
rect 5675 10268 5731 10324
rect 5799 10268 5855 10324
rect 5923 10268 5979 10324
rect 6047 10268 6103 10324
rect 6171 10268 6227 10324
rect 4435 10144 4491 10200
rect 4559 10144 4615 10200
rect 4683 10144 4739 10200
rect 4807 10144 4863 10200
rect 4931 10144 4987 10200
rect 5055 10144 5111 10200
rect 5179 10144 5235 10200
rect 5303 10144 5359 10200
rect 5427 10144 5483 10200
rect 5551 10144 5607 10200
rect 5675 10144 5731 10200
rect 5799 10144 5855 10200
rect 5923 10144 5979 10200
rect 6047 10144 6103 10200
rect 6171 10144 6227 10200
rect 4435 10020 4491 10076
rect 4559 10020 4615 10076
rect 4683 10020 4739 10076
rect 4807 10020 4863 10076
rect 4931 10020 4987 10076
rect 5055 10020 5111 10076
rect 5179 10020 5235 10076
rect 5303 10020 5359 10076
rect 5427 10020 5483 10076
rect 5551 10020 5607 10076
rect 5675 10020 5731 10076
rect 5799 10020 5855 10076
rect 5923 10020 5979 10076
rect 6047 10020 6103 10076
rect 6171 10020 6227 10076
rect 4435 9896 4491 9952
rect 4559 9896 4615 9952
rect 4683 9896 4739 9952
rect 4807 9896 4863 9952
rect 4931 9896 4987 9952
rect 5055 9896 5111 9952
rect 5179 9896 5235 9952
rect 5303 9896 5359 9952
rect 5427 9896 5483 9952
rect 5551 9896 5607 9952
rect 5675 9896 5731 9952
rect 5799 9896 5855 9952
rect 5923 9896 5979 9952
rect 6047 9896 6103 9952
rect 6171 9896 6227 9952
rect 4435 9772 4491 9828
rect 4559 9772 4615 9828
rect 4683 9772 4739 9828
rect 4807 9772 4863 9828
rect 4931 9772 4987 9828
rect 5055 9772 5111 9828
rect 5179 9772 5235 9828
rect 5303 9772 5359 9828
rect 5427 9772 5483 9828
rect 5551 9772 5607 9828
rect 5675 9772 5731 9828
rect 5799 9772 5855 9828
rect 5923 9772 5979 9828
rect 6047 9772 6103 9828
rect 6171 9772 6227 9828
rect 4435 9648 4491 9704
rect 4559 9648 4615 9704
rect 4683 9648 4739 9704
rect 4807 9648 4863 9704
rect 4931 9648 4987 9704
rect 5055 9648 5111 9704
rect 5179 9648 5235 9704
rect 5303 9648 5359 9704
rect 5427 9648 5483 9704
rect 5551 9648 5607 9704
rect 5675 9648 5731 9704
rect 5799 9648 5855 9704
rect 5923 9648 5979 9704
rect 6047 9648 6103 9704
rect 6171 9648 6227 9704
rect 7562 10888 7618 10944
rect 7686 10888 7742 10944
rect 7810 10888 7866 10944
rect 7934 10888 7990 10944
rect 8058 10888 8114 10944
rect 8182 10888 8238 10944
rect 8306 10888 8362 10944
rect 8430 10888 8486 10944
rect 8554 10888 8610 10944
rect 7562 10764 7618 10820
rect 7686 10764 7742 10820
rect 7810 10764 7866 10820
rect 7934 10764 7990 10820
rect 8058 10764 8114 10820
rect 8182 10764 8238 10820
rect 8306 10764 8362 10820
rect 8430 10764 8486 10820
rect 8554 10764 8610 10820
rect 7562 10640 7618 10696
rect 7686 10640 7742 10696
rect 7810 10640 7866 10696
rect 7934 10640 7990 10696
rect 8058 10640 8114 10696
rect 8182 10640 8238 10696
rect 8306 10640 8362 10696
rect 8430 10640 8486 10696
rect 8554 10640 8610 10696
rect 7562 10516 7618 10572
rect 7686 10516 7742 10572
rect 7810 10516 7866 10572
rect 7934 10516 7990 10572
rect 8058 10516 8114 10572
rect 8182 10516 8238 10572
rect 8306 10516 8362 10572
rect 8430 10516 8486 10572
rect 8554 10516 8610 10572
rect 7562 10392 7618 10448
rect 7686 10392 7742 10448
rect 7810 10392 7866 10448
rect 7934 10392 7990 10448
rect 8058 10392 8114 10448
rect 8182 10392 8238 10448
rect 8306 10392 8362 10448
rect 8430 10392 8486 10448
rect 8554 10392 8610 10448
rect 7562 10268 7618 10324
rect 7686 10268 7742 10324
rect 7810 10268 7866 10324
rect 7934 10268 7990 10324
rect 8058 10268 8114 10324
rect 8182 10268 8238 10324
rect 8306 10268 8362 10324
rect 8430 10268 8486 10324
rect 8554 10268 8610 10324
rect 7562 10144 7618 10200
rect 7686 10144 7742 10200
rect 7810 10144 7866 10200
rect 7934 10144 7990 10200
rect 8058 10144 8114 10200
rect 8182 10144 8238 10200
rect 8306 10144 8362 10200
rect 8430 10144 8486 10200
rect 8554 10144 8610 10200
rect 7562 10020 7618 10076
rect 7686 10020 7742 10076
rect 7810 10020 7866 10076
rect 7934 10020 7990 10076
rect 8058 10020 8114 10076
rect 8182 10020 8238 10076
rect 8306 10020 8362 10076
rect 8430 10020 8486 10076
rect 8554 10020 8610 10076
rect 7562 9896 7618 9952
rect 7686 9896 7742 9952
rect 7810 9896 7866 9952
rect 7934 9896 7990 9952
rect 8058 9896 8114 9952
rect 8182 9896 8238 9952
rect 8306 9896 8362 9952
rect 8430 9896 8486 9952
rect 8554 9896 8610 9952
rect 7562 9772 7618 9828
rect 7686 9772 7742 9828
rect 7810 9772 7866 9828
rect 7934 9772 7990 9828
rect 8058 9772 8114 9828
rect 8182 9772 8238 9828
rect 8306 9772 8362 9828
rect 8430 9772 8486 9828
rect 8554 9772 8610 9828
rect 7562 9648 7618 9704
rect 7686 9648 7742 9704
rect 7810 9648 7866 9704
rect 7934 9648 7990 9704
rect 8058 9648 8114 9704
rect 8182 9648 8238 9704
rect 8306 9648 8362 9704
rect 8430 9648 8486 9704
rect 8554 9648 8610 9704
rect 10679 10888 10735 10944
rect 10803 10888 10859 10944
rect 10927 10888 10983 10944
rect 11051 10888 11107 10944
rect 11175 10888 11231 10944
rect 11299 10888 11355 10944
rect 11423 10888 11479 10944
rect 11547 10888 11603 10944
rect 11671 10888 11727 10944
rect 11795 10888 11851 10944
rect 11919 10888 11975 10944
rect 12043 10888 12099 10944
rect 12167 10888 12223 10944
rect 12291 10888 12347 10944
rect 12415 10888 12471 10944
rect 10679 10764 10735 10820
rect 10803 10764 10859 10820
rect 10927 10764 10983 10820
rect 11051 10764 11107 10820
rect 11175 10764 11231 10820
rect 11299 10764 11355 10820
rect 11423 10764 11479 10820
rect 11547 10764 11603 10820
rect 11671 10764 11727 10820
rect 11795 10764 11851 10820
rect 11919 10764 11975 10820
rect 12043 10764 12099 10820
rect 12167 10764 12223 10820
rect 12291 10764 12347 10820
rect 12415 10764 12471 10820
rect 10679 10640 10735 10696
rect 10803 10640 10859 10696
rect 10927 10640 10983 10696
rect 11051 10640 11107 10696
rect 11175 10640 11231 10696
rect 11299 10640 11355 10696
rect 11423 10640 11479 10696
rect 11547 10640 11603 10696
rect 11671 10640 11727 10696
rect 11795 10640 11851 10696
rect 11919 10640 11975 10696
rect 12043 10640 12099 10696
rect 12167 10640 12223 10696
rect 12291 10640 12347 10696
rect 12415 10640 12471 10696
rect 10679 10516 10735 10572
rect 10803 10516 10859 10572
rect 10927 10516 10983 10572
rect 11051 10516 11107 10572
rect 11175 10516 11231 10572
rect 11299 10516 11355 10572
rect 11423 10516 11479 10572
rect 11547 10516 11603 10572
rect 11671 10516 11727 10572
rect 11795 10516 11851 10572
rect 11919 10516 11975 10572
rect 12043 10516 12099 10572
rect 12167 10516 12223 10572
rect 12291 10516 12347 10572
rect 12415 10516 12471 10572
rect 10679 10392 10735 10448
rect 10803 10392 10859 10448
rect 10927 10392 10983 10448
rect 11051 10392 11107 10448
rect 11175 10392 11231 10448
rect 11299 10392 11355 10448
rect 11423 10392 11479 10448
rect 11547 10392 11603 10448
rect 11671 10392 11727 10448
rect 11795 10392 11851 10448
rect 11919 10392 11975 10448
rect 12043 10392 12099 10448
rect 12167 10392 12223 10448
rect 12291 10392 12347 10448
rect 12415 10392 12471 10448
rect 10679 10268 10735 10324
rect 10803 10268 10859 10324
rect 10927 10268 10983 10324
rect 11051 10268 11107 10324
rect 11175 10268 11231 10324
rect 11299 10268 11355 10324
rect 11423 10268 11479 10324
rect 11547 10268 11603 10324
rect 11671 10268 11727 10324
rect 11795 10268 11851 10324
rect 11919 10268 11975 10324
rect 12043 10268 12099 10324
rect 12167 10268 12223 10324
rect 12291 10268 12347 10324
rect 12415 10268 12471 10324
rect 10679 10144 10735 10200
rect 10803 10144 10859 10200
rect 10927 10144 10983 10200
rect 11051 10144 11107 10200
rect 11175 10144 11231 10200
rect 11299 10144 11355 10200
rect 11423 10144 11479 10200
rect 11547 10144 11603 10200
rect 11671 10144 11727 10200
rect 11795 10144 11851 10200
rect 11919 10144 11975 10200
rect 12043 10144 12099 10200
rect 12167 10144 12223 10200
rect 12291 10144 12347 10200
rect 12415 10144 12471 10200
rect 10679 10020 10735 10076
rect 10803 10020 10859 10076
rect 10927 10020 10983 10076
rect 11051 10020 11107 10076
rect 11175 10020 11231 10076
rect 11299 10020 11355 10076
rect 11423 10020 11479 10076
rect 11547 10020 11603 10076
rect 11671 10020 11727 10076
rect 11795 10020 11851 10076
rect 11919 10020 11975 10076
rect 12043 10020 12099 10076
rect 12167 10020 12223 10076
rect 12291 10020 12347 10076
rect 12415 10020 12471 10076
rect 10679 9896 10735 9952
rect 10803 9896 10859 9952
rect 10927 9896 10983 9952
rect 11051 9896 11107 9952
rect 11175 9896 11231 9952
rect 11299 9896 11355 9952
rect 11423 9896 11479 9952
rect 11547 9896 11603 9952
rect 11671 9896 11727 9952
rect 11795 9896 11851 9952
rect 11919 9896 11975 9952
rect 12043 9896 12099 9952
rect 12167 9896 12223 9952
rect 12291 9896 12347 9952
rect 12415 9896 12471 9952
rect 10679 9772 10735 9828
rect 10803 9772 10859 9828
rect 10927 9772 10983 9828
rect 11051 9772 11107 9828
rect 11175 9772 11231 9828
rect 11299 9772 11355 9828
rect 11423 9772 11479 9828
rect 11547 9772 11603 9828
rect 11671 9772 11727 9828
rect 11795 9772 11851 9828
rect 11919 9772 11975 9828
rect 12043 9772 12099 9828
rect 12167 9772 12223 9828
rect 12291 9772 12347 9828
rect 12415 9772 12471 9828
rect 10679 9648 10735 9704
rect 10803 9648 10859 9704
rect 10927 9648 10983 9704
rect 11051 9648 11107 9704
rect 11175 9648 11231 9704
rect 11299 9648 11355 9704
rect 11423 9648 11479 9704
rect 11547 9648 11603 9704
rect 11671 9648 11727 9704
rect 11795 9648 11851 9704
rect 11919 9648 11975 9704
rect 12043 9648 12099 9704
rect 12167 9648 12223 9704
rect 12291 9648 12347 9704
rect 12415 9648 12471 9704
rect 2507 9294 2563 9350
rect 2631 9294 2687 9350
rect 2755 9294 2811 9350
rect 2879 9294 2935 9350
rect 3003 9294 3059 9350
rect 3127 9294 3183 9350
rect 3251 9294 3307 9350
rect 3375 9294 3431 9350
rect 3499 9294 3555 9350
rect 3623 9294 3679 9350
rect 3747 9294 3803 9350
rect 3871 9294 3927 9350
rect 3995 9294 4051 9350
rect 4119 9294 4175 9350
rect 4243 9294 4299 9350
rect 2507 9170 2563 9226
rect 2631 9170 2687 9226
rect 2755 9170 2811 9226
rect 2879 9170 2935 9226
rect 3003 9170 3059 9226
rect 3127 9170 3183 9226
rect 3251 9170 3307 9226
rect 3375 9170 3431 9226
rect 3499 9170 3555 9226
rect 3623 9170 3679 9226
rect 3747 9170 3803 9226
rect 3871 9170 3927 9226
rect 3995 9170 4051 9226
rect 4119 9170 4175 9226
rect 4243 9170 4299 9226
rect 2507 9046 2563 9102
rect 2631 9046 2687 9102
rect 2755 9046 2811 9102
rect 2879 9046 2935 9102
rect 3003 9046 3059 9102
rect 3127 9046 3183 9102
rect 3251 9046 3307 9102
rect 3375 9046 3431 9102
rect 3499 9046 3555 9102
rect 3623 9046 3679 9102
rect 3747 9046 3803 9102
rect 3871 9046 3927 9102
rect 3995 9046 4051 9102
rect 4119 9046 4175 9102
rect 4243 9046 4299 9102
rect 2507 8922 2563 8978
rect 2631 8922 2687 8978
rect 2755 8922 2811 8978
rect 2879 8922 2935 8978
rect 3003 8922 3059 8978
rect 3127 8922 3183 8978
rect 3251 8922 3307 8978
rect 3375 8922 3431 8978
rect 3499 8922 3555 8978
rect 3623 8922 3679 8978
rect 3747 8922 3803 8978
rect 3871 8922 3927 8978
rect 3995 8922 4051 8978
rect 4119 8922 4175 8978
rect 4243 8922 4299 8978
rect 2507 8798 2563 8854
rect 2631 8798 2687 8854
rect 2755 8798 2811 8854
rect 2879 8798 2935 8854
rect 3003 8798 3059 8854
rect 3127 8798 3183 8854
rect 3251 8798 3307 8854
rect 3375 8798 3431 8854
rect 3499 8798 3555 8854
rect 3623 8798 3679 8854
rect 3747 8798 3803 8854
rect 3871 8798 3927 8854
rect 3995 8798 4051 8854
rect 4119 8798 4175 8854
rect 4243 8798 4299 8854
rect 2507 8674 2563 8730
rect 2631 8674 2687 8730
rect 2755 8674 2811 8730
rect 2879 8674 2935 8730
rect 3003 8674 3059 8730
rect 3127 8674 3183 8730
rect 3251 8674 3307 8730
rect 3375 8674 3431 8730
rect 3499 8674 3555 8730
rect 3623 8674 3679 8730
rect 3747 8674 3803 8730
rect 3871 8674 3927 8730
rect 3995 8674 4051 8730
rect 4119 8674 4175 8730
rect 4243 8674 4299 8730
rect 2507 8550 2563 8606
rect 2631 8550 2687 8606
rect 2755 8550 2811 8606
rect 2879 8550 2935 8606
rect 3003 8550 3059 8606
rect 3127 8550 3183 8606
rect 3251 8550 3307 8606
rect 3375 8550 3431 8606
rect 3499 8550 3555 8606
rect 3623 8550 3679 8606
rect 3747 8550 3803 8606
rect 3871 8550 3927 8606
rect 3995 8550 4051 8606
rect 4119 8550 4175 8606
rect 4243 8550 4299 8606
rect 2507 8426 2563 8482
rect 2631 8426 2687 8482
rect 2755 8426 2811 8482
rect 2879 8426 2935 8482
rect 3003 8426 3059 8482
rect 3127 8426 3183 8482
rect 3251 8426 3307 8482
rect 3375 8426 3431 8482
rect 3499 8426 3555 8482
rect 3623 8426 3679 8482
rect 3747 8426 3803 8482
rect 3871 8426 3927 8482
rect 3995 8426 4051 8482
rect 4119 8426 4175 8482
rect 4243 8426 4299 8482
rect 2507 8302 2563 8358
rect 2631 8302 2687 8358
rect 2755 8302 2811 8358
rect 2879 8302 2935 8358
rect 3003 8302 3059 8358
rect 3127 8302 3183 8358
rect 3251 8302 3307 8358
rect 3375 8302 3431 8358
rect 3499 8302 3555 8358
rect 3623 8302 3679 8358
rect 3747 8302 3803 8358
rect 3871 8302 3927 8358
rect 3995 8302 4051 8358
rect 4119 8302 4175 8358
rect 4243 8302 4299 8358
rect 2507 8178 2563 8234
rect 2631 8178 2687 8234
rect 2755 8178 2811 8234
rect 2879 8178 2935 8234
rect 3003 8178 3059 8234
rect 3127 8178 3183 8234
rect 3251 8178 3307 8234
rect 3375 8178 3431 8234
rect 3499 8178 3555 8234
rect 3623 8178 3679 8234
rect 3747 8178 3803 8234
rect 3871 8178 3927 8234
rect 3995 8178 4051 8234
rect 4119 8178 4175 8234
rect 4243 8178 4299 8234
rect 2507 8054 2563 8110
rect 2631 8054 2687 8110
rect 2755 8054 2811 8110
rect 2879 8054 2935 8110
rect 3003 8054 3059 8110
rect 3127 8054 3183 8110
rect 3251 8054 3307 8110
rect 3375 8054 3431 8110
rect 3499 8054 3555 8110
rect 3623 8054 3679 8110
rect 3747 8054 3803 8110
rect 3871 8054 3927 8110
rect 3995 8054 4051 8110
rect 4119 8054 4175 8110
rect 4243 8054 4299 8110
rect 2507 7930 2563 7986
rect 2631 7930 2687 7986
rect 2755 7930 2811 7986
rect 2879 7930 2935 7986
rect 3003 7930 3059 7986
rect 3127 7930 3183 7986
rect 3251 7930 3307 7986
rect 3375 7930 3431 7986
rect 3499 7930 3555 7986
rect 3623 7930 3679 7986
rect 3747 7930 3803 7986
rect 3871 7930 3927 7986
rect 3995 7930 4051 7986
rect 4119 7930 4175 7986
rect 4243 7930 4299 7986
rect 2507 7806 2563 7862
rect 2631 7806 2687 7862
rect 2755 7806 2811 7862
rect 2879 7806 2935 7862
rect 3003 7806 3059 7862
rect 3127 7806 3183 7862
rect 3251 7806 3307 7862
rect 3375 7806 3431 7862
rect 3499 7806 3555 7862
rect 3623 7806 3679 7862
rect 3747 7806 3803 7862
rect 3871 7806 3927 7862
rect 3995 7806 4051 7862
rect 4119 7806 4175 7862
rect 4243 7806 4299 7862
rect 2507 7682 2563 7738
rect 2631 7682 2687 7738
rect 2755 7682 2811 7738
rect 2879 7682 2935 7738
rect 3003 7682 3059 7738
rect 3127 7682 3183 7738
rect 3251 7682 3307 7738
rect 3375 7682 3431 7738
rect 3499 7682 3555 7738
rect 3623 7682 3679 7738
rect 3747 7682 3803 7738
rect 3871 7682 3927 7738
rect 3995 7682 4051 7738
rect 4119 7682 4175 7738
rect 4243 7682 4299 7738
rect 2507 7558 2563 7614
rect 2631 7558 2687 7614
rect 2755 7558 2811 7614
rect 2879 7558 2935 7614
rect 3003 7558 3059 7614
rect 3127 7558 3183 7614
rect 3251 7558 3307 7614
rect 3375 7558 3431 7614
rect 3499 7558 3555 7614
rect 3623 7558 3679 7614
rect 3747 7558 3803 7614
rect 3871 7558 3927 7614
rect 3995 7558 4051 7614
rect 4119 7558 4175 7614
rect 4243 7558 4299 7614
rect 2507 7434 2563 7490
rect 2631 7434 2687 7490
rect 2755 7434 2811 7490
rect 2879 7434 2935 7490
rect 3003 7434 3059 7490
rect 3127 7434 3183 7490
rect 3251 7434 3307 7490
rect 3375 7434 3431 7490
rect 3499 7434 3555 7490
rect 3623 7434 3679 7490
rect 3747 7434 3803 7490
rect 3871 7434 3927 7490
rect 3995 7434 4051 7490
rect 4119 7434 4175 7490
rect 4243 7434 4299 7490
rect 2507 7310 2563 7366
rect 2631 7310 2687 7366
rect 2755 7310 2811 7366
rect 2879 7310 2935 7366
rect 3003 7310 3059 7366
rect 3127 7310 3183 7366
rect 3251 7310 3307 7366
rect 3375 7310 3431 7366
rect 3499 7310 3555 7366
rect 3623 7310 3679 7366
rect 3747 7310 3803 7366
rect 3871 7310 3927 7366
rect 3995 7310 4051 7366
rect 4119 7310 4175 7366
rect 4243 7310 4299 7366
rect 2507 7186 2563 7242
rect 2631 7186 2687 7242
rect 2755 7186 2811 7242
rect 2879 7186 2935 7242
rect 3003 7186 3059 7242
rect 3127 7186 3183 7242
rect 3251 7186 3307 7242
rect 3375 7186 3431 7242
rect 3499 7186 3555 7242
rect 3623 7186 3679 7242
rect 3747 7186 3803 7242
rect 3871 7186 3927 7242
rect 3995 7186 4051 7242
rect 4119 7186 4175 7242
rect 4243 7186 4299 7242
rect 2507 7062 2563 7118
rect 2631 7062 2687 7118
rect 2755 7062 2811 7118
rect 2879 7062 2935 7118
rect 3003 7062 3059 7118
rect 3127 7062 3183 7118
rect 3251 7062 3307 7118
rect 3375 7062 3431 7118
rect 3499 7062 3555 7118
rect 3623 7062 3679 7118
rect 3747 7062 3803 7118
rect 3871 7062 3927 7118
rect 3995 7062 4051 7118
rect 4119 7062 4175 7118
rect 4243 7062 4299 7118
rect 2507 6938 2563 6994
rect 2631 6938 2687 6994
rect 2755 6938 2811 6994
rect 2879 6938 2935 6994
rect 3003 6938 3059 6994
rect 3127 6938 3183 6994
rect 3251 6938 3307 6994
rect 3375 6938 3431 6994
rect 3499 6938 3555 6994
rect 3623 6938 3679 6994
rect 3747 6938 3803 6994
rect 3871 6938 3927 6994
rect 3995 6938 4051 6994
rect 4119 6938 4175 6994
rect 4243 6938 4299 6994
rect 2507 6814 2563 6870
rect 2631 6814 2687 6870
rect 2755 6814 2811 6870
rect 2879 6814 2935 6870
rect 3003 6814 3059 6870
rect 3127 6814 3183 6870
rect 3251 6814 3307 6870
rect 3375 6814 3431 6870
rect 3499 6814 3555 6870
rect 3623 6814 3679 6870
rect 3747 6814 3803 6870
rect 3871 6814 3927 6870
rect 3995 6814 4051 6870
rect 4119 6814 4175 6870
rect 4243 6814 4299 6870
rect 2507 6690 2563 6746
rect 2631 6690 2687 6746
rect 2755 6690 2811 6746
rect 2879 6690 2935 6746
rect 3003 6690 3059 6746
rect 3127 6690 3183 6746
rect 3251 6690 3307 6746
rect 3375 6690 3431 6746
rect 3499 6690 3555 6746
rect 3623 6690 3679 6746
rect 3747 6690 3803 6746
rect 3871 6690 3927 6746
rect 3995 6690 4051 6746
rect 4119 6690 4175 6746
rect 4243 6690 4299 6746
rect 2507 6566 2563 6622
rect 2631 6566 2687 6622
rect 2755 6566 2811 6622
rect 2879 6566 2935 6622
rect 3003 6566 3059 6622
rect 3127 6566 3183 6622
rect 3251 6566 3307 6622
rect 3375 6566 3431 6622
rect 3499 6566 3555 6622
rect 3623 6566 3679 6622
rect 3747 6566 3803 6622
rect 3871 6566 3927 6622
rect 3995 6566 4051 6622
rect 4119 6566 4175 6622
rect 4243 6566 4299 6622
rect 2507 6442 2563 6498
rect 2631 6442 2687 6498
rect 2755 6442 2811 6498
rect 2879 6442 2935 6498
rect 3003 6442 3059 6498
rect 3127 6442 3183 6498
rect 3251 6442 3307 6498
rect 3375 6442 3431 6498
rect 3499 6442 3555 6498
rect 3623 6442 3679 6498
rect 3747 6442 3803 6498
rect 3871 6442 3927 6498
rect 3995 6442 4051 6498
rect 4119 6442 4175 6498
rect 4243 6442 4299 6498
rect 6368 9294 6424 9350
rect 6492 9294 6548 9350
rect 6616 9294 6672 9350
rect 6740 9294 6796 9350
rect 6864 9294 6920 9350
rect 6988 9294 7044 9350
rect 7112 9294 7168 9350
rect 7236 9294 7292 9350
rect 7360 9294 7416 9350
rect 6368 9170 6424 9226
rect 6492 9170 6548 9226
rect 6616 9170 6672 9226
rect 6740 9170 6796 9226
rect 6864 9170 6920 9226
rect 6988 9170 7044 9226
rect 7112 9170 7168 9226
rect 7236 9170 7292 9226
rect 7360 9170 7416 9226
rect 6368 9046 6424 9102
rect 6492 9046 6548 9102
rect 6616 9046 6672 9102
rect 6740 9046 6796 9102
rect 6864 9046 6920 9102
rect 6988 9046 7044 9102
rect 7112 9046 7168 9102
rect 7236 9046 7292 9102
rect 7360 9046 7416 9102
rect 6368 8922 6424 8978
rect 6492 8922 6548 8978
rect 6616 8922 6672 8978
rect 6740 8922 6796 8978
rect 6864 8922 6920 8978
rect 6988 8922 7044 8978
rect 7112 8922 7168 8978
rect 7236 8922 7292 8978
rect 7360 8922 7416 8978
rect 6368 8798 6424 8854
rect 6492 8798 6548 8854
rect 6616 8798 6672 8854
rect 6740 8798 6796 8854
rect 6864 8798 6920 8854
rect 6988 8798 7044 8854
rect 7112 8798 7168 8854
rect 7236 8798 7292 8854
rect 7360 8798 7416 8854
rect 6368 8674 6424 8730
rect 6492 8674 6548 8730
rect 6616 8674 6672 8730
rect 6740 8674 6796 8730
rect 6864 8674 6920 8730
rect 6988 8674 7044 8730
rect 7112 8674 7168 8730
rect 7236 8674 7292 8730
rect 7360 8674 7416 8730
rect 6368 8550 6424 8606
rect 6492 8550 6548 8606
rect 6616 8550 6672 8606
rect 6740 8550 6796 8606
rect 6864 8550 6920 8606
rect 6988 8550 7044 8606
rect 7112 8550 7168 8606
rect 7236 8550 7292 8606
rect 7360 8550 7416 8606
rect 6368 8426 6424 8482
rect 6492 8426 6548 8482
rect 6616 8426 6672 8482
rect 6740 8426 6796 8482
rect 6864 8426 6920 8482
rect 6988 8426 7044 8482
rect 7112 8426 7168 8482
rect 7236 8426 7292 8482
rect 7360 8426 7416 8482
rect 6368 8302 6424 8358
rect 6492 8302 6548 8358
rect 6616 8302 6672 8358
rect 6740 8302 6796 8358
rect 6864 8302 6920 8358
rect 6988 8302 7044 8358
rect 7112 8302 7168 8358
rect 7236 8302 7292 8358
rect 7360 8302 7416 8358
rect 6368 8178 6424 8234
rect 6492 8178 6548 8234
rect 6616 8178 6672 8234
rect 6740 8178 6796 8234
rect 6864 8178 6920 8234
rect 6988 8178 7044 8234
rect 7112 8178 7168 8234
rect 7236 8178 7292 8234
rect 7360 8178 7416 8234
rect 6368 8054 6424 8110
rect 6492 8054 6548 8110
rect 6616 8054 6672 8110
rect 6740 8054 6796 8110
rect 6864 8054 6920 8110
rect 6988 8054 7044 8110
rect 7112 8054 7168 8110
rect 7236 8054 7292 8110
rect 7360 8054 7416 8110
rect 6368 7930 6424 7986
rect 6492 7930 6548 7986
rect 6616 7930 6672 7986
rect 6740 7930 6796 7986
rect 6864 7930 6920 7986
rect 6988 7930 7044 7986
rect 7112 7930 7168 7986
rect 7236 7930 7292 7986
rect 7360 7930 7416 7986
rect 6368 7806 6424 7862
rect 6492 7806 6548 7862
rect 6616 7806 6672 7862
rect 6740 7806 6796 7862
rect 6864 7806 6920 7862
rect 6988 7806 7044 7862
rect 7112 7806 7168 7862
rect 7236 7806 7292 7862
rect 7360 7806 7416 7862
rect 6368 7682 6424 7738
rect 6492 7682 6548 7738
rect 6616 7682 6672 7738
rect 6740 7682 6796 7738
rect 6864 7682 6920 7738
rect 6988 7682 7044 7738
rect 7112 7682 7168 7738
rect 7236 7682 7292 7738
rect 7360 7682 7416 7738
rect 6368 7558 6424 7614
rect 6492 7558 6548 7614
rect 6616 7558 6672 7614
rect 6740 7558 6796 7614
rect 6864 7558 6920 7614
rect 6988 7558 7044 7614
rect 7112 7558 7168 7614
rect 7236 7558 7292 7614
rect 7360 7558 7416 7614
rect 6368 7434 6424 7490
rect 6492 7434 6548 7490
rect 6616 7434 6672 7490
rect 6740 7434 6796 7490
rect 6864 7434 6920 7490
rect 6988 7434 7044 7490
rect 7112 7434 7168 7490
rect 7236 7434 7292 7490
rect 7360 7434 7416 7490
rect 6368 7310 6424 7366
rect 6492 7310 6548 7366
rect 6616 7310 6672 7366
rect 6740 7310 6796 7366
rect 6864 7310 6920 7366
rect 6988 7310 7044 7366
rect 7112 7310 7168 7366
rect 7236 7310 7292 7366
rect 7360 7310 7416 7366
rect 6368 7186 6424 7242
rect 6492 7186 6548 7242
rect 6616 7186 6672 7242
rect 6740 7186 6796 7242
rect 6864 7186 6920 7242
rect 6988 7186 7044 7242
rect 7112 7186 7168 7242
rect 7236 7186 7292 7242
rect 7360 7186 7416 7242
rect 6368 7062 6424 7118
rect 6492 7062 6548 7118
rect 6616 7062 6672 7118
rect 6740 7062 6796 7118
rect 6864 7062 6920 7118
rect 6988 7062 7044 7118
rect 7112 7062 7168 7118
rect 7236 7062 7292 7118
rect 7360 7062 7416 7118
rect 6368 6938 6424 6994
rect 6492 6938 6548 6994
rect 6616 6938 6672 6994
rect 6740 6938 6796 6994
rect 6864 6938 6920 6994
rect 6988 6938 7044 6994
rect 7112 6938 7168 6994
rect 7236 6938 7292 6994
rect 7360 6938 7416 6994
rect 6368 6814 6424 6870
rect 6492 6814 6548 6870
rect 6616 6814 6672 6870
rect 6740 6814 6796 6870
rect 6864 6814 6920 6870
rect 6988 6814 7044 6870
rect 7112 6814 7168 6870
rect 7236 6814 7292 6870
rect 7360 6814 7416 6870
rect 6368 6690 6424 6746
rect 6492 6690 6548 6746
rect 6616 6690 6672 6746
rect 6740 6690 6796 6746
rect 6864 6690 6920 6746
rect 6988 6690 7044 6746
rect 7112 6690 7168 6746
rect 7236 6690 7292 6746
rect 7360 6690 7416 6746
rect 6368 6566 6424 6622
rect 6492 6566 6548 6622
rect 6616 6566 6672 6622
rect 6740 6566 6796 6622
rect 6864 6566 6920 6622
rect 6988 6566 7044 6622
rect 7112 6566 7168 6622
rect 7236 6566 7292 6622
rect 7360 6566 7416 6622
rect 6368 6442 6424 6498
rect 6492 6442 6548 6498
rect 6616 6442 6672 6498
rect 6740 6442 6796 6498
rect 6864 6442 6920 6498
rect 6988 6442 7044 6498
rect 7112 6442 7168 6498
rect 7236 6442 7292 6498
rect 7360 6442 7416 6498
rect 8751 9294 8807 9350
rect 8875 9294 8931 9350
rect 8999 9294 9055 9350
rect 9123 9294 9179 9350
rect 9247 9294 9303 9350
rect 9371 9294 9427 9350
rect 9495 9294 9551 9350
rect 9619 9294 9675 9350
rect 9743 9294 9799 9350
rect 9867 9294 9923 9350
rect 9991 9294 10047 9350
rect 10115 9294 10171 9350
rect 10239 9294 10295 9350
rect 10363 9294 10419 9350
rect 10487 9294 10543 9350
rect 8751 9170 8807 9226
rect 8875 9170 8931 9226
rect 8999 9170 9055 9226
rect 9123 9170 9179 9226
rect 9247 9170 9303 9226
rect 9371 9170 9427 9226
rect 9495 9170 9551 9226
rect 9619 9170 9675 9226
rect 9743 9170 9799 9226
rect 9867 9170 9923 9226
rect 9991 9170 10047 9226
rect 10115 9170 10171 9226
rect 10239 9170 10295 9226
rect 10363 9170 10419 9226
rect 10487 9170 10543 9226
rect 8751 9046 8807 9102
rect 8875 9046 8931 9102
rect 8999 9046 9055 9102
rect 9123 9046 9179 9102
rect 9247 9046 9303 9102
rect 9371 9046 9427 9102
rect 9495 9046 9551 9102
rect 9619 9046 9675 9102
rect 9743 9046 9799 9102
rect 9867 9046 9923 9102
rect 9991 9046 10047 9102
rect 10115 9046 10171 9102
rect 10239 9046 10295 9102
rect 10363 9046 10419 9102
rect 10487 9046 10543 9102
rect 8751 8922 8807 8978
rect 8875 8922 8931 8978
rect 8999 8922 9055 8978
rect 9123 8922 9179 8978
rect 9247 8922 9303 8978
rect 9371 8922 9427 8978
rect 9495 8922 9551 8978
rect 9619 8922 9675 8978
rect 9743 8922 9799 8978
rect 9867 8922 9923 8978
rect 9991 8922 10047 8978
rect 10115 8922 10171 8978
rect 10239 8922 10295 8978
rect 10363 8922 10419 8978
rect 10487 8922 10543 8978
rect 8751 8798 8807 8854
rect 8875 8798 8931 8854
rect 8999 8798 9055 8854
rect 9123 8798 9179 8854
rect 9247 8798 9303 8854
rect 9371 8798 9427 8854
rect 9495 8798 9551 8854
rect 9619 8798 9675 8854
rect 9743 8798 9799 8854
rect 9867 8798 9923 8854
rect 9991 8798 10047 8854
rect 10115 8798 10171 8854
rect 10239 8798 10295 8854
rect 10363 8798 10419 8854
rect 10487 8798 10543 8854
rect 8751 8674 8807 8730
rect 8875 8674 8931 8730
rect 8999 8674 9055 8730
rect 9123 8674 9179 8730
rect 9247 8674 9303 8730
rect 9371 8674 9427 8730
rect 9495 8674 9551 8730
rect 9619 8674 9675 8730
rect 9743 8674 9799 8730
rect 9867 8674 9923 8730
rect 9991 8674 10047 8730
rect 10115 8674 10171 8730
rect 10239 8674 10295 8730
rect 10363 8674 10419 8730
rect 10487 8674 10543 8730
rect 8751 8550 8807 8606
rect 8875 8550 8931 8606
rect 8999 8550 9055 8606
rect 9123 8550 9179 8606
rect 9247 8550 9303 8606
rect 9371 8550 9427 8606
rect 9495 8550 9551 8606
rect 9619 8550 9675 8606
rect 9743 8550 9799 8606
rect 9867 8550 9923 8606
rect 9991 8550 10047 8606
rect 10115 8550 10171 8606
rect 10239 8550 10295 8606
rect 10363 8550 10419 8606
rect 10487 8550 10543 8606
rect 8751 8426 8807 8482
rect 8875 8426 8931 8482
rect 8999 8426 9055 8482
rect 9123 8426 9179 8482
rect 9247 8426 9303 8482
rect 9371 8426 9427 8482
rect 9495 8426 9551 8482
rect 9619 8426 9675 8482
rect 9743 8426 9799 8482
rect 9867 8426 9923 8482
rect 9991 8426 10047 8482
rect 10115 8426 10171 8482
rect 10239 8426 10295 8482
rect 10363 8426 10419 8482
rect 10487 8426 10543 8482
rect 8751 8302 8807 8358
rect 8875 8302 8931 8358
rect 8999 8302 9055 8358
rect 9123 8302 9179 8358
rect 9247 8302 9303 8358
rect 9371 8302 9427 8358
rect 9495 8302 9551 8358
rect 9619 8302 9675 8358
rect 9743 8302 9799 8358
rect 9867 8302 9923 8358
rect 9991 8302 10047 8358
rect 10115 8302 10171 8358
rect 10239 8302 10295 8358
rect 10363 8302 10419 8358
rect 10487 8302 10543 8358
rect 8751 8178 8807 8234
rect 8875 8178 8931 8234
rect 8999 8178 9055 8234
rect 9123 8178 9179 8234
rect 9247 8178 9303 8234
rect 9371 8178 9427 8234
rect 9495 8178 9551 8234
rect 9619 8178 9675 8234
rect 9743 8178 9799 8234
rect 9867 8178 9923 8234
rect 9991 8178 10047 8234
rect 10115 8178 10171 8234
rect 10239 8178 10295 8234
rect 10363 8178 10419 8234
rect 10487 8178 10543 8234
rect 8751 8054 8807 8110
rect 8875 8054 8931 8110
rect 8999 8054 9055 8110
rect 9123 8054 9179 8110
rect 9247 8054 9303 8110
rect 9371 8054 9427 8110
rect 9495 8054 9551 8110
rect 9619 8054 9675 8110
rect 9743 8054 9799 8110
rect 9867 8054 9923 8110
rect 9991 8054 10047 8110
rect 10115 8054 10171 8110
rect 10239 8054 10295 8110
rect 10363 8054 10419 8110
rect 10487 8054 10543 8110
rect 8751 7930 8807 7986
rect 8875 7930 8931 7986
rect 8999 7930 9055 7986
rect 9123 7930 9179 7986
rect 9247 7930 9303 7986
rect 9371 7930 9427 7986
rect 9495 7930 9551 7986
rect 9619 7930 9675 7986
rect 9743 7930 9799 7986
rect 9867 7930 9923 7986
rect 9991 7930 10047 7986
rect 10115 7930 10171 7986
rect 10239 7930 10295 7986
rect 10363 7930 10419 7986
rect 10487 7930 10543 7986
rect 8751 7806 8807 7862
rect 8875 7806 8931 7862
rect 8999 7806 9055 7862
rect 9123 7806 9179 7862
rect 9247 7806 9303 7862
rect 9371 7806 9427 7862
rect 9495 7806 9551 7862
rect 9619 7806 9675 7862
rect 9743 7806 9799 7862
rect 9867 7806 9923 7862
rect 9991 7806 10047 7862
rect 10115 7806 10171 7862
rect 10239 7806 10295 7862
rect 10363 7806 10419 7862
rect 10487 7806 10543 7862
rect 8751 7682 8807 7738
rect 8875 7682 8931 7738
rect 8999 7682 9055 7738
rect 9123 7682 9179 7738
rect 9247 7682 9303 7738
rect 9371 7682 9427 7738
rect 9495 7682 9551 7738
rect 9619 7682 9675 7738
rect 9743 7682 9799 7738
rect 9867 7682 9923 7738
rect 9991 7682 10047 7738
rect 10115 7682 10171 7738
rect 10239 7682 10295 7738
rect 10363 7682 10419 7738
rect 10487 7682 10543 7738
rect 8751 7558 8807 7614
rect 8875 7558 8931 7614
rect 8999 7558 9055 7614
rect 9123 7558 9179 7614
rect 9247 7558 9303 7614
rect 9371 7558 9427 7614
rect 9495 7558 9551 7614
rect 9619 7558 9675 7614
rect 9743 7558 9799 7614
rect 9867 7558 9923 7614
rect 9991 7558 10047 7614
rect 10115 7558 10171 7614
rect 10239 7558 10295 7614
rect 10363 7558 10419 7614
rect 10487 7558 10543 7614
rect 8751 7434 8807 7490
rect 8875 7434 8931 7490
rect 8999 7434 9055 7490
rect 9123 7434 9179 7490
rect 9247 7434 9303 7490
rect 9371 7434 9427 7490
rect 9495 7434 9551 7490
rect 9619 7434 9675 7490
rect 9743 7434 9799 7490
rect 9867 7434 9923 7490
rect 9991 7434 10047 7490
rect 10115 7434 10171 7490
rect 10239 7434 10295 7490
rect 10363 7434 10419 7490
rect 10487 7434 10543 7490
rect 8751 7310 8807 7366
rect 8875 7310 8931 7366
rect 8999 7310 9055 7366
rect 9123 7310 9179 7366
rect 9247 7310 9303 7366
rect 9371 7310 9427 7366
rect 9495 7310 9551 7366
rect 9619 7310 9675 7366
rect 9743 7310 9799 7366
rect 9867 7310 9923 7366
rect 9991 7310 10047 7366
rect 10115 7310 10171 7366
rect 10239 7310 10295 7366
rect 10363 7310 10419 7366
rect 10487 7310 10543 7366
rect 8751 7186 8807 7242
rect 8875 7186 8931 7242
rect 8999 7186 9055 7242
rect 9123 7186 9179 7242
rect 9247 7186 9303 7242
rect 9371 7186 9427 7242
rect 9495 7186 9551 7242
rect 9619 7186 9675 7242
rect 9743 7186 9799 7242
rect 9867 7186 9923 7242
rect 9991 7186 10047 7242
rect 10115 7186 10171 7242
rect 10239 7186 10295 7242
rect 10363 7186 10419 7242
rect 10487 7186 10543 7242
rect 8751 7062 8807 7118
rect 8875 7062 8931 7118
rect 8999 7062 9055 7118
rect 9123 7062 9179 7118
rect 9247 7062 9303 7118
rect 9371 7062 9427 7118
rect 9495 7062 9551 7118
rect 9619 7062 9675 7118
rect 9743 7062 9799 7118
rect 9867 7062 9923 7118
rect 9991 7062 10047 7118
rect 10115 7062 10171 7118
rect 10239 7062 10295 7118
rect 10363 7062 10419 7118
rect 10487 7062 10543 7118
rect 8751 6938 8807 6994
rect 8875 6938 8931 6994
rect 8999 6938 9055 6994
rect 9123 6938 9179 6994
rect 9247 6938 9303 6994
rect 9371 6938 9427 6994
rect 9495 6938 9551 6994
rect 9619 6938 9675 6994
rect 9743 6938 9799 6994
rect 9867 6938 9923 6994
rect 9991 6938 10047 6994
rect 10115 6938 10171 6994
rect 10239 6938 10295 6994
rect 10363 6938 10419 6994
rect 10487 6938 10543 6994
rect 8751 6814 8807 6870
rect 8875 6814 8931 6870
rect 8999 6814 9055 6870
rect 9123 6814 9179 6870
rect 9247 6814 9303 6870
rect 9371 6814 9427 6870
rect 9495 6814 9551 6870
rect 9619 6814 9675 6870
rect 9743 6814 9799 6870
rect 9867 6814 9923 6870
rect 9991 6814 10047 6870
rect 10115 6814 10171 6870
rect 10239 6814 10295 6870
rect 10363 6814 10419 6870
rect 10487 6814 10543 6870
rect 8751 6690 8807 6746
rect 8875 6690 8931 6746
rect 8999 6690 9055 6746
rect 9123 6690 9179 6746
rect 9247 6690 9303 6746
rect 9371 6690 9427 6746
rect 9495 6690 9551 6746
rect 9619 6690 9675 6746
rect 9743 6690 9799 6746
rect 9867 6690 9923 6746
rect 9991 6690 10047 6746
rect 10115 6690 10171 6746
rect 10239 6690 10295 6746
rect 10363 6690 10419 6746
rect 10487 6690 10543 6746
rect 8751 6566 8807 6622
rect 8875 6566 8931 6622
rect 8999 6566 9055 6622
rect 9123 6566 9179 6622
rect 9247 6566 9303 6622
rect 9371 6566 9427 6622
rect 9495 6566 9551 6622
rect 9619 6566 9675 6622
rect 9743 6566 9799 6622
rect 9867 6566 9923 6622
rect 9991 6566 10047 6622
rect 10115 6566 10171 6622
rect 10239 6566 10295 6622
rect 10363 6566 10419 6622
rect 10487 6566 10543 6622
rect 8751 6442 8807 6498
rect 8875 6442 8931 6498
rect 8999 6442 9055 6498
rect 9123 6442 9179 6498
rect 9247 6442 9303 6498
rect 9371 6442 9427 6498
rect 9495 6442 9551 6498
rect 9619 6442 9675 6498
rect 9743 6442 9799 6498
rect 9867 6442 9923 6498
rect 9991 6442 10047 6498
rect 10115 6442 10171 6498
rect 10239 6442 10295 6498
rect 10363 6442 10419 6498
rect 10487 6442 10543 6498
rect 12852 9294 12908 9350
rect 12976 9294 13032 9350
rect 13100 9294 13156 9350
rect 13224 9294 13280 9350
rect 13348 9294 13404 9350
rect 13472 9294 13528 9350
rect 13596 9294 13652 9350
rect 13720 9294 13776 9350
rect 13844 9294 13900 9350
rect 12852 9170 12908 9226
rect 12976 9170 13032 9226
rect 13100 9170 13156 9226
rect 13224 9170 13280 9226
rect 13348 9170 13404 9226
rect 13472 9170 13528 9226
rect 13596 9170 13652 9226
rect 13720 9170 13776 9226
rect 13844 9170 13900 9226
rect 12852 9046 12908 9102
rect 12976 9046 13032 9102
rect 13100 9046 13156 9102
rect 13224 9046 13280 9102
rect 13348 9046 13404 9102
rect 13472 9046 13528 9102
rect 13596 9046 13652 9102
rect 13720 9046 13776 9102
rect 13844 9046 13900 9102
rect 12852 8922 12908 8978
rect 12976 8922 13032 8978
rect 13100 8922 13156 8978
rect 13224 8922 13280 8978
rect 13348 8922 13404 8978
rect 13472 8922 13528 8978
rect 13596 8922 13652 8978
rect 13720 8922 13776 8978
rect 13844 8922 13900 8978
rect 12852 8798 12908 8854
rect 12976 8798 13032 8854
rect 13100 8798 13156 8854
rect 13224 8798 13280 8854
rect 13348 8798 13404 8854
rect 13472 8798 13528 8854
rect 13596 8798 13652 8854
rect 13720 8798 13776 8854
rect 13844 8798 13900 8854
rect 12852 8674 12908 8730
rect 12976 8674 13032 8730
rect 13100 8674 13156 8730
rect 13224 8674 13280 8730
rect 13348 8674 13404 8730
rect 13472 8674 13528 8730
rect 13596 8674 13652 8730
rect 13720 8674 13776 8730
rect 13844 8674 13900 8730
rect 12852 8550 12908 8606
rect 12976 8550 13032 8606
rect 13100 8550 13156 8606
rect 13224 8550 13280 8606
rect 13348 8550 13404 8606
rect 13472 8550 13528 8606
rect 13596 8550 13652 8606
rect 13720 8550 13776 8606
rect 13844 8550 13900 8606
rect 12852 8426 12908 8482
rect 12976 8426 13032 8482
rect 13100 8426 13156 8482
rect 13224 8426 13280 8482
rect 13348 8426 13404 8482
rect 13472 8426 13528 8482
rect 13596 8426 13652 8482
rect 13720 8426 13776 8482
rect 13844 8426 13900 8482
rect 12852 8302 12908 8358
rect 12976 8302 13032 8358
rect 13100 8302 13156 8358
rect 13224 8302 13280 8358
rect 13348 8302 13404 8358
rect 13472 8302 13528 8358
rect 13596 8302 13652 8358
rect 13720 8302 13776 8358
rect 13844 8302 13900 8358
rect 12852 8178 12908 8234
rect 12976 8178 13032 8234
rect 13100 8178 13156 8234
rect 13224 8178 13280 8234
rect 13348 8178 13404 8234
rect 13472 8178 13528 8234
rect 13596 8178 13652 8234
rect 13720 8178 13776 8234
rect 13844 8178 13900 8234
rect 12852 8054 12908 8110
rect 12976 8054 13032 8110
rect 13100 8054 13156 8110
rect 13224 8054 13280 8110
rect 13348 8054 13404 8110
rect 13472 8054 13528 8110
rect 13596 8054 13652 8110
rect 13720 8054 13776 8110
rect 13844 8054 13900 8110
rect 12852 7930 12908 7986
rect 12976 7930 13032 7986
rect 13100 7930 13156 7986
rect 13224 7930 13280 7986
rect 13348 7930 13404 7986
rect 13472 7930 13528 7986
rect 13596 7930 13652 7986
rect 13720 7930 13776 7986
rect 13844 7930 13900 7986
rect 12852 7806 12908 7862
rect 12976 7806 13032 7862
rect 13100 7806 13156 7862
rect 13224 7806 13280 7862
rect 13348 7806 13404 7862
rect 13472 7806 13528 7862
rect 13596 7806 13652 7862
rect 13720 7806 13776 7862
rect 13844 7806 13900 7862
rect 12852 7682 12908 7738
rect 12976 7682 13032 7738
rect 13100 7682 13156 7738
rect 13224 7682 13280 7738
rect 13348 7682 13404 7738
rect 13472 7682 13528 7738
rect 13596 7682 13652 7738
rect 13720 7682 13776 7738
rect 13844 7682 13900 7738
rect 12852 7558 12908 7614
rect 12976 7558 13032 7614
rect 13100 7558 13156 7614
rect 13224 7558 13280 7614
rect 13348 7558 13404 7614
rect 13472 7558 13528 7614
rect 13596 7558 13652 7614
rect 13720 7558 13776 7614
rect 13844 7558 13900 7614
rect 12852 7434 12908 7490
rect 12976 7434 13032 7490
rect 13100 7434 13156 7490
rect 13224 7434 13280 7490
rect 13348 7434 13404 7490
rect 13472 7434 13528 7490
rect 13596 7434 13652 7490
rect 13720 7434 13776 7490
rect 13844 7434 13900 7490
rect 12852 7310 12908 7366
rect 12976 7310 13032 7366
rect 13100 7310 13156 7366
rect 13224 7310 13280 7366
rect 13348 7310 13404 7366
rect 13472 7310 13528 7366
rect 13596 7310 13652 7366
rect 13720 7310 13776 7366
rect 13844 7310 13900 7366
rect 12852 7186 12908 7242
rect 12976 7186 13032 7242
rect 13100 7186 13156 7242
rect 13224 7186 13280 7242
rect 13348 7186 13404 7242
rect 13472 7186 13528 7242
rect 13596 7186 13652 7242
rect 13720 7186 13776 7242
rect 13844 7186 13900 7242
rect 12852 7062 12908 7118
rect 12976 7062 13032 7118
rect 13100 7062 13156 7118
rect 13224 7062 13280 7118
rect 13348 7062 13404 7118
rect 13472 7062 13528 7118
rect 13596 7062 13652 7118
rect 13720 7062 13776 7118
rect 13844 7062 13900 7118
rect 12852 6938 12908 6994
rect 12976 6938 13032 6994
rect 13100 6938 13156 6994
rect 13224 6938 13280 6994
rect 13348 6938 13404 6994
rect 13472 6938 13528 6994
rect 13596 6938 13652 6994
rect 13720 6938 13776 6994
rect 13844 6938 13900 6994
rect 12852 6814 12908 6870
rect 12976 6814 13032 6870
rect 13100 6814 13156 6870
rect 13224 6814 13280 6870
rect 13348 6814 13404 6870
rect 13472 6814 13528 6870
rect 13596 6814 13652 6870
rect 13720 6814 13776 6870
rect 13844 6814 13900 6870
rect 12852 6690 12908 6746
rect 12976 6690 13032 6746
rect 13100 6690 13156 6746
rect 13224 6690 13280 6746
rect 13348 6690 13404 6746
rect 13472 6690 13528 6746
rect 13596 6690 13652 6746
rect 13720 6690 13776 6746
rect 13844 6690 13900 6746
rect 12852 6566 12908 6622
rect 12976 6566 13032 6622
rect 13100 6566 13156 6622
rect 13224 6566 13280 6622
rect 13348 6566 13404 6622
rect 13472 6566 13528 6622
rect 13596 6566 13652 6622
rect 13720 6566 13776 6622
rect 13844 6566 13900 6622
rect 12852 6442 12908 6498
rect 12976 6442 13032 6498
rect 13100 6442 13156 6498
rect 13224 6442 13280 6498
rect 13348 6442 13404 6498
rect 13472 6442 13528 6498
rect 13596 6442 13652 6498
rect 13720 6442 13776 6498
rect 13844 6442 13900 6498
rect 2507 6094 2563 6150
rect 2631 6094 2687 6150
rect 2755 6094 2811 6150
rect 2879 6094 2935 6150
rect 3003 6094 3059 6150
rect 3127 6094 3183 6150
rect 3251 6094 3307 6150
rect 3375 6094 3431 6150
rect 3499 6094 3555 6150
rect 3623 6094 3679 6150
rect 3747 6094 3803 6150
rect 3871 6094 3927 6150
rect 3995 6094 4051 6150
rect 4119 6094 4175 6150
rect 4243 6094 4299 6150
rect 2507 5970 2563 6026
rect 2631 5970 2687 6026
rect 2755 5970 2811 6026
rect 2879 5970 2935 6026
rect 3003 5970 3059 6026
rect 3127 5970 3183 6026
rect 3251 5970 3307 6026
rect 3375 5970 3431 6026
rect 3499 5970 3555 6026
rect 3623 5970 3679 6026
rect 3747 5970 3803 6026
rect 3871 5970 3927 6026
rect 3995 5970 4051 6026
rect 4119 5970 4175 6026
rect 4243 5970 4299 6026
rect 2507 5846 2563 5902
rect 2631 5846 2687 5902
rect 2755 5846 2811 5902
rect 2879 5846 2935 5902
rect 3003 5846 3059 5902
rect 3127 5846 3183 5902
rect 3251 5846 3307 5902
rect 3375 5846 3431 5902
rect 3499 5846 3555 5902
rect 3623 5846 3679 5902
rect 3747 5846 3803 5902
rect 3871 5846 3927 5902
rect 3995 5846 4051 5902
rect 4119 5846 4175 5902
rect 4243 5846 4299 5902
rect 2507 5722 2563 5778
rect 2631 5722 2687 5778
rect 2755 5722 2811 5778
rect 2879 5722 2935 5778
rect 3003 5722 3059 5778
rect 3127 5722 3183 5778
rect 3251 5722 3307 5778
rect 3375 5722 3431 5778
rect 3499 5722 3555 5778
rect 3623 5722 3679 5778
rect 3747 5722 3803 5778
rect 3871 5722 3927 5778
rect 3995 5722 4051 5778
rect 4119 5722 4175 5778
rect 4243 5722 4299 5778
rect 2507 5598 2563 5654
rect 2631 5598 2687 5654
rect 2755 5598 2811 5654
rect 2879 5598 2935 5654
rect 3003 5598 3059 5654
rect 3127 5598 3183 5654
rect 3251 5598 3307 5654
rect 3375 5598 3431 5654
rect 3499 5598 3555 5654
rect 3623 5598 3679 5654
rect 3747 5598 3803 5654
rect 3871 5598 3927 5654
rect 3995 5598 4051 5654
rect 4119 5598 4175 5654
rect 4243 5598 4299 5654
rect 2507 5474 2563 5530
rect 2631 5474 2687 5530
rect 2755 5474 2811 5530
rect 2879 5474 2935 5530
rect 3003 5474 3059 5530
rect 3127 5474 3183 5530
rect 3251 5474 3307 5530
rect 3375 5474 3431 5530
rect 3499 5474 3555 5530
rect 3623 5474 3679 5530
rect 3747 5474 3803 5530
rect 3871 5474 3927 5530
rect 3995 5474 4051 5530
rect 4119 5474 4175 5530
rect 4243 5474 4299 5530
rect 2507 5350 2563 5406
rect 2631 5350 2687 5406
rect 2755 5350 2811 5406
rect 2879 5350 2935 5406
rect 3003 5350 3059 5406
rect 3127 5350 3183 5406
rect 3251 5350 3307 5406
rect 3375 5350 3431 5406
rect 3499 5350 3555 5406
rect 3623 5350 3679 5406
rect 3747 5350 3803 5406
rect 3871 5350 3927 5406
rect 3995 5350 4051 5406
rect 4119 5350 4175 5406
rect 4243 5350 4299 5406
rect 2507 5226 2563 5282
rect 2631 5226 2687 5282
rect 2755 5226 2811 5282
rect 2879 5226 2935 5282
rect 3003 5226 3059 5282
rect 3127 5226 3183 5282
rect 3251 5226 3307 5282
rect 3375 5226 3431 5282
rect 3499 5226 3555 5282
rect 3623 5226 3679 5282
rect 3747 5226 3803 5282
rect 3871 5226 3927 5282
rect 3995 5226 4051 5282
rect 4119 5226 4175 5282
rect 4243 5226 4299 5282
rect 2507 5102 2563 5158
rect 2631 5102 2687 5158
rect 2755 5102 2811 5158
rect 2879 5102 2935 5158
rect 3003 5102 3059 5158
rect 3127 5102 3183 5158
rect 3251 5102 3307 5158
rect 3375 5102 3431 5158
rect 3499 5102 3555 5158
rect 3623 5102 3679 5158
rect 3747 5102 3803 5158
rect 3871 5102 3927 5158
rect 3995 5102 4051 5158
rect 4119 5102 4175 5158
rect 4243 5102 4299 5158
rect 2507 4978 2563 5034
rect 2631 4978 2687 5034
rect 2755 4978 2811 5034
rect 2879 4978 2935 5034
rect 3003 4978 3059 5034
rect 3127 4978 3183 5034
rect 3251 4978 3307 5034
rect 3375 4978 3431 5034
rect 3499 4978 3555 5034
rect 3623 4978 3679 5034
rect 3747 4978 3803 5034
rect 3871 4978 3927 5034
rect 3995 4978 4051 5034
rect 4119 4978 4175 5034
rect 4243 4978 4299 5034
rect 2507 4854 2563 4910
rect 2631 4854 2687 4910
rect 2755 4854 2811 4910
rect 2879 4854 2935 4910
rect 3003 4854 3059 4910
rect 3127 4854 3183 4910
rect 3251 4854 3307 4910
rect 3375 4854 3431 4910
rect 3499 4854 3555 4910
rect 3623 4854 3679 4910
rect 3747 4854 3803 4910
rect 3871 4854 3927 4910
rect 3995 4854 4051 4910
rect 4119 4854 4175 4910
rect 4243 4854 4299 4910
rect 2507 4730 2563 4786
rect 2631 4730 2687 4786
rect 2755 4730 2811 4786
rect 2879 4730 2935 4786
rect 3003 4730 3059 4786
rect 3127 4730 3183 4786
rect 3251 4730 3307 4786
rect 3375 4730 3431 4786
rect 3499 4730 3555 4786
rect 3623 4730 3679 4786
rect 3747 4730 3803 4786
rect 3871 4730 3927 4786
rect 3995 4730 4051 4786
rect 4119 4730 4175 4786
rect 4243 4730 4299 4786
rect 2507 4606 2563 4662
rect 2631 4606 2687 4662
rect 2755 4606 2811 4662
rect 2879 4606 2935 4662
rect 3003 4606 3059 4662
rect 3127 4606 3183 4662
rect 3251 4606 3307 4662
rect 3375 4606 3431 4662
rect 3499 4606 3555 4662
rect 3623 4606 3679 4662
rect 3747 4606 3803 4662
rect 3871 4606 3927 4662
rect 3995 4606 4051 4662
rect 4119 4606 4175 4662
rect 4243 4606 4299 4662
rect 2507 4482 2563 4538
rect 2631 4482 2687 4538
rect 2755 4482 2811 4538
rect 2879 4482 2935 4538
rect 3003 4482 3059 4538
rect 3127 4482 3183 4538
rect 3251 4482 3307 4538
rect 3375 4482 3431 4538
rect 3499 4482 3555 4538
rect 3623 4482 3679 4538
rect 3747 4482 3803 4538
rect 3871 4482 3927 4538
rect 3995 4482 4051 4538
rect 4119 4482 4175 4538
rect 4243 4482 4299 4538
rect 2507 4358 2563 4414
rect 2631 4358 2687 4414
rect 2755 4358 2811 4414
rect 2879 4358 2935 4414
rect 3003 4358 3059 4414
rect 3127 4358 3183 4414
rect 3251 4358 3307 4414
rect 3375 4358 3431 4414
rect 3499 4358 3555 4414
rect 3623 4358 3679 4414
rect 3747 4358 3803 4414
rect 3871 4358 3927 4414
rect 3995 4358 4051 4414
rect 4119 4358 4175 4414
rect 4243 4358 4299 4414
rect 2507 4234 2563 4290
rect 2631 4234 2687 4290
rect 2755 4234 2811 4290
rect 2879 4234 2935 4290
rect 3003 4234 3059 4290
rect 3127 4234 3183 4290
rect 3251 4234 3307 4290
rect 3375 4234 3431 4290
rect 3499 4234 3555 4290
rect 3623 4234 3679 4290
rect 3747 4234 3803 4290
rect 3871 4234 3927 4290
rect 3995 4234 4051 4290
rect 4119 4234 4175 4290
rect 4243 4234 4299 4290
rect 2507 4110 2563 4166
rect 2631 4110 2687 4166
rect 2755 4110 2811 4166
rect 2879 4110 2935 4166
rect 3003 4110 3059 4166
rect 3127 4110 3183 4166
rect 3251 4110 3307 4166
rect 3375 4110 3431 4166
rect 3499 4110 3555 4166
rect 3623 4110 3679 4166
rect 3747 4110 3803 4166
rect 3871 4110 3927 4166
rect 3995 4110 4051 4166
rect 4119 4110 4175 4166
rect 4243 4110 4299 4166
rect 2507 3986 2563 4042
rect 2631 3986 2687 4042
rect 2755 3986 2811 4042
rect 2879 3986 2935 4042
rect 3003 3986 3059 4042
rect 3127 3986 3183 4042
rect 3251 3986 3307 4042
rect 3375 3986 3431 4042
rect 3499 3986 3555 4042
rect 3623 3986 3679 4042
rect 3747 3986 3803 4042
rect 3871 3986 3927 4042
rect 3995 3986 4051 4042
rect 4119 3986 4175 4042
rect 4243 3986 4299 4042
rect 2507 3862 2563 3918
rect 2631 3862 2687 3918
rect 2755 3862 2811 3918
rect 2879 3862 2935 3918
rect 3003 3862 3059 3918
rect 3127 3862 3183 3918
rect 3251 3862 3307 3918
rect 3375 3862 3431 3918
rect 3499 3862 3555 3918
rect 3623 3862 3679 3918
rect 3747 3862 3803 3918
rect 3871 3862 3927 3918
rect 3995 3862 4051 3918
rect 4119 3862 4175 3918
rect 4243 3862 4299 3918
rect 2507 3738 2563 3794
rect 2631 3738 2687 3794
rect 2755 3738 2811 3794
rect 2879 3738 2935 3794
rect 3003 3738 3059 3794
rect 3127 3738 3183 3794
rect 3251 3738 3307 3794
rect 3375 3738 3431 3794
rect 3499 3738 3555 3794
rect 3623 3738 3679 3794
rect 3747 3738 3803 3794
rect 3871 3738 3927 3794
rect 3995 3738 4051 3794
rect 4119 3738 4175 3794
rect 4243 3738 4299 3794
rect 2507 3614 2563 3670
rect 2631 3614 2687 3670
rect 2755 3614 2811 3670
rect 2879 3614 2935 3670
rect 3003 3614 3059 3670
rect 3127 3614 3183 3670
rect 3251 3614 3307 3670
rect 3375 3614 3431 3670
rect 3499 3614 3555 3670
rect 3623 3614 3679 3670
rect 3747 3614 3803 3670
rect 3871 3614 3927 3670
rect 3995 3614 4051 3670
rect 4119 3614 4175 3670
rect 4243 3614 4299 3670
rect 2507 3490 2563 3546
rect 2631 3490 2687 3546
rect 2755 3490 2811 3546
rect 2879 3490 2935 3546
rect 3003 3490 3059 3546
rect 3127 3490 3183 3546
rect 3251 3490 3307 3546
rect 3375 3490 3431 3546
rect 3499 3490 3555 3546
rect 3623 3490 3679 3546
rect 3747 3490 3803 3546
rect 3871 3490 3927 3546
rect 3995 3490 4051 3546
rect 4119 3490 4175 3546
rect 4243 3490 4299 3546
rect 2507 3366 2563 3422
rect 2631 3366 2687 3422
rect 2755 3366 2811 3422
rect 2879 3366 2935 3422
rect 3003 3366 3059 3422
rect 3127 3366 3183 3422
rect 3251 3366 3307 3422
rect 3375 3366 3431 3422
rect 3499 3366 3555 3422
rect 3623 3366 3679 3422
rect 3747 3366 3803 3422
rect 3871 3366 3927 3422
rect 3995 3366 4051 3422
rect 4119 3366 4175 3422
rect 4243 3366 4299 3422
rect 2507 3242 2563 3298
rect 2631 3242 2687 3298
rect 2755 3242 2811 3298
rect 2879 3242 2935 3298
rect 3003 3242 3059 3298
rect 3127 3242 3183 3298
rect 3251 3242 3307 3298
rect 3375 3242 3431 3298
rect 3499 3242 3555 3298
rect 3623 3242 3679 3298
rect 3747 3242 3803 3298
rect 3871 3242 3927 3298
rect 3995 3242 4051 3298
rect 4119 3242 4175 3298
rect 4243 3242 4299 3298
rect 6368 6094 6424 6150
rect 6492 6094 6548 6150
rect 6616 6094 6672 6150
rect 6740 6094 6796 6150
rect 6864 6094 6920 6150
rect 6988 6094 7044 6150
rect 7112 6094 7168 6150
rect 7236 6094 7292 6150
rect 7360 6094 7416 6150
rect 6368 5970 6424 6026
rect 6492 5970 6548 6026
rect 6616 5970 6672 6026
rect 6740 5970 6796 6026
rect 6864 5970 6920 6026
rect 6988 5970 7044 6026
rect 7112 5970 7168 6026
rect 7236 5970 7292 6026
rect 7360 5970 7416 6026
rect 6368 5846 6424 5902
rect 6492 5846 6548 5902
rect 6616 5846 6672 5902
rect 6740 5846 6796 5902
rect 6864 5846 6920 5902
rect 6988 5846 7044 5902
rect 7112 5846 7168 5902
rect 7236 5846 7292 5902
rect 7360 5846 7416 5902
rect 6368 5722 6424 5778
rect 6492 5722 6548 5778
rect 6616 5722 6672 5778
rect 6740 5722 6796 5778
rect 6864 5722 6920 5778
rect 6988 5722 7044 5778
rect 7112 5722 7168 5778
rect 7236 5722 7292 5778
rect 7360 5722 7416 5778
rect 6368 5598 6424 5654
rect 6492 5598 6548 5654
rect 6616 5598 6672 5654
rect 6740 5598 6796 5654
rect 6864 5598 6920 5654
rect 6988 5598 7044 5654
rect 7112 5598 7168 5654
rect 7236 5598 7292 5654
rect 7360 5598 7416 5654
rect 6368 5474 6424 5530
rect 6492 5474 6548 5530
rect 6616 5474 6672 5530
rect 6740 5474 6796 5530
rect 6864 5474 6920 5530
rect 6988 5474 7044 5530
rect 7112 5474 7168 5530
rect 7236 5474 7292 5530
rect 7360 5474 7416 5530
rect 6368 5350 6424 5406
rect 6492 5350 6548 5406
rect 6616 5350 6672 5406
rect 6740 5350 6796 5406
rect 6864 5350 6920 5406
rect 6988 5350 7044 5406
rect 7112 5350 7168 5406
rect 7236 5350 7292 5406
rect 7360 5350 7416 5406
rect 6368 5226 6424 5282
rect 6492 5226 6548 5282
rect 6616 5226 6672 5282
rect 6740 5226 6796 5282
rect 6864 5226 6920 5282
rect 6988 5226 7044 5282
rect 7112 5226 7168 5282
rect 7236 5226 7292 5282
rect 7360 5226 7416 5282
rect 6368 5102 6424 5158
rect 6492 5102 6548 5158
rect 6616 5102 6672 5158
rect 6740 5102 6796 5158
rect 6864 5102 6920 5158
rect 6988 5102 7044 5158
rect 7112 5102 7168 5158
rect 7236 5102 7292 5158
rect 7360 5102 7416 5158
rect 6368 4978 6424 5034
rect 6492 4978 6548 5034
rect 6616 4978 6672 5034
rect 6740 4978 6796 5034
rect 6864 4978 6920 5034
rect 6988 4978 7044 5034
rect 7112 4978 7168 5034
rect 7236 4978 7292 5034
rect 7360 4978 7416 5034
rect 6368 4854 6424 4910
rect 6492 4854 6548 4910
rect 6616 4854 6672 4910
rect 6740 4854 6796 4910
rect 6864 4854 6920 4910
rect 6988 4854 7044 4910
rect 7112 4854 7168 4910
rect 7236 4854 7292 4910
rect 7360 4854 7416 4910
rect 6368 4730 6424 4786
rect 6492 4730 6548 4786
rect 6616 4730 6672 4786
rect 6740 4730 6796 4786
rect 6864 4730 6920 4786
rect 6988 4730 7044 4786
rect 7112 4730 7168 4786
rect 7236 4730 7292 4786
rect 7360 4730 7416 4786
rect 6368 4606 6424 4662
rect 6492 4606 6548 4662
rect 6616 4606 6672 4662
rect 6740 4606 6796 4662
rect 6864 4606 6920 4662
rect 6988 4606 7044 4662
rect 7112 4606 7168 4662
rect 7236 4606 7292 4662
rect 7360 4606 7416 4662
rect 6368 4482 6424 4538
rect 6492 4482 6548 4538
rect 6616 4482 6672 4538
rect 6740 4482 6796 4538
rect 6864 4482 6920 4538
rect 6988 4482 7044 4538
rect 7112 4482 7168 4538
rect 7236 4482 7292 4538
rect 7360 4482 7416 4538
rect 6368 4358 6424 4414
rect 6492 4358 6548 4414
rect 6616 4358 6672 4414
rect 6740 4358 6796 4414
rect 6864 4358 6920 4414
rect 6988 4358 7044 4414
rect 7112 4358 7168 4414
rect 7236 4358 7292 4414
rect 7360 4358 7416 4414
rect 6368 4234 6424 4290
rect 6492 4234 6548 4290
rect 6616 4234 6672 4290
rect 6740 4234 6796 4290
rect 6864 4234 6920 4290
rect 6988 4234 7044 4290
rect 7112 4234 7168 4290
rect 7236 4234 7292 4290
rect 7360 4234 7416 4290
rect 6368 4110 6424 4166
rect 6492 4110 6548 4166
rect 6616 4110 6672 4166
rect 6740 4110 6796 4166
rect 6864 4110 6920 4166
rect 6988 4110 7044 4166
rect 7112 4110 7168 4166
rect 7236 4110 7292 4166
rect 7360 4110 7416 4166
rect 6368 3986 6424 4042
rect 6492 3986 6548 4042
rect 6616 3986 6672 4042
rect 6740 3986 6796 4042
rect 6864 3986 6920 4042
rect 6988 3986 7044 4042
rect 7112 3986 7168 4042
rect 7236 3986 7292 4042
rect 7360 3986 7416 4042
rect 6368 3862 6424 3918
rect 6492 3862 6548 3918
rect 6616 3862 6672 3918
rect 6740 3862 6796 3918
rect 6864 3862 6920 3918
rect 6988 3862 7044 3918
rect 7112 3862 7168 3918
rect 7236 3862 7292 3918
rect 7360 3862 7416 3918
rect 6368 3738 6424 3794
rect 6492 3738 6548 3794
rect 6616 3738 6672 3794
rect 6740 3738 6796 3794
rect 6864 3738 6920 3794
rect 6988 3738 7044 3794
rect 7112 3738 7168 3794
rect 7236 3738 7292 3794
rect 7360 3738 7416 3794
rect 6368 3614 6424 3670
rect 6492 3614 6548 3670
rect 6616 3614 6672 3670
rect 6740 3614 6796 3670
rect 6864 3614 6920 3670
rect 6988 3614 7044 3670
rect 7112 3614 7168 3670
rect 7236 3614 7292 3670
rect 7360 3614 7416 3670
rect 6368 3490 6424 3546
rect 6492 3490 6548 3546
rect 6616 3490 6672 3546
rect 6740 3490 6796 3546
rect 6864 3490 6920 3546
rect 6988 3490 7044 3546
rect 7112 3490 7168 3546
rect 7236 3490 7292 3546
rect 7360 3490 7416 3546
rect 6368 3366 6424 3422
rect 6492 3366 6548 3422
rect 6616 3366 6672 3422
rect 6740 3366 6796 3422
rect 6864 3366 6920 3422
rect 6988 3366 7044 3422
rect 7112 3366 7168 3422
rect 7236 3366 7292 3422
rect 7360 3366 7416 3422
rect 6368 3242 6424 3298
rect 6492 3242 6548 3298
rect 6616 3242 6672 3298
rect 6740 3242 6796 3298
rect 6864 3242 6920 3298
rect 6988 3242 7044 3298
rect 7112 3242 7168 3298
rect 7236 3242 7292 3298
rect 7360 3242 7416 3298
rect 8751 6094 8807 6150
rect 8875 6094 8931 6150
rect 8999 6094 9055 6150
rect 9123 6094 9179 6150
rect 9247 6094 9303 6150
rect 9371 6094 9427 6150
rect 9495 6094 9551 6150
rect 9619 6094 9675 6150
rect 9743 6094 9799 6150
rect 9867 6094 9923 6150
rect 9991 6094 10047 6150
rect 10115 6094 10171 6150
rect 10239 6094 10295 6150
rect 10363 6094 10419 6150
rect 10487 6094 10543 6150
rect 8751 5970 8807 6026
rect 8875 5970 8931 6026
rect 8999 5970 9055 6026
rect 9123 5970 9179 6026
rect 9247 5970 9303 6026
rect 9371 5970 9427 6026
rect 9495 5970 9551 6026
rect 9619 5970 9675 6026
rect 9743 5970 9799 6026
rect 9867 5970 9923 6026
rect 9991 5970 10047 6026
rect 10115 5970 10171 6026
rect 10239 5970 10295 6026
rect 10363 5970 10419 6026
rect 10487 5970 10543 6026
rect 8751 5846 8807 5902
rect 8875 5846 8931 5902
rect 8999 5846 9055 5902
rect 9123 5846 9179 5902
rect 9247 5846 9303 5902
rect 9371 5846 9427 5902
rect 9495 5846 9551 5902
rect 9619 5846 9675 5902
rect 9743 5846 9799 5902
rect 9867 5846 9923 5902
rect 9991 5846 10047 5902
rect 10115 5846 10171 5902
rect 10239 5846 10295 5902
rect 10363 5846 10419 5902
rect 10487 5846 10543 5902
rect 8751 5722 8807 5778
rect 8875 5722 8931 5778
rect 8999 5722 9055 5778
rect 9123 5722 9179 5778
rect 9247 5722 9303 5778
rect 9371 5722 9427 5778
rect 9495 5722 9551 5778
rect 9619 5722 9675 5778
rect 9743 5722 9799 5778
rect 9867 5722 9923 5778
rect 9991 5722 10047 5778
rect 10115 5722 10171 5778
rect 10239 5722 10295 5778
rect 10363 5722 10419 5778
rect 10487 5722 10543 5778
rect 8751 5598 8807 5654
rect 8875 5598 8931 5654
rect 8999 5598 9055 5654
rect 9123 5598 9179 5654
rect 9247 5598 9303 5654
rect 9371 5598 9427 5654
rect 9495 5598 9551 5654
rect 9619 5598 9675 5654
rect 9743 5598 9799 5654
rect 9867 5598 9923 5654
rect 9991 5598 10047 5654
rect 10115 5598 10171 5654
rect 10239 5598 10295 5654
rect 10363 5598 10419 5654
rect 10487 5598 10543 5654
rect 8751 5474 8807 5530
rect 8875 5474 8931 5530
rect 8999 5474 9055 5530
rect 9123 5474 9179 5530
rect 9247 5474 9303 5530
rect 9371 5474 9427 5530
rect 9495 5474 9551 5530
rect 9619 5474 9675 5530
rect 9743 5474 9799 5530
rect 9867 5474 9923 5530
rect 9991 5474 10047 5530
rect 10115 5474 10171 5530
rect 10239 5474 10295 5530
rect 10363 5474 10419 5530
rect 10487 5474 10543 5530
rect 8751 5350 8807 5406
rect 8875 5350 8931 5406
rect 8999 5350 9055 5406
rect 9123 5350 9179 5406
rect 9247 5350 9303 5406
rect 9371 5350 9427 5406
rect 9495 5350 9551 5406
rect 9619 5350 9675 5406
rect 9743 5350 9799 5406
rect 9867 5350 9923 5406
rect 9991 5350 10047 5406
rect 10115 5350 10171 5406
rect 10239 5350 10295 5406
rect 10363 5350 10419 5406
rect 10487 5350 10543 5406
rect 8751 5226 8807 5282
rect 8875 5226 8931 5282
rect 8999 5226 9055 5282
rect 9123 5226 9179 5282
rect 9247 5226 9303 5282
rect 9371 5226 9427 5282
rect 9495 5226 9551 5282
rect 9619 5226 9675 5282
rect 9743 5226 9799 5282
rect 9867 5226 9923 5282
rect 9991 5226 10047 5282
rect 10115 5226 10171 5282
rect 10239 5226 10295 5282
rect 10363 5226 10419 5282
rect 10487 5226 10543 5282
rect 8751 5102 8807 5158
rect 8875 5102 8931 5158
rect 8999 5102 9055 5158
rect 9123 5102 9179 5158
rect 9247 5102 9303 5158
rect 9371 5102 9427 5158
rect 9495 5102 9551 5158
rect 9619 5102 9675 5158
rect 9743 5102 9799 5158
rect 9867 5102 9923 5158
rect 9991 5102 10047 5158
rect 10115 5102 10171 5158
rect 10239 5102 10295 5158
rect 10363 5102 10419 5158
rect 10487 5102 10543 5158
rect 8751 4978 8807 5034
rect 8875 4978 8931 5034
rect 8999 4978 9055 5034
rect 9123 4978 9179 5034
rect 9247 4978 9303 5034
rect 9371 4978 9427 5034
rect 9495 4978 9551 5034
rect 9619 4978 9675 5034
rect 9743 4978 9799 5034
rect 9867 4978 9923 5034
rect 9991 4978 10047 5034
rect 10115 4978 10171 5034
rect 10239 4978 10295 5034
rect 10363 4978 10419 5034
rect 10487 4978 10543 5034
rect 8751 4854 8807 4910
rect 8875 4854 8931 4910
rect 8999 4854 9055 4910
rect 9123 4854 9179 4910
rect 9247 4854 9303 4910
rect 9371 4854 9427 4910
rect 9495 4854 9551 4910
rect 9619 4854 9675 4910
rect 9743 4854 9799 4910
rect 9867 4854 9923 4910
rect 9991 4854 10047 4910
rect 10115 4854 10171 4910
rect 10239 4854 10295 4910
rect 10363 4854 10419 4910
rect 10487 4854 10543 4910
rect 8751 4730 8807 4786
rect 8875 4730 8931 4786
rect 8999 4730 9055 4786
rect 9123 4730 9179 4786
rect 9247 4730 9303 4786
rect 9371 4730 9427 4786
rect 9495 4730 9551 4786
rect 9619 4730 9675 4786
rect 9743 4730 9799 4786
rect 9867 4730 9923 4786
rect 9991 4730 10047 4786
rect 10115 4730 10171 4786
rect 10239 4730 10295 4786
rect 10363 4730 10419 4786
rect 10487 4730 10543 4786
rect 8751 4606 8807 4662
rect 8875 4606 8931 4662
rect 8999 4606 9055 4662
rect 9123 4606 9179 4662
rect 9247 4606 9303 4662
rect 9371 4606 9427 4662
rect 9495 4606 9551 4662
rect 9619 4606 9675 4662
rect 9743 4606 9799 4662
rect 9867 4606 9923 4662
rect 9991 4606 10047 4662
rect 10115 4606 10171 4662
rect 10239 4606 10295 4662
rect 10363 4606 10419 4662
rect 10487 4606 10543 4662
rect 8751 4482 8807 4538
rect 8875 4482 8931 4538
rect 8999 4482 9055 4538
rect 9123 4482 9179 4538
rect 9247 4482 9303 4538
rect 9371 4482 9427 4538
rect 9495 4482 9551 4538
rect 9619 4482 9675 4538
rect 9743 4482 9799 4538
rect 9867 4482 9923 4538
rect 9991 4482 10047 4538
rect 10115 4482 10171 4538
rect 10239 4482 10295 4538
rect 10363 4482 10419 4538
rect 10487 4482 10543 4538
rect 8751 4358 8807 4414
rect 8875 4358 8931 4414
rect 8999 4358 9055 4414
rect 9123 4358 9179 4414
rect 9247 4358 9303 4414
rect 9371 4358 9427 4414
rect 9495 4358 9551 4414
rect 9619 4358 9675 4414
rect 9743 4358 9799 4414
rect 9867 4358 9923 4414
rect 9991 4358 10047 4414
rect 10115 4358 10171 4414
rect 10239 4358 10295 4414
rect 10363 4358 10419 4414
rect 10487 4358 10543 4414
rect 8751 4234 8807 4290
rect 8875 4234 8931 4290
rect 8999 4234 9055 4290
rect 9123 4234 9179 4290
rect 9247 4234 9303 4290
rect 9371 4234 9427 4290
rect 9495 4234 9551 4290
rect 9619 4234 9675 4290
rect 9743 4234 9799 4290
rect 9867 4234 9923 4290
rect 9991 4234 10047 4290
rect 10115 4234 10171 4290
rect 10239 4234 10295 4290
rect 10363 4234 10419 4290
rect 10487 4234 10543 4290
rect 8751 4110 8807 4166
rect 8875 4110 8931 4166
rect 8999 4110 9055 4166
rect 9123 4110 9179 4166
rect 9247 4110 9303 4166
rect 9371 4110 9427 4166
rect 9495 4110 9551 4166
rect 9619 4110 9675 4166
rect 9743 4110 9799 4166
rect 9867 4110 9923 4166
rect 9991 4110 10047 4166
rect 10115 4110 10171 4166
rect 10239 4110 10295 4166
rect 10363 4110 10419 4166
rect 10487 4110 10543 4166
rect 8751 3986 8807 4042
rect 8875 3986 8931 4042
rect 8999 3986 9055 4042
rect 9123 3986 9179 4042
rect 9247 3986 9303 4042
rect 9371 3986 9427 4042
rect 9495 3986 9551 4042
rect 9619 3986 9675 4042
rect 9743 3986 9799 4042
rect 9867 3986 9923 4042
rect 9991 3986 10047 4042
rect 10115 3986 10171 4042
rect 10239 3986 10295 4042
rect 10363 3986 10419 4042
rect 10487 3986 10543 4042
rect 8751 3862 8807 3918
rect 8875 3862 8931 3918
rect 8999 3862 9055 3918
rect 9123 3862 9179 3918
rect 9247 3862 9303 3918
rect 9371 3862 9427 3918
rect 9495 3862 9551 3918
rect 9619 3862 9675 3918
rect 9743 3862 9799 3918
rect 9867 3862 9923 3918
rect 9991 3862 10047 3918
rect 10115 3862 10171 3918
rect 10239 3862 10295 3918
rect 10363 3862 10419 3918
rect 10487 3862 10543 3918
rect 8751 3738 8807 3794
rect 8875 3738 8931 3794
rect 8999 3738 9055 3794
rect 9123 3738 9179 3794
rect 9247 3738 9303 3794
rect 9371 3738 9427 3794
rect 9495 3738 9551 3794
rect 9619 3738 9675 3794
rect 9743 3738 9799 3794
rect 9867 3738 9923 3794
rect 9991 3738 10047 3794
rect 10115 3738 10171 3794
rect 10239 3738 10295 3794
rect 10363 3738 10419 3794
rect 10487 3738 10543 3794
rect 8751 3614 8807 3670
rect 8875 3614 8931 3670
rect 8999 3614 9055 3670
rect 9123 3614 9179 3670
rect 9247 3614 9303 3670
rect 9371 3614 9427 3670
rect 9495 3614 9551 3670
rect 9619 3614 9675 3670
rect 9743 3614 9799 3670
rect 9867 3614 9923 3670
rect 9991 3614 10047 3670
rect 10115 3614 10171 3670
rect 10239 3614 10295 3670
rect 10363 3614 10419 3670
rect 10487 3614 10543 3670
rect 8751 3490 8807 3546
rect 8875 3490 8931 3546
rect 8999 3490 9055 3546
rect 9123 3490 9179 3546
rect 9247 3490 9303 3546
rect 9371 3490 9427 3546
rect 9495 3490 9551 3546
rect 9619 3490 9675 3546
rect 9743 3490 9799 3546
rect 9867 3490 9923 3546
rect 9991 3490 10047 3546
rect 10115 3490 10171 3546
rect 10239 3490 10295 3546
rect 10363 3490 10419 3546
rect 10487 3490 10543 3546
rect 8751 3366 8807 3422
rect 8875 3366 8931 3422
rect 8999 3366 9055 3422
rect 9123 3366 9179 3422
rect 9247 3366 9303 3422
rect 9371 3366 9427 3422
rect 9495 3366 9551 3422
rect 9619 3366 9675 3422
rect 9743 3366 9799 3422
rect 9867 3366 9923 3422
rect 9991 3366 10047 3422
rect 10115 3366 10171 3422
rect 10239 3366 10295 3422
rect 10363 3366 10419 3422
rect 10487 3366 10543 3422
rect 8751 3242 8807 3298
rect 8875 3242 8931 3298
rect 8999 3242 9055 3298
rect 9123 3242 9179 3298
rect 9247 3242 9303 3298
rect 9371 3242 9427 3298
rect 9495 3242 9551 3298
rect 9619 3242 9675 3298
rect 9743 3242 9799 3298
rect 9867 3242 9923 3298
rect 9991 3242 10047 3298
rect 10115 3242 10171 3298
rect 10239 3242 10295 3298
rect 10363 3242 10419 3298
rect 10487 3242 10543 3298
rect 12852 6094 12908 6150
rect 12976 6094 13032 6150
rect 13100 6094 13156 6150
rect 13224 6094 13280 6150
rect 13348 6094 13404 6150
rect 13472 6094 13528 6150
rect 13596 6094 13652 6150
rect 13720 6094 13776 6150
rect 13844 6094 13900 6150
rect 12852 5970 12908 6026
rect 12976 5970 13032 6026
rect 13100 5970 13156 6026
rect 13224 5970 13280 6026
rect 13348 5970 13404 6026
rect 13472 5970 13528 6026
rect 13596 5970 13652 6026
rect 13720 5970 13776 6026
rect 13844 5970 13900 6026
rect 12852 5846 12908 5902
rect 12976 5846 13032 5902
rect 13100 5846 13156 5902
rect 13224 5846 13280 5902
rect 13348 5846 13404 5902
rect 13472 5846 13528 5902
rect 13596 5846 13652 5902
rect 13720 5846 13776 5902
rect 13844 5846 13900 5902
rect 12852 5722 12908 5778
rect 12976 5722 13032 5778
rect 13100 5722 13156 5778
rect 13224 5722 13280 5778
rect 13348 5722 13404 5778
rect 13472 5722 13528 5778
rect 13596 5722 13652 5778
rect 13720 5722 13776 5778
rect 13844 5722 13900 5778
rect 12852 5598 12908 5654
rect 12976 5598 13032 5654
rect 13100 5598 13156 5654
rect 13224 5598 13280 5654
rect 13348 5598 13404 5654
rect 13472 5598 13528 5654
rect 13596 5598 13652 5654
rect 13720 5598 13776 5654
rect 13844 5598 13900 5654
rect 12852 5474 12908 5530
rect 12976 5474 13032 5530
rect 13100 5474 13156 5530
rect 13224 5474 13280 5530
rect 13348 5474 13404 5530
rect 13472 5474 13528 5530
rect 13596 5474 13652 5530
rect 13720 5474 13776 5530
rect 13844 5474 13900 5530
rect 12852 5350 12908 5406
rect 12976 5350 13032 5406
rect 13100 5350 13156 5406
rect 13224 5350 13280 5406
rect 13348 5350 13404 5406
rect 13472 5350 13528 5406
rect 13596 5350 13652 5406
rect 13720 5350 13776 5406
rect 13844 5350 13900 5406
rect 12852 5226 12908 5282
rect 12976 5226 13032 5282
rect 13100 5226 13156 5282
rect 13224 5226 13280 5282
rect 13348 5226 13404 5282
rect 13472 5226 13528 5282
rect 13596 5226 13652 5282
rect 13720 5226 13776 5282
rect 13844 5226 13900 5282
rect 12852 5102 12908 5158
rect 12976 5102 13032 5158
rect 13100 5102 13156 5158
rect 13224 5102 13280 5158
rect 13348 5102 13404 5158
rect 13472 5102 13528 5158
rect 13596 5102 13652 5158
rect 13720 5102 13776 5158
rect 13844 5102 13900 5158
rect 12852 4978 12908 5034
rect 12976 4978 13032 5034
rect 13100 4978 13156 5034
rect 13224 4978 13280 5034
rect 13348 4978 13404 5034
rect 13472 4978 13528 5034
rect 13596 4978 13652 5034
rect 13720 4978 13776 5034
rect 13844 4978 13900 5034
rect 12852 4854 12908 4910
rect 12976 4854 13032 4910
rect 13100 4854 13156 4910
rect 13224 4854 13280 4910
rect 13348 4854 13404 4910
rect 13472 4854 13528 4910
rect 13596 4854 13652 4910
rect 13720 4854 13776 4910
rect 13844 4854 13900 4910
rect 12852 4730 12908 4786
rect 12976 4730 13032 4786
rect 13100 4730 13156 4786
rect 13224 4730 13280 4786
rect 13348 4730 13404 4786
rect 13472 4730 13528 4786
rect 13596 4730 13652 4786
rect 13720 4730 13776 4786
rect 13844 4730 13900 4786
rect 12852 4606 12908 4662
rect 12976 4606 13032 4662
rect 13100 4606 13156 4662
rect 13224 4606 13280 4662
rect 13348 4606 13404 4662
rect 13472 4606 13528 4662
rect 13596 4606 13652 4662
rect 13720 4606 13776 4662
rect 13844 4606 13900 4662
rect 12852 4482 12908 4538
rect 12976 4482 13032 4538
rect 13100 4482 13156 4538
rect 13224 4482 13280 4538
rect 13348 4482 13404 4538
rect 13472 4482 13528 4538
rect 13596 4482 13652 4538
rect 13720 4482 13776 4538
rect 13844 4482 13900 4538
rect 12852 4358 12908 4414
rect 12976 4358 13032 4414
rect 13100 4358 13156 4414
rect 13224 4358 13280 4414
rect 13348 4358 13404 4414
rect 13472 4358 13528 4414
rect 13596 4358 13652 4414
rect 13720 4358 13776 4414
rect 13844 4358 13900 4414
rect 12852 4234 12908 4290
rect 12976 4234 13032 4290
rect 13100 4234 13156 4290
rect 13224 4234 13280 4290
rect 13348 4234 13404 4290
rect 13472 4234 13528 4290
rect 13596 4234 13652 4290
rect 13720 4234 13776 4290
rect 13844 4234 13900 4290
rect 12852 4110 12908 4166
rect 12976 4110 13032 4166
rect 13100 4110 13156 4166
rect 13224 4110 13280 4166
rect 13348 4110 13404 4166
rect 13472 4110 13528 4166
rect 13596 4110 13652 4166
rect 13720 4110 13776 4166
rect 13844 4110 13900 4166
rect 12852 3986 12908 4042
rect 12976 3986 13032 4042
rect 13100 3986 13156 4042
rect 13224 3986 13280 4042
rect 13348 3986 13404 4042
rect 13472 3986 13528 4042
rect 13596 3986 13652 4042
rect 13720 3986 13776 4042
rect 13844 3986 13900 4042
rect 12852 3862 12908 3918
rect 12976 3862 13032 3918
rect 13100 3862 13156 3918
rect 13224 3862 13280 3918
rect 13348 3862 13404 3918
rect 13472 3862 13528 3918
rect 13596 3862 13652 3918
rect 13720 3862 13776 3918
rect 13844 3862 13900 3918
rect 12852 3738 12908 3794
rect 12976 3738 13032 3794
rect 13100 3738 13156 3794
rect 13224 3738 13280 3794
rect 13348 3738 13404 3794
rect 13472 3738 13528 3794
rect 13596 3738 13652 3794
rect 13720 3738 13776 3794
rect 13844 3738 13900 3794
rect 12852 3614 12908 3670
rect 12976 3614 13032 3670
rect 13100 3614 13156 3670
rect 13224 3614 13280 3670
rect 13348 3614 13404 3670
rect 13472 3614 13528 3670
rect 13596 3614 13652 3670
rect 13720 3614 13776 3670
rect 13844 3614 13900 3670
rect 12852 3490 12908 3546
rect 12976 3490 13032 3546
rect 13100 3490 13156 3546
rect 13224 3490 13280 3546
rect 13348 3490 13404 3546
rect 13472 3490 13528 3546
rect 13596 3490 13652 3546
rect 13720 3490 13776 3546
rect 13844 3490 13900 3546
rect 12852 3366 12908 3422
rect 12976 3366 13032 3422
rect 13100 3366 13156 3422
rect 13224 3366 13280 3422
rect 13348 3366 13404 3422
rect 13472 3366 13528 3422
rect 13596 3366 13652 3422
rect 13720 3366 13776 3422
rect 13844 3366 13900 3422
rect 12852 3242 12908 3298
rect 12976 3242 13032 3298
rect 13100 3242 13156 3298
rect 13224 3242 13280 3298
rect 13348 3242 13404 3298
rect 13472 3242 13528 3298
rect 13596 3242 13652 3298
rect 13720 3242 13776 3298
rect 13844 3242 13900 3298
rect 2507 2894 2563 2950
rect 2631 2894 2687 2950
rect 2755 2894 2811 2950
rect 2879 2894 2935 2950
rect 3003 2894 3059 2950
rect 3127 2894 3183 2950
rect 3251 2894 3307 2950
rect 3375 2894 3431 2950
rect 3499 2894 3555 2950
rect 3623 2894 3679 2950
rect 3747 2894 3803 2950
rect 3871 2894 3927 2950
rect 3995 2894 4051 2950
rect 4119 2894 4175 2950
rect 4243 2894 4299 2950
rect 2507 2770 2563 2826
rect 2631 2770 2687 2826
rect 2755 2770 2811 2826
rect 2879 2770 2935 2826
rect 3003 2770 3059 2826
rect 3127 2770 3183 2826
rect 3251 2770 3307 2826
rect 3375 2770 3431 2826
rect 3499 2770 3555 2826
rect 3623 2770 3679 2826
rect 3747 2770 3803 2826
rect 3871 2770 3927 2826
rect 3995 2770 4051 2826
rect 4119 2770 4175 2826
rect 4243 2770 4299 2826
rect 2507 2646 2563 2702
rect 2631 2646 2687 2702
rect 2755 2646 2811 2702
rect 2879 2646 2935 2702
rect 3003 2646 3059 2702
rect 3127 2646 3183 2702
rect 3251 2646 3307 2702
rect 3375 2646 3431 2702
rect 3499 2646 3555 2702
rect 3623 2646 3679 2702
rect 3747 2646 3803 2702
rect 3871 2646 3927 2702
rect 3995 2646 4051 2702
rect 4119 2646 4175 2702
rect 4243 2646 4299 2702
rect 2507 2522 2563 2578
rect 2631 2522 2687 2578
rect 2755 2522 2811 2578
rect 2879 2522 2935 2578
rect 3003 2522 3059 2578
rect 3127 2522 3183 2578
rect 3251 2522 3307 2578
rect 3375 2522 3431 2578
rect 3499 2522 3555 2578
rect 3623 2522 3679 2578
rect 3747 2522 3803 2578
rect 3871 2522 3927 2578
rect 3995 2522 4051 2578
rect 4119 2522 4175 2578
rect 4243 2522 4299 2578
rect 2507 2398 2563 2454
rect 2631 2398 2687 2454
rect 2755 2398 2811 2454
rect 2879 2398 2935 2454
rect 3003 2398 3059 2454
rect 3127 2398 3183 2454
rect 3251 2398 3307 2454
rect 3375 2398 3431 2454
rect 3499 2398 3555 2454
rect 3623 2398 3679 2454
rect 3747 2398 3803 2454
rect 3871 2398 3927 2454
rect 3995 2398 4051 2454
rect 4119 2398 4175 2454
rect 4243 2398 4299 2454
rect 2507 2274 2563 2330
rect 2631 2274 2687 2330
rect 2755 2274 2811 2330
rect 2879 2274 2935 2330
rect 3003 2274 3059 2330
rect 3127 2274 3183 2330
rect 3251 2274 3307 2330
rect 3375 2274 3431 2330
rect 3499 2274 3555 2330
rect 3623 2274 3679 2330
rect 3747 2274 3803 2330
rect 3871 2274 3927 2330
rect 3995 2274 4051 2330
rect 4119 2274 4175 2330
rect 4243 2274 4299 2330
rect 2507 2150 2563 2206
rect 2631 2150 2687 2206
rect 2755 2150 2811 2206
rect 2879 2150 2935 2206
rect 3003 2150 3059 2206
rect 3127 2150 3183 2206
rect 3251 2150 3307 2206
rect 3375 2150 3431 2206
rect 3499 2150 3555 2206
rect 3623 2150 3679 2206
rect 3747 2150 3803 2206
rect 3871 2150 3927 2206
rect 3995 2150 4051 2206
rect 4119 2150 4175 2206
rect 4243 2150 4299 2206
rect 2507 2026 2563 2082
rect 2631 2026 2687 2082
rect 2755 2026 2811 2082
rect 2879 2026 2935 2082
rect 3003 2026 3059 2082
rect 3127 2026 3183 2082
rect 3251 2026 3307 2082
rect 3375 2026 3431 2082
rect 3499 2026 3555 2082
rect 3623 2026 3679 2082
rect 3747 2026 3803 2082
rect 3871 2026 3927 2082
rect 3995 2026 4051 2082
rect 4119 2026 4175 2082
rect 4243 2026 4299 2082
rect 2507 1902 2563 1958
rect 2631 1902 2687 1958
rect 2755 1902 2811 1958
rect 2879 1902 2935 1958
rect 3003 1902 3059 1958
rect 3127 1902 3183 1958
rect 3251 1902 3307 1958
rect 3375 1902 3431 1958
rect 3499 1902 3555 1958
rect 3623 1902 3679 1958
rect 3747 1902 3803 1958
rect 3871 1902 3927 1958
rect 3995 1902 4051 1958
rect 4119 1902 4175 1958
rect 4243 1902 4299 1958
rect 2507 1778 2563 1834
rect 2631 1778 2687 1834
rect 2755 1778 2811 1834
rect 2879 1778 2935 1834
rect 3003 1778 3059 1834
rect 3127 1778 3183 1834
rect 3251 1778 3307 1834
rect 3375 1778 3431 1834
rect 3499 1778 3555 1834
rect 3623 1778 3679 1834
rect 3747 1778 3803 1834
rect 3871 1778 3927 1834
rect 3995 1778 4051 1834
rect 4119 1778 4175 1834
rect 4243 1778 4299 1834
rect 2507 1654 2563 1710
rect 2631 1654 2687 1710
rect 2755 1654 2811 1710
rect 2879 1654 2935 1710
rect 3003 1654 3059 1710
rect 3127 1654 3183 1710
rect 3251 1654 3307 1710
rect 3375 1654 3431 1710
rect 3499 1654 3555 1710
rect 3623 1654 3679 1710
rect 3747 1654 3803 1710
rect 3871 1654 3927 1710
rect 3995 1654 4051 1710
rect 4119 1654 4175 1710
rect 4243 1654 4299 1710
rect 2507 1530 2563 1586
rect 2631 1530 2687 1586
rect 2755 1530 2811 1586
rect 2879 1530 2935 1586
rect 3003 1530 3059 1586
rect 3127 1530 3183 1586
rect 3251 1530 3307 1586
rect 3375 1530 3431 1586
rect 3499 1530 3555 1586
rect 3623 1530 3679 1586
rect 3747 1530 3803 1586
rect 3871 1530 3927 1586
rect 3995 1530 4051 1586
rect 4119 1530 4175 1586
rect 4243 1530 4299 1586
rect 2507 1406 2563 1462
rect 2631 1406 2687 1462
rect 2755 1406 2811 1462
rect 2879 1406 2935 1462
rect 3003 1406 3059 1462
rect 3127 1406 3183 1462
rect 3251 1406 3307 1462
rect 3375 1406 3431 1462
rect 3499 1406 3555 1462
rect 3623 1406 3679 1462
rect 3747 1406 3803 1462
rect 3871 1406 3927 1462
rect 3995 1406 4051 1462
rect 4119 1406 4175 1462
rect 4243 1406 4299 1462
rect 2507 1282 2563 1338
rect 2631 1282 2687 1338
rect 2755 1282 2811 1338
rect 2879 1282 2935 1338
rect 3003 1282 3059 1338
rect 3127 1282 3183 1338
rect 3251 1282 3307 1338
rect 3375 1282 3431 1338
rect 3499 1282 3555 1338
rect 3623 1282 3679 1338
rect 3747 1282 3803 1338
rect 3871 1282 3927 1338
rect 3995 1282 4051 1338
rect 4119 1282 4175 1338
rect 4243 1282 4299 1338
rect 2507 1158 2563 1214
rect 2631 1158 2687 1214
rect 2755 1158 2811 1214
rect 2879 1158 2935 1214
rect 3003 1158 3059 1214
rect 3127 1158 3183 1214
rect 3251 1158 3307 1214
rect 3375 1158 3431 1214
rect 3499 1158 3555 1214
rect 3623 1158 3679 1214
rect 3747 1158 3803 1214
rect 3871 1158 3927 1214
rect 3995 1158 4051 1214
rect 4119 1158 4175 1214
rect 4243 1158 4299 1214
rect 2507 1034 2563 1090
rect 2631 1034 2687 1090
rect 2755 1034 2811 1090
rect 2879 1034 2935 1090
rect 3003 1034 3059 1090
rect 3127 1034 3183 1090
rect 3251 1034 3307 1090
rect 3375 1034 3431 1090
rect 3499 1034 3555 1090
rect 3623 1034 3679 1090
rect 3747 1034 3803 1090
rect 3871 1034 3927 1090
rect 3995 1034 4051 1090
rect 4119 1034 4175 1090
rect 4243 1034 4299 1090
rect 2507 910 2563 966
rect 2631 910 2687 966
rect 2755 910 2811 966
rect 2879 910 2935 966
rect 3003 910 3059 966
rect 3127 910 3183 966
rect 3251 910 3307 966
rect 3375 910 3431 966
rect 3499 910 3555 966
rect 3623 910 3679 966
rect 3747 910 3803 966
rect 3871 910 3927 966
rect 3995 910 4051 966
rect 4119 910 4175 966
rect 4243 910 4299 966
rect 2507 786 2563 842
rect 2631 786 2687 842
rect 2755 786 2811 842
rect 2879 786 2935 842
rect 3003 786 3059 842
rect 3127 786 3183 842
rect 3251 786 3307 842
rect 3375 786 3431 842
rect 3499 786 3555 842
rect 3623 786 3679 842
rect 3747 786 3803 842
rect 3871 786 3927 842
rect 3995 786 4051 842
rect 4119 786 4175 842
rect 4243 786 4299 842
rect 2507 662 2563 718
rect 2631 662 2687 718
rect 2755 662 2811 718
rect 2879 662 2935 718
rect 3003 662 3059 718
rect 3127 662 3183 718
rect 3251 662 3307 718
rect 3375 662 3431 718
rect 3499 662 3555 718
rect 3623 662 3679 718
rect 3747 662 3803 718
rect 3871 662 3927 718
rect 3995 662 4051 718
rect 4119 662 4175 718
rect 4243 662 4299 718
rect 2507 538 2563 594
rect 2631 538 2687 594
rect 2755 538 2811 594
rect 2879 538 2935 594
rect 3003 538 3059 594
rect 3127 538 3183 594
rect 3251 538 3307 594
rect 3375 538 3431 594
rect 3499 538 3555 594
rect 3623 538 3679 594
rect 3747 538 3803 594
rect 3871 538 3927 594
rect 3995 538 4051 594
rect 4119 538 4175 594
rect 4243 538 4299 594
rect 2507 414 2563 470
rect 2631 414 2687 470
rect 2755 414 2811 470
rect 2879 414 2935 470
rect 3003 414 3059 470
rect 3127 414 3183 470
rect 3251 414 3307 470
rect 3375 414 3431 470
rect 3499 414 3555 470
rect 3623 414 3679 470
rect 3747 414 3803 470
rect 3871 414 3927 470
rect 3995 414 4051 470
rect 4119 414 4175 470
rect 4243 414 4299 470
rect 2507 290 2563 346
rect 2631 290 2687 346
rect 2755 290 2811 346
rect 2879 290 2935 346
rect 3003 290 3059 346
rect 3127 290 3183 346
rect 3251 290 3307 346
rect 3375 290 3431 346
rect 3499 290 3555 346
rect 3623 290 3679 346
rect 3747 290 3803 346
rect 3871 290 3927 346
rect 3995 290 4051 346
rect 4119 290 4175 346
rect 4243 290 4299 346
rect 2507 166 2563 222
rect 2631 166 2687 222
rect 2755 166 2811 222
rect 2879 166 2935 222
rect 3003 166 3059 222
rect 3127 166 3183 222
rect 3251 166 3307 222
rect 3375 166 3431 222
rect 3499 166 3555 222
rect 3623 166 3679 222
rect 3747 166 3803 222
rect 3871 166 3927 222
rect 3995 166 4051 222
rect 4119 166 4175 222
rect 4243 166 4299 222
rect 2507 42 2563 98
rect 2631 42 2687 98
rect 2755 42 2811 98
rect 2879 42 2935 98
rect 3003 42 3059 98
rect 3127 42 3183 98
rect 3251 42 3307 98
rect 3375 42 3431 98
rect 3499 42 3555 98
rect 3623 42 3679 98
rect 3747 42 3803 98
rect 3871 42 3927 98
rect 3995 42 4051 98
rect 4119 42 4175 98
rect 4243 42 4299 98
rect 6368 2894 6424 2950
rect 6492 2894 6548 2950
rect 6616 2894 6672 2950
rect 6740 2894 6796 2950
rect 6864 2894 6920 2950
rect 6988 2894 7044 2950
rect 7112 2894 7168 2950
rect 7236 2894 7292 2950
rect 7360 2894 7416 2950
rect 6368 2770 6424 2826
rect 6492 2770 6548 2826
rect 6616 2770 6672 2826
rect 6740 2770 6796 2826
rect 6864 2770 6920 2826
rect 6988 2770 7044 2826
rect 7112 2770 7168 2826
rect 7236 2770 7292 2826
rect 7360 2770 7416 2826
rect 6368 2646 6424 2702
rect 6492 2646 6548 2702
rect 6616 2646 6672 2702
rect 6740 2646 6796 2702
rect 6864 2646 6920 2702
rect 6988 2646 7044 2702
rect 7112 2646 7168 2702
rect 7236 2646 7292 2702
rect 7360 2646 7416 2702
rect 6368 2522 6424 2578
rect 6492 2522 6548 2578
rect 6616 2522 6672 2578
rect 6740 2522 6796 2578
rect 6864 2522 6920 2578
rect 6988 2522 7044 2578
rect 7112 2522 7168 2578
rect 7236 2522 7292 2578
rect 7360 2522 7416 2578
rect 6368 2398 6424 2454
rect 6492 2398 6548 2454
rect 6616 2398 6672 2454
rect 6740 2398 6796 2454
rect 6864 2398 6920 2454
rect 6988 2398 7044 2454
rect 7112 2398 7168 2454
rect 7236 2398 7292 2454
rect 7360 2398 7416 2454
rect 6368 2274 6424 2330
rect 6492 2274 6548 2330
rect 6616 2274 6672 2330
rect 6740 2274 6796 2330
rect 6864 2274 6920 2330
rect 6988 2274 7044 2330
rect 7112 2274 7168 2330
rect 7236 2274 7292 2330
rect 7360 2274 7416 2330
rect 6368 2150 6424 2206
rect 6492 2150 6548 2206
rect 6616 2150 6672 2206
rect 6740 2150 6796 2206
rect 6864 2150 6920 2206
rect 6988 2150 7044 2206
rect 7112 2150 7168 2206
rect 7236 2150 7292 2206
rect 7360 2150 7416 2206
rect 6368 2026 6424 2082
rect 6492 2026 6548 2082
rect 6616 2026 6672 2082
rect 6740 2026 6796 2082
rect 6864 2026 6920 2082
rect 6988 2026 7044 2082
rect 7112 2026 7168 2082
rect 7236 2026 7292 2082
rect 7360 2026 7416 2082
rect 6368 1902 6424 1958
rect 6492 1902 6548 1958
rect 6616 1902 6672 1958
rect 6740 1902 6796 1958
rect 6864 1902 6920 1958
rect 6988 1902 7044 1958
rect 7112 1902 7168 1958
rect 7236 1902 7292 1958
rect 7360 1902 7416 1958
rect 6368 1778 6424 1834
rect 6492 1778 6548 1834
rect 6616 1778 6672 1834
rect 6740 1778 6796 1834
rect 6864 1778 6920 1834
rect 6988 1778 7044 1834
rect 7112 1778 7168 1834
rect 7236 1778 7292 1834
rect 7360 1778 7416 1834
rect 6368 1654 6424 1710
rect 6492 1654 6548 1710
rect 6616 1654 6672 1710
rect 6740 1654 6796 1710
rect 6864 1654 6920 1710
rect 6988 1654 7044 1710
rect 7112 1654 7168 1710
rect 7236 1654 7292 1710
rect 7360 1654 7416 1710
rect 6368 1530 6424 1586
rect 6492 1530 6548 1586
rect 6616 1530 6672 1586
rect 6740 1530 6796 1586
rect 6864 1530 6920 1586
rect 6988 1530 7044 1586
rect 7112 1530 7168 1586
rect 7236 1530 7292 1586
rect 7360 1530 7416 1586
rect 6368 1406 6424 1462
rect 6492 1406 6548 1462
rect 6616 1406 6672 1462
rect 6740 1406 6796 1462
rect 6864 1406 6920 1462
rect 6988 1406 7044 1462
rect 7112 1406 7168 1462
rect 7236 1406 7292 1462
rect 7360 1406 7416 1462
rect 6368 1282 6424 1338
rect 6492 1282 6548 1338
rect 6616 1282 6672 1338
rect 6740 1282 6796 1338
rect 6864 1282 6920 1338
rect 6988 1282 7044 1338
rect 7112 1282 7168 1338
rect 7236 1282 7292 1338
rect 7360 1282 7416 1338
rect 6368 1158 6424 1214
rect 6492 1158 6548 1214
rect 6616 1158 6672 1214
rect 6740 1158 6796 1214
rect 6864 1158 6920 1214
rect 6988 1158 7044 1214
rect 7112 1158 7168 1214
rect 7236 1158 7292 1214
rect 7360 1158 7416 1214
rect 6368 1034 6424 1090
rect 6492 1034 6548 1090
rect 6616 1034 6672 1090
rect 6740 1034 6796 1090
rect 6864 1034 6920 1090
rect 6988 1034 7044 1090
rect 7112 1034 7168 1090
rect 7236 1034 7292 1090
rect 7360 1034 7416 1090
rect 6368 910 6424 966
rect 6492 910 6548 966
rect 6616 910 6672 966
rect 6740 910 6796 966
rect 6864 910 6920 966
rect 6988 910 7044 966
rect 7112 910 7168 966
rect 7236 910 7292 966
rect 7360 910 7416 966
rect 6368 786 6424 842
rect 6492 786 6548 842
rect 6616 786 6672 842
rect 6740 786 6796 842
rect 6864 786 6920 842
rect 6988 786 7044 842
rect 7112 786 7168 842
rect 7236 786 7292 842
rect 7360 786 7416 842
rect 6368 662 6424 718
rect 6492 662 6548 718
rect 6616 662 6672 718
rect 6740 662 6796 718
rect 6864 662 6920 718
rect 6988 662 7044 718
rect 7112 662 7168 718
rect 7236 662 7292 718
rect 7360 662 7416 718
rect 6368 538 6424 594
rect 6492 538 6548 594
rect 6616 538 6672 594
rect 6740 538 6796 594
rect 6864 538 6920 594
rect 6988 538 7044 594
rect 7112 538 7168 594
rect 7236 538 7292 594
rect 7360 538 7416 594
rect 6368 414 6424 470
rect 6492 414 6548 470
rect 6616 414 6672 470
rect 6740 414 6796 470
rect 6864 414 6920 470
rect 6988 414 7044 470
rect 7112 414 7168 470
rect 7236 414 7292 470
rect 7360 414 7416 470
rect 6368 290 6424 346
rect 6492 290 6548 346
rect 6616 290 6672 346
rect 6740 290 6796 346
rect 6864 290 6920 346
rect 6988 290 7044 346
rect 7112 290 7168 346
rect 7236 290 7292 346
rect 7360 290 7416 346
rect 6368 166 6424 222
rect 6492 166 6548 222
rect 6616 166 6672 222
rect 6740 166 6796 222
rect 6864 166 6920 222
rect 6988 166 7044 222
rect 7112 166 7168 222
rect 7236 166 7292 222
rect 7360 166 7416 222
rect 6368 42 6424 98
rect 6492 42 6548 98
rect 6616 42 6672 98
rect 6740 42 6796 98
rect 6864 42 6920 98
rect 6988 42 7044 98
rect 7112 42 7168 98
rect 7236 42 7292 98
rect 7360 42 7416 98
rect 8751 2894 8807 2950
rect 8875 2894 8931 2950
rect 8999 2894 9055 2950
rect 9123 2894 9179 2950
rect 9247 2894 9303 2950
rect 9371 2894 9427 2950
rect 9495 2894 9551 2950
rect 9619 2894 9675 2950
rect 9743 2894 9799 2950
rect 9867 2894 9923 2950
rect 9991 2894 10047 2950
rect 10115 2894 10171 2950
rect 10239 2894 10295 2950
rect 10363 2894 10419 2950
rect 10487 2894 10543 2950
rect 8751 2770 8807 2826
rect 8875 2770 8931 2826
rect 8999 2770 9055 2826
rect 9123 2770 9179 2826
rect 9247 2770 9303 2826
rect 9371 2770 9427 2826
rect 9495 2770 9551 2826
rect 9619 2770 9675 2826
rect 9743 2770 9799 2826
rect 9867 2770 9923 2826
rect 9991 2770 10047 2826
rect 10115 2770 10171 2826
rect 10239 2770 10295 2826
rect 10363 2770 10419 2826
rect 10487 2770 10543 2826
rect 8751 2646 8807 2702
rect 8875 2646 8931 2702
rect 8999 2646 9055 2702
rect 9123 2646 9179 2702
rect 9247 2646 9303 2702
rect 9371 2646 9427 2702
rect 9495 2646 9551 2702
rect 9619 2646 9675 2702
rect 9743 2646 9799 2702
rect 9867 2646 9923 2702
rect 9991 2646 10047 2702
rect 10115 2646 10171 2702
rect 10239 2646 10295 2702
rect 10363 2646 10419 2702
rect 10487 2646 10543 2702
rect 8751 2522 8807 2578
rect 8875 2522 8931 2578
rect 8999 2522 9055 2578
rect 9123 2522 9179 2578
rect 9247 2522 9303 2578
rect 9371 2522 9427 2578
rect 9495 2522 9551 2578
rect 9619 2522 9675 2578
rect 9743 2522 9799 2578
rect 9867 2522 9923 2578
rect 9991 2522 10047 2578
rect 10115 2522 10171 2578
rect 10239 2522 10295 2578
rect 10363 2522 10419 2578
rect 10487 2522 10543 2578
rect 8751 2398 8807 2454
rect 8875 2398 8931 2454
rect 8999 2398 9055 2454
rect 9123 2398 9179 2454
rect 9247 2398 9303 2454
rect 9371 2398 9427 2454
rect 9495 2398 9551 2454
rect 9619 2398 9675 2454
rect 9743 2398 9799 2454
rect 9867 2398 9923 2454
rect 9991 2398 10047 2454
rect 10115 2398 10171 2454
rect 10239 2398 10295 2454
rect 10363 2398 10419 2454
rect 10487 2398 10543 2454
rect 8751 2274 8807 2330
rect 8875 2274 8931 2330
rect 8999 2274 9055 2330
rect 9123 2274 9179 2330
rect 9247 2274 9303 2330
rect 9371 2274 9427 2330
rect 9495 2274 9551 2330
rect 9619 2274 9675 2330
rect 9743 2274 9799 2330
rect 9867 2274 9923 2330
rect 9991 2274 10047 2330
rect 10115 2274 10171 2330
rect 10239 2274 10295 2330
rect 10363 2274 10419 2330
rect 10487 2274 10543 2330
rect 8751 2150 8807 2206
rect 8875 2150 8931 2206
rect 8999 2150 9055 2206
rect 9123 2150 9179 2206
rect 9247 2150 9303 2206
rect 9371 2150 9427 2206
rect 9495 2150 9551 2206
rect 9619 2150 9675 2206
rect 9743 2150 9799 2206
rect 9867 2150 9923 2206
rect 9991 2150 10047 2206
rect 10115 2150 10171 2206
rect 10239 2150 10295 2206
rect 10363 2150 10419 2206
rect 10487 2150 10543 2206
rect 8751 2026 8807 2082
rect 8875 2026 8931 2082
rect 8999 2026 9055 2082
rect 9123 2026 9179 2082
rect 9247 2026 9303 2082
rect 9371 2026 9427 2082
rect 9495 2026 9551 2082
rect 9619 2026 9675 2082
rect 9743 2026 9799 2082
rect 9867 2026 9923 2082
rect 9991 2026 10047 2082
rect 10115 2026 10171 2082
rect 10239 2026 10295 2082
rect 10363 2026 10419 2082
rect 10487 2026 10543 2082
rect 8751 1902 8807 1958
rect 8875 1902 8931 1958
rect 8999 1902 9055 1958
rect 9123 1902 9179 1958
rect 9247 1902 9303 1958
rect 9371 1902 9427 1958
rect 9495 1902 9551 1958
rect 9619 1902 9675 1958
rect 9743 1902 9799 1958
rect 9867 1902 9923 1958
rect 9991 1902 10047 1958
rect 10115 1902 10171 1958
rect 10239 1902 10295 1958
rect 10363 1902 10419 1958
rect 10487 1902 10543 1958
rect 8751 1778 8807 1834
rect 8875 1778 8931 1834
rect 8999 1778 9055 1834
rect 9123 1778 9179 1834
rect 9247 1778 9303 1834
rect 9371 1778 9427 1834
rect 9495 1778 9551 1834
rect 9619 1778 9675 1834
rect 9743 1778 9799 1834
rect 9867 1778 9923 1834
rect 9991 1778 10047 1834
rect 10115 1778 10171 1834
rect 10239 1778 10295 1834
rect 10363 1778 10419 1834
rect 10487 1778 10543 1834
rect 8751 1654 8807 1710
rect 8875 1654 8931 1710
rect 8999 1654 9055 1710
rect 9123 1654 9179 1710
rect 9247 1654 9303 1710
rect 9371 1654 9427 1710
rect 9495 1654 9551 1710
rect 9619 1654 9675 1710
rect 9743 1654 9799 1710
rect 9867 1654 9923 1710
rect 9991 1654 10047 1710
rect 10115 1654 10171 1710
rect 10239 1654 10295 1710
rect 10363 1654 10419 1710
rect 10487 1654 10543 1710
rect 8751 1530 8807 1586
rect 8875 1530 8931 1586
rect 8999 1530 9055 1586
rect 9123 1530 9179 1586
rect 9247 1530 9303 1586
rect 9371 1530 9427 1586
rect 9495 1530 9551 1586
rect 9619 1530 9675 1586
rect 9743 1530 9799 1586
rect 9867 1530 9923 1586
rect 9991 1530 10047 1586
rect 10115 1530 10171 1586
rect 10239 1530 10295 1586
rect 10363 1530 10419 1586
rect 10487 1530 10543 1586
rect 8751 1406 8807 1462
rect 8875 1406 8931 1462
rect 8999 1406 9055 1462
rect 9123 1406 9179 1462
rect 9247 1406 9303 1462
rect 9371 1406 9427 1462
rect 9495 1406 9551 1462
rect 9619 1406 9675 1462
rect 9743 1406 9799 1462
rect 9867 1406 9923 1462
rect 9991 1406 10047 1462
rect 10115 1406 10171 1462
rect 10239 1406 10295 1462
rect 10363 1406 10419 1462
rect 10487 1406 10543 1462
rect 8751 1282 8807 1338
rect 8875 1282 8931 1338
rect 8999 1282 9055 1338
rect 9123 1282 9179 1338
rect 9247 1282 9303 1338
rect 9371 1282 9427 1338
rect 9495 1282 9551 1338
rect 9619 1282 9675 1338
rect 9743 1282 9799 1338
rect 9867 1282 9923 1338
rect 9991 1282 10047 1338
rect 10115 1282 10171 1338
rect 10239 1282 10295 1338
rect 10363 1282 10419 1338
rect 10487 1282 10543 1338
rect 8751 1158 8807 1214
rect 8875 1158 8931 1214
rect 8999 1158 9055 1214
rect 9123 1158 9179 1214
rect 9247 1158 9303 1214
rect 9371 1158 9427 1214
rect 9495 1158 9551 1214
rect 9619 1158 9675 1214
rect 9743 1158 9799 1214
rect 9867 1158 9923 1214
rect 9991 1158 10047 1214
rect 10115 1158 10171 1214
rect 10239 1158 10295 1214
rect 10363 1158 10419 1214
rect 10487 1158 10543 1214
rect 8751 1034 8807 1090
rect 8875 1034 8931 1090
rect 8999 1034 9055 1090
rect 9123 1034 9179 1090
rect 9247 1034 9303 1090
rect 9371 1034 9427 1090
rect 9495 1034 9551 1090
rect 9619 1034 9675 1090
rect 9743 1034 9799 1090
rect 9867 1034 9923 1090
rect 9991 1034 10047 1090
rect 10115 1034 10171 1090
rect 10239 1034 10295 1090
rect 10363 1034 10419 1090
rect 10487 1034 10543 1090
rect 8751 910 8807 966
rect 8875 910 8931 966
rect 8999 910 9055 966
rect 9123 910 9179 966
rect 9247 910 9303 966
rect 9371 910 9427 966
rect 9495 910 9551 966
rect 9619 910 9675 966
rect 9743 910 9799 966
rect 9867 910 9923 966
rect 9991 910 10047 966
rect 10115 910 10171 966
rect 10239 910 10295 966
rect 10363 910 10419 966
rect 10487 910 10543 966
rect 8751 786 8807 842
rect 8875 786 8931 842
rect 8999 786 9055 842
rect 9123 786 9179 842
rect 9247 786 9303 842
rect 9371 786 9427 842
rect 9495 786 9551 842
rect 9619 786 9675 842
rect 9743 786 9799 842
rect 9867 786 9923 842
rect 9991 786 10047 842
rect 10115 786 10171 842
rect 10239 786 10295 842
rect 10363 786 10419 842
rect 10487 786 10543 842
rect 8751 662 8807 718
rect 8875 662 8931 718
rect 8999 662 9055 718
rect 9123 662 9179 718
rect 9247 662 9303 718
rect 9371 662 9427 718
rect 9495 662 9551 718
rect 9619 662 9675 718
rect 9743 662 9799 718
rect 9867 662 9923 718
rect 9991 662 10047 718
rect 10115 662 10171 718
rect 10239 662 10295 718
rect 10363 662 10419 718
rect 10487 662 10543 718
rect 8751 538 8807 594
rect 8875 538 8931 594
rect 8999 538 9055 594
rect 9123 538 9179 594
rect 9247 538 9303 594
rect 9371 538 9427 594
rect 9495 538 9551 594
rect 9619 538 9675 594
rect 9743 538 9799 594
rect 9867 538 9923 594
rect 9991 538 10047 594
rect 10115 538 10171 594
rect 10239 538 10295 594
rect 10363 538 10419 594
rect 10487 538 10543 594
rect 8751 414 8807 470
rect 8875 414 8931 470
rect 8999 414 9055 470
rect 9123 414 9179 470
rect 9247 414 9303 470
rect 9371 414 9427 470
rect 9495 414 9551 470
rect 9619 414 9675 470
rect 9743 414 9799 470
rect 9867 414 9923 470
rect 9991 414 10047 470
rect 10115 414 10171 470
rect 10239 414 10295 470
rect 10363 414 10419 470
rect 10487 414 10543 470
rect 8751 290 8807 346
rect 8875 290 8931 346
rect 8999 290 9055 346
rect 9123 290 9179 346
rect 9247 290 9303 346
rect 9371 290 9427 346
rect 9495 290 9551 346
rect 9619 290 9675 346
rect 9743 290 9799 346
rect 9867 290 9923 346
rect 9991 290 10047 346
rect 10115 290 10171 346
rect 10239 290 10295 346
rect 10363 290 10419 346
rect 10487 290 10543 346
rect 8751 166 8807 222
rect 8875 166 8931 222
rect 8999 166 9055 222
rect 9123 166 9179 222
rect 9247 166 9303 222
rect 9371 166 9427 222
rect 9495 166 9551 222
rect 9619 166 9675 222
rect 9743 166 9799 222
rect 9867 166 9923 222
rect 9991 166 10047 222
rect 10115 166 10171 222
rect 10239 166 10295 222
rect 10363 166 10419 222
rect 10487 166 10543 222
rect 8751 42 8807 98
rect 8875 42 8931 98
rect 8999 42 9055 98
rect 9123 42 9179 98
rect 9247 42 9303 98
rect 9371 42 9427 98
rect 9495 42 9551 98
rect 9619 42 9675 98
rect 9743 42 9799 98
rect 9867 42 9923 98
rect 9991 42 10047 98
rect 10115 42 10171 98
rect 10239 42 10295 98
rect 10363 42 10419 98
rect 10487 42 10543 98
rect 12852 2894 12908 2950
rect 12976 2894 13032 2950
rect 13100 2894 13156 2950
rect 13224 2894 13280 2950
rect 13348 2894 13404 2950
rect 13472 2894 13528 2950
rect 13596 2894 13652 2950
rect 13720 2894 13776 2950
rect 13844 2894 13900 2950
rect 12852 2770 12908 2826
rect 12976 2770 13032 2826
rect 13100 2770 13156 2826
rect 13224 2770 13280 2826
rect 13348 2770 13404 2826
rect 13472 2770 13528 2826
rect 13596 2770 13652 2826
rect 13720 2770 13776 2826
rect 13844 2770 13900 2826
rect 12852 2646 12908 2702
rect 12976 2646 13032 2702
rect 13100 2646 13156 2702
rect 13224 2646 13280 2702
rect 13348 2646 13404 2702
rect 13472 2646 13528 2702
rect 13596 2646 13652 2702
rect 13720 2646 13776 2702
rect 13844 2646 13900 2702
rect 12852 2522 12908 2578
rect 12976 2522 13032 2578
rect 13100 2522 13156 2578
rect 13224 2522 13280 2578
rect 13348 2522 13404 2578
rect 13472 2522 13528 2578
rect 13596 2522 13652 2578
rect 13720 2522 13776 2578
rect 13844 2522 13900 2578
rect 12852 2398 12908 2454
rect 12976 2398 13032 2454
rect 13100 2398 13156 2454
rect 13224 2398 13280 2454
rect 13348 2398 13404 2454
rect 13472 2398 13528 2454
rect 13596 2398 13652 2454
rect 13720 2398 13776 2454
rect 13844 2398 13900 2454
rect 12852 2274 12908 2330
rect 12976 2274 13032 2330
rect 13100 2274 13156 2330
rect 13224 2274 13280 2330
rect 13348 2274 13404 2330
rect 13472 2274 13528 2330
rect 13596 2274 13652 2330
rect 13720 2274 13776 2330
rect 13844 2274 13900 2330
rect 12852 2150 12908 2206
rect 12976 2150 13032 2206
rect 13100 2150 13156 2206
rect 13224 2150 13280 2206
rect 13348 2150 13404 2206
rect 13472 2150 13528 2206
rect 13596 2150 13652 2206
rect 13720 2150 13776 2206
rect 13844 2150 13900 2206
rect 12852 2026 12908 2082
rect 12976 2026 13032 2082
rect 13100 2026 13156 2082
rect 13224 2026 13280 2082
rect 13348 2026 13404 2082
rect 13472 2026 13528 2082
rect 13596 2026 13652 2082
rect 13720 2026 13776 2082
rect 13844 2026 13900 2082
rect 12852 1902 12908 1958
rect 12976 1902 13032 1958
rect 13100 1902 13156 1958
rect 13224 1902 13280 1958
rect 13348 1902 13404 1958
rect 13472 1902 13528 1958
rect 13596 1902 13652 1958
rect 13720 1902 13776 1958
rect 13844 1902 13900 1958
rect 12852 1778 12908 1834
rect 12976 1778 13032 1834
rect 13100 1778 13156 1834
rect 13224 1778 13280 1834
rect 13348 1778 13404 1834
rect 13472 1778 13528 1834
rect 13596 1778 13652 1834
rect 13720 1778 13776 1834
rect 13844 1778 13900 1834
rect 12852 1654 12908 1710
rect 12976 1654 13032 1710
rect 13100 1654 13156 1710
rect 13224 1654 13280 1710
rect 13348 1654 13404 1710
rect 13472 1654 13528 1710
rect 13596 1654 13652 1710
rect 13720 1654 13776 1710
rect 13844 1654 13900 1710
rect 12852 1530 12908 1586
rect 12976 1530 13032 1586
rect 13100 1530 13156 1586
rect 13224 1530 13280 1586
rect 13348 1530 13404 1586
rect 13472 1530 13528 1586
rect 13596 1530 13652 1586
rect 13720 1530 13776 1586
rect 13844 1530 13900 1586
rect 12852 1406 12908 1462
rect 12976 1406 13032 1462
rect 13100 1406 13156 1462
rect 13224 1406 13280 1462
rect 13348 1406 13404 1462
rect 13472 1406 13528 1462
rect 13596 1406 13652 1462
rect 13720 1406 13776 1462
rect 13844 1406 13900 1462
rect 12852 1282 12908 1338
rect 12976 1282 13032 1338
rect 13100 1282 13156 1338
rect 13224 1282 13280 1338
rect 13348 1282 13404 1338
rect 13472 1282 13528 1338
rect 13596 1282 13652 1338
rect 13720 1282 13776 1338
rect 13844 1282 13900 1338
rect 12852 1158 12908 1214
rect 12976 1158 13032 1214
rect 13100 1158 13156 1214
rect 13224 1158 13280 1214
rect 13348 1158 13404 1214
rect 13472 1158 13528 1214
rect 13596 1158 13652 1214
rect 13720 1158 13776 1214
rect 13844 1158 13900 1214
rect 12852 1034 12908 1090
rect 12976 1034 13032 1090
rect 13100 1034 13156 1090
rect 13224 1034 13280 1090
rect 13348 1034 13404 1090
rect 13472 1034 13528 1090
rect 13596 1034 13652 1090
rect 13720 1034 13776 1090
rect 13844 1034 13900 1090
rect 12852 910 12908 966
rect 12976 910 13032 966
rect 13100 910 13156 966
rect 13224 910 13280 966
rect 13348 910 13404 966
rect 13472 910 13528 966
rect 13596 910 13652 966
rect 13720 910 13776 966
rect 13844 910 13900 966
rect 12852 786 12908 842
rect 12976 786 13032 842
rect 13100 786 13156 842
rect 13224 786 13280 842
rect 13348 786 13404 842
rect 13472 786 13528 842
rect 13596 786 13652 842
rect 13720 786 13776 842
rect 13844 786 13900 842
rect 12852 662 12908 718
rect 12976 662 13032 718
rect 13100 662 13156 718
rect 13224 662 13280 718
rect 13348 662 13404 718
rect 13472 662 13528 718
rect 13596 662 13652 718
rect 13720 662 13776 718
rect 13844 662 13900 718
rect 12852 538 12908 594
rect 12976 538 13032 594
rect 13100 538 13156 594
rect 13224 538 13280 594
rect 13348 538 13404 594
rect 13472 538 13528 594
rect 13596 538 13652 594
rect 13720 538 13776 594
rect 13844 538 13900 594
rect 12852 414 12908 470
rect 12976 414 13032 470
rect 13100 414 13156 470
rect 13224 414 13280 470
rect 13348 414 13404 470
rect 13472 414 13528 470
rect 13596 414 13652 470
rect 13720 414 13776 470
rect 13844 414 13900 470
rect 12852 290 12908 346
rect 12976 290 13032 346
rect 13100 290 13156 346
rect 13224 290 13280 346
rect 13348 290 13404 346
rect 13472 290 13528 346
rect 13596 290 13652 346
rect 13720 290 13776 346
rect 13844 290 13900 346
rect 12852 166 12908 222
rect 12976 166 13032 222
rect 13100 166 13156 222
rect 13224 166 13280 222
rect 13348 166 13404 222
rect 13472 166 13528 222
rect 13596 166 13652 222
rect 13720 166 13776 222
rect 13844 166 13900 222
rect 12852 42 12908 98
rect 12976 42 13032 98
rect 13100 42 13156 98
rect 13224 42 13280 98
rect 13348 42 13404 98
rect 13472 42 13528 98
rect 13596 42 13652 98
rect 13720 42 13776 98
rect 13844 42 13900 98
<< metal3 >>
rect 14757 50972 14833 50982
rect 14757 49620 14767 50972
rect 14823 49620 14833 50972
rect 14757 49610 14833 49620
rect 6384 46670 6460 46680
rect 6384 46614 6394 46670
rect 6450 46614 6460 46670
rect 6384 46546 6460 46614
rect 6384 46490 6394 46546
rect 6450 46490 6460 46546
rect 6384 46422 6460 46490
rect 6384 46366 6394 46422
rect 6450 46366 6460 46422
rect 4460 46323 4536 46333
rect 4460 46267 4470 46323
rect 4526 46267 4536 46323
rect 4460 46199 4536 46267
rect 6384 46298 6460 46366
rect 6384 46242 6394 46298
rect 6450 46242 6460 46298
rect 4460 46143 4470 46199
rect 4526 46143 4536 46199
rect 4460 46075 4536 46143
rect 4460 46019 4470 46075
rect 4526 46019 4536 46075
rect 4460 45951 4536 46019
rect 4460 45895 4470 45951
rect 4526 45895 4536 45951
rect 4460 45827 4536 45895
rect 4460 45771 4470 45827
rect 4526 45771 4536 45827
rect 4460 45703 4536 45771
rect 4460 45647 4470 45703
rect 4526 45647 4536 45703
rect 4460 45579 4536 45647
rect 4460 45523 4470 45579
rect 4526 45523 4536 45579
rect 4460 45455 4536 45523
rect 4460 45399 4470 45455
rect 4526 45399 4536 45455
rect 4460 45331 4536 45399
rect 4460 45275 4470 45331
rect 4526 45275 4536 45331
rect 1094 45255 1170 45265
rect 1094 45199 1104 45255
rect 1160 45199 1170 45255
rect 1094 45131 1170 45199
rect 4460 45207 4536 45275
rect 4460 45151 4470 45207
rect 4526 45151 4536 45207
rect 1094 45075 1104 45131
rect 1160 45075 1170 45131
rect 1094 45007 1170 45075
rect 1094 44951 1104 45007
rect 1160 44951 1170 45007
rect 1094 44883 1170 44951
rect 1094 44827 1104 44883
rect 1160 44827 1170 44883
rect 1094 44759 1170 44827
rect 1094 44703 1104 44759
rect 1160 44703 1170 44759
rect 1094 44635 1170 44703
rect 1094 44579 1104 44635
rect 1160 44579 1170 44635
rect 1094 44511 1170 44579
rect 1094 44455 1104 44511
rect 1160 44455 1170 44511
rect 1094 44387 1170 44455
rect 1094 44331 1104 44387
rect 1160 44331 1170 44387
rect 1094 44263 1170 44331
rect 1094 44207 1104 44263
rect 1160 44207 1170 44263
rect 1094 44139 1170 44207
rect 1094 44083 1104 44139
rect 1160 44083 1170 44139
rect 1094 44015 1170 44083
rect 1094 43959 1104 44015
rect 1160 43959 1170 44015
rect 1094 43891 1170 43959
rect 1094 43835 1104 43891
rect 1160 43835 1170 43891
rect 1094 43767 1170 43835
rect 1094 43711 1104 43767
rect 1160 43711 1170 43767
rect 1094 43643 1170 43711
rect 1094 43587 1104 43643
rect 1160 43587 1170 43643
rect 1094 43519 1170 43587
rect 1094 43463 1104 43519
rect 1160 43463 1170 43519
rect 1094 43453 1170 43463
rect 1218 45131 1294 45141
rect 1218 45075 1228 45131
rect 1284 45075 1294 45131
rect 1218 45007 1294 45075
rect 4460 45083 4536 45151
rect 4460 45027 4470 45083
rect 4526 45027 4536 45083
rect 1218 44951 1228 45007
rect 1284 44951 1294 45007
rect 1218 44883 1294 44951
rect 1218 44827 1228 44883
rect 1284 44827 1294 44883
rect 1218 44759 1294 44827
rect 1218 44703 1228 44759
rect 1284 44703 1294 44759
rect 1218 44635 1294 44703
rect 1218 44579 1228 44635
rect 1284 44579 1294 44635
rect 1218 44511 1294 44579
rect 1218 44455 1228 44511
rect 1284 44455 1294 44511
rect 1218 44387 1294 44455
rect 1218 44331 1228 44387
rect 1284 44331 1294 44387
rect 1218 44263 1294 44331
rect 1218 44207 1228 44263
rect 1284 44207 1294 44263
rect 1218 44139 1294 44207
rect 1218 44083 1228 44139
rect 1284 44083 1294 44139
rect 1218 44015 1294 44083
rect 1218 43959 1228 44015
rect 1284 43959 1294 44015
rect 1218 43891 1294 43959
rect 1218 43835 1228 43891
rect 1284 43835 1294 43891
rect 1218 43767 1294 43835
rect 1218 43711 1228 43767
rect 1284 43711 1294 43767
rect 1218 43643 1294 43711
rect 1218 43587 1228 43643
rect 1284 43587 1294 43643
rect 1218 43519 1294 43587
rect 1218 43463 1228 43519
rect 1284 43463 1294 43519
rect 1218 43395 1294 43463
rect 1218 43339 1228 43395
rect 1284 43339 1294 43395
rect 1218 43329 1294 43339
rect 1342 45007 1418 45017
rect 1342 44951 1352 45007
rect 1408 44951 1418 45007
rect 1342 44883 1418 44951
rect 4460 44959 4536 45027
rect 4460 44903 4470 44959
rect 4526 44903 4536 44959
rect 1342 44827 1352 44883
rect 1408 44827 1418 44883
rect 1342 44759 1418 44827
rect 1342 44703 1352 44759
rect 1408 44703 1418 44759
rect 1342 44635 1418 44703
rect 1342 44579 1352 44635
rect 1408 44579 1418 44635
rect 1342 44511 1418 44579
rect 1342 44455 1352 44511
rect 1408 44455 1418 44511
rect 1342 44387 1418 44455
rect 1342 44331 1352 44387
rect 1408 44331 1418 44387
rect 1342 44263 1418 44331
rect 1342 44207 1352 44263
rect 1408 44207 1418 44263
rect 1342 44139 1418 44207
rect 1342 44083 1352 44139
rect 1408 44083 1418 44139
rect 1342 44015 1418 44083
rect 1342 43959 1352 44015
rect 1408 43959 1418 44015
rect 1342 43891 1418 43959
rect 1342 43835 1352 43891
rect 1408 43835 1418 43891
rect 1342 43767 1418 43835
rect 1342 43711 1352 43767
rect 1408 43711 1418 43767
rect 1342 43643 1418 43711
rect 1342 43587 1352 43643
rect 1408 43587 1418 43643
rect 1342 43519 1418 43587
rect 1342 43463 1352 43519
rect 1408 43463 1418 43519
rect 1342 43395 1418 43463
rect 1342 43339 1352 43395
rect 1408 43339 1418 43395
rect 1342 43271 1418 43339
rect 1342 43215 1352 43271
rect 1408 43215 1418 43271
rect 1342 43205 1418 43215
rect 1466 44883 1542 44893
rect 1466 44827 1476 44883
rect 1532 44827 1542 44883
rect 1466 44759 1542 44827
rect 4460 44835 4536 44903
rect 4460 44779 4470 44835
rect 4526 44779 4536 44835
rect 1466 44703 1476 44759
rect 1532 44703 1542 44759
rect 1466 44635 1542 44703
rect 1466 44579 1476 44635
rect 1532 44579 1542 44635
rect 1466 44511 1542 44579
rect 1466 44455 1476 44511
rect 1532 44455 1542 44511
rect 1466 44387 1542 44455
rect 1466 44331 1476 44387
rect 1532 44331 1542 44387
rect 1466 44263 1542 44331
rect 1466 44207 1476 44263
rect 1532 44207 1542 44263
rect 1466 44139 1542 44207
rect 1466 44083 1476 44139
rect 1532 44083 1542 44139
rect 1466 44015 1542 44083
rect 1466 43959 1476 44015
rect 1532 43959 1542 44015
rect 1466 43891 1542 43959
rect 1466 43835 1476 43891
rect 1532 43835 1542 43891
rect 1466 43767 1542 43835
rect 1466 43711 1476 43767
rect 1532 43711 1542 43767
rect 1466 43643 1542 43711
rect 1466 43587 1476 43643
rect 1532 43587 1542 43643
rect 1466 43519 1542 43587
rect 1466 43463 1476 43519
rect 1532 43463 1542 43519
rect 1466 43395 1542 43463
rect 1466 43339 1476 43395
rect 1532 43339 1542 43395
rect 1466 43271 1542 43339
rect 1466 43215 1476 43271
rect 1532 43215 1542 43271
rect 1466 43147 1542 43215
rect 1466 43091 1476 43147
rect 1532 43091 1542 43147
rect 1466 43081 1542 43091
rect 1590 44759 1666 44769
rect 1590 44703 1600 44759
rect 1656 44703 1666 44759
rect 1590 44635 1666 44703
rect 4460 44711 4536 44779
rect 4460 44655 4470 44711
rect 4526 44655 4536 44711
rect 4460 44645 4536 44655
rect 4584 46199 4660 46209
rect 4584 46143 4594 46199
rect 4650 46143 4660 46199
rect 4584 46075 4660 46143
rect 6384 46174 6460 46242
rect 6384 46118 6394 46174
rect 6450 46118 6460 46174
rect 4584 46019 4594 46075
rect 4650 46019 4660 46075
rect 4584 45951 4660 46019
rect 4584 45895 4594 45951
rect 4650 45895 4660 45951
rect 4584 45827 4660 45895
rect 4584 45771 4594 45827
rect 4650 45771 4660 45827
rect 4584 45703 4660 45771
rect 4584 45647 4594 45703
rect 4650 45647 4660 45703
rect 4584 45579 4660 45647
rect 4584 45523 4594 45579
rect 4650 45523 4660 45579
rect 4584 45455 4660 45523
rect 4584 45399 4594 45455
rect 4650 45399 4660 45455
rect 4584 45331 4660 45399
rect 4584 45275 4594 45331
rect 4650 45275 4660 45331
rect 4584 45207 4660 45275
rect 4584 45151 4594 45207
rect 4650 45151 4660 45207
rect 4584 45083 4660 45151
rect 4584 45027 4594 45083
rect 4650 45027 4660 45083
rect 4584 44959 4660 45027
rect 4584 44903 4594 44959
rect 4650 44903 4660 44959
rect 4584 44835 4660 44903
rect 4584 44779 4594 44835
rect 4650 44779 4660 44835
rect 4584 44711 4660 44779
rect 4584 44655 4594 44711
rect 4650 44655 4660 44711
rect 1590 44579 1600 44635
rect 1656 44579 1666 44635
rect 1590 44511 1666 44579
rect 1590 44455 1600 44511
rect 1656 44455 1666 44511
rect 1590 44387 1666 44455
rect 1590 44331 1600 44387
rect 1656 44331 1666 44387
rect 1590 44263 1666 44331
rect 1590 44207 1600 44263
rect 1656 44207 1666 44263
rect 1590 44139 1666 44207
rect 1590 44083 1600 44139
rect 1656 44083 1666 44139
rect 1590 44015 1666 44083
rect 1590 43959 1600 44015
rect 1656 43959 1666 44015
rect 1590 43891 1666 43959
rect 1590 43835 1600 43891
rect 1656 43835 1666 43891
rect 1590 43767 1666 43835
rect 1590 43711 1600 43767
rect 1656 43711 1666 43767
rect 1590 43643 1666 43711
rect 1590 43587 1600 43643
rect 1656 43587 1666 43643
rect 1590 43519 1666 43587
rect 1590 43463 1600 43519
rect 1656 43463 1666 43519
rect 1590 43395 1666 43463
rect 1590 43339 1600 43395
rect 1656 43339 1666 43395
rect 1590 43271 1666 43339
rect 1590 43215 1600 43271
rect 1656 43215 1666 43271
rect 1590 43147 1666 43215
rect 1590 43091 1600 43147
rect 1656 43091 1666 43147
rect 1590 43023 1666 43091
rect 1590 42967 1600 43023
rect 1656 42967 1666 43023
rect 1590 42957 1666 42967
rect 1714 44635 1790 44645
rect 1714 44579 1724 44635
rect 1780 44579 1790 44635
rect 1714 44511 1790 44579
rect 4584 44587 4660 44655
rect 4584 44531 4594 44587
rect 4650 44531 4660 44587
rect 4584 44521 4660 44531
rect 4708 46075 4784 46085
rect 4708 46019 4718 46075
rect 4774 46019 4784 46075
rect 4708 45951 4784 46019
rect 6384 46050 6460 46118
rect 6384 45994 6394 46050
rect 6450 45994 6460 46050
rect 4708 45895 4718 45951
rect 4774 45895 4784 45951
rect 4708 45827 4784 45895
rect 4708 45771 4718 45827
rect 4774 45771 4784 45827
rect 4708 45703 4784 45771
rect 4708 45647 4718 45703
rect 4774 45647 4784 45703
rect 4708 45579 4784 45647
rect 4708 45523 4718 45579
rect 4774 45523 4784 45579
rect 4708 45455 4784 45523
rect 4708 45399 4718 45455
rect 4774 45399 4784 45455
rect 4708 45331 4784 45399
rect 4708 45275 4718 45331
rect 4774 45275 4784 45331
rect 4708 45207 4784 45275
rect 4708 45151 4718 45207
rect 4774 45151 4784 45207
rect 4708 45083 4784 45151
rect 4708 45027 4718 45083
rect 4774 45027 4784 45083
rect 4708 44959 4784 45027
rect 4708 44903 4718 44959
rect 4774 44903 4784 44959
rect 4708 44835 4784 44903
rect 4708 44779 4718 44835
rect 4774 44779 4784 44835
rect 4708 44711 4784 44779
rect 4708 44655 4718 44711
rect 4774 44655 4784 44711
rect 4708 44587 4784 44655
rect 4708 44531 4718 44587
rect 4774 44531 4784 44587
rect 1714 44455 1724 44511
rect 1780 44455 1790 44511
rect 1714 44387 1790 44455
rect 1714 44331 1724 44387
rect 1780 44331 1790 44387
rect 1714 44263 1790 44331
rect 1714 44207 1724 44263
rect 1780 44207 1790 44263
rect 1714 44139 1790 44207
rect 1714 44083 1724 44139
rect 1780 44083 1790 44139
rect 1714 44015 1790 44083
rect 1714 43959 1724 44015
rect 1780 43959 1790 44015
rect 1714 43891 1790 43959
rect 1714 43835 1724 43891
rect 1780 43835 1790 43891
rect 1714 43767 1790 43835
rect 1714 43711 1724 43767
rect 1780 43711 1790 43767
rect 1714 43643 1790 43711
rect 1714 43587 1724 43643
rect 1780 43587 1790 43643
rect 1714 43519 1790 43587
rect 1714 43463 1724 43519
rect 1780 43463 1790 43519
rect 1714 43395 1790 43463
rect 1714 43339 1724 43395
rect 1780 43339 1790 43395
rect 1714 43271 1790 43339
rect 1714 43215 1724 43271
rect 1780 43215 1790 43271
rect 1714 43147 1790 43215
rect 1714 43091 1724 43147
rect 1780 43091 1790 43147
rect 1714 43023 1790 43091
rect 1714 42967 1724 43023
rect 1780 42967 1790 43023
rect 1714 42899 1790 42967
rect 1714 42843 1724 42899
rect 1780 42843 1790 42899
rect 1714 42833 1790 42843
rect 1838 44511 1914 44521
rect 1838 44455 1848 44511
rect 1904 44455 1914 44511
rect 1838 44387 1914 44455
rect 4708 44463 4784 44531
rect 4708 44407 4718 44463
rect 4774 44407 4784 44463
rect 4708 44397 4784 44407
rect 4832 45951 4908 45961
rect 4832 45895 4842 45951
rect 4898 45895 4908 45951
rect 4832 45827 4908 45895
rect 6384 45926 6460 45994
rect 6384 45870 6394 45926
rect 6450 45870 6460 45926
rect 4832 45771 4842 45827
rect 4898 45771 4908 45827
rect 4832 45703 4908 45771
rect 4832 45647 4842 45703
rect 4898 45647 4908 45703
rect 4832 45579 4908 45647
rect 4832 45523 4842 45579
rect 4898 45523 4908 45579
rect 4832 45455 4908 45523
rect 4832 45399 4842 45455
rect 4898 45399 4908 45455
rect 4832 45331 4908 45399
rect 4832 45275 4842 45331
rect 4898 45275 4908 45331
rect 4832 45207 4908 45275
rect 4832 45151 4842 45207
rect 4898 45151 4908 45207
rect 4832 45083 4908 45151
rect 4832 45027 4842 45083
rect 4898 45027 4908 45083
rect 4832 44959 4908 45027
rect 4832 44903 4842 44959
rect 4898 44903 4908 44959
rect 4832 44835 4908 44903
rect 4832 44779 4842 44835
rect 4898 44779 4908 44835
rect 4832 44711 4908 44779
rect 4832 44655 4842 44711
rect 4898 44655 4908 44711
rect 4832 44587 4908 44655
rect 4832 44531 4842 44587
rect 4898 44531 4908 44587
rect 4832 44463 4908 44531
rect 4832 44407 4842 44463
rect 4898 44407 4908 44463
rect 1838 44331 1848 44387
rect 1904 44331 1914 44387
rect 1838 44263 1914 44331
rect 1838 44207 1848 44263
rect 1904 44207 1914 44263
rect 1838 44139 1914 44207
rect 1838 44083 1848 44139
rect 1904 44083 1914 44139
rect 1838 44015 1914 44083
rect 1838 43959 1848 44015
rect 1904 43959 1914 44015
rect 1838 43891 1914 43959
rect 1838 43835 1848 43891
rect 1904 43835 1914 43891
rect 1838 43767 1914 43835
rect 1838 43711 1848 43767
rect 1904 43711 1914 43767
rect 1838 43643 1914 43711
rect 1838 43587 1848 43643
rect 1904 43587 1914 43643
rect 1838 43519 1914 43587
rect 1838 43463 1848 43519
rect 1904 43463 1914 43519
rect 1838 43395 1914 43463
rect 1838 43339 1848 43395
rect 1904 43339 1914 43395
rect 1838 43271 1914 43339
rect 1838 43215 1848 43271
rect 1904 43215 1914 43271
rect 1838 43147 1914 43215
rect 1838 43091 1848 43147
rect 1904 43091 1914 43147
rect 1838 43023 1914 43091
rect 1838 42967 1848 43023
rect 1904 42967 1914 43023
rect 1838 42899 1914 42967
rect 1838 42843 1848 42899
rect 1904 42843 1914 42899
rect 1838 42775 1914 42843
rect 1838 42719 1848 42775
rect 1904 42719 1914 42775
rect 1838 42709 1914 42719
rect 1962 44387 2038 44397
rect 1962 44331 1972 44387
rect 2028 44331 2038 44387
rect 1962 44263 2038 44331
rect 4832 44339 4908 44407
rect 4832 44283 4842 44339
rect 4898 44283 4908 44339
rect 4832 44273 4908 44283
rect 4956 45827 5032 45837
rect 4956 45771 4966 45827
rect 5022 45771 5032 45827
rect 4956 45703 5032 45771
rect 6384 45802 6460 45870
rect 6384 45746 6394 45802
rect 6450 45746 6460 45802
rect 4956 45647 4966 45703
rect 5022 45647 5032 45703
rect 4956 45579 5032 45647
rect 4956 45523 4966 45579
rect 5022 45523 5032 45579
rect 4956 45455 5032 45523
rect 4956 45399 4966 45455
rect 5022 45399 5032 45455
rect 4956 45331 5032 45399
rect 4956 45275 4966 45331
rect 5022 45275 5032 45331
rect 4956 45207 5032 45275
rect 4956 45151 4966 45207
rect 5022 45151 5032 45207
rect 4956 45083 5032 45151
rect 4956 45027 4966 45083
rect 5022 45027 5032 45083
rect 4956 44959 5032 45027
rect 4956 44903 4966 44959
rect 5022 44903 5032 44959
rect 4956 44835 5032 44903
rect 4956 44779 4966 44835
rect 5022 44779 5032 44835
rect 4956 44711 5032 44779
rect 4956 44655 4966 44711
rect 5022 44655 5032 44711
rect 4956 44587 5032 44655
rect 4956 44531 4966 44587
rect 5022 44531 5032 44587
rect 4956 44463 5032 44531
rect 4956 44407 4966 44463
rect 5022 44407 5032 44463
rect 4956 44339 5032 44407
rect 4956 44283 4966 44339
rect 5022 44283 5032 44339
rect 1962 44207 1972 44263
rect 2028 44207 2038 44263
rect 1962 44139 2038 44207
rect 4956 44215 5032 44283
rect 4956 44159 4966 44215
rect 5022 44159 5032 44215
rect 4956 44149 5032 44159
rect 5080 45703 5156 45713
rect 5080 45647 5090 45703
rect 5146 45647 5156 45703
rect 5080 45579 5156 45647
rect 6384 45678 6460 45746
rect 6384 45622 6394 45678
rect 6450 45622 6460 45678
rect 5080 45523 5090 45579
rect 5146 45523 5156 45579
rect 5080 45455 5156 45523
rect 5080 45399 5090 45455
rect 5146 45399 5156 45455
rect 5080 45331 5156 45399
rect 5080 45275 5090 45331
rect 5146 45275 5156 45331
rect 5080 45207 5156 45275
rect 5080 45151 5090 45207
rect 5146 45151 5156 45207
rect 5080 45083 5156 45151
rect 5080 45027 5090 45083
rect 5146 45027 5156 45083
rect 5080 44959 5156 45027
rect 5080 44903 5090 44959
rect 5146 44903 5156 44959
rect 5080 44835 5156 44903
rect 5080 44779 5090 44835
rect 5146 44779 5156 44835
rect 5080 44711 5156 44779
rect 5080 44655 5090 44711
rect 5146 44655 5156 44711
rect 5080 44587 5156 44655
rect 5080 44531 5090 44587
rect 5146 44531 5156 44587
rect 5080 44463 5156 44531
rect 5080 44407 5090 44463
rect 5146 44407 5156 44463
rect 5080 44339 5156 44407
rect 5080 44283 5090 44339
rect 5146 44283 5156 44339
rect 5080 44215 5156 44283
rect 5080 44159 5090 44215
rect 5146 44159 5156 44215
rect 1962 44083 1972 44139
rect 2028 44083 2038 44139
rect 1962 44015 2038 44083
rect 5080 44091 5156 44159
rect 5080 44035 5090 44091
rect 5146 44035 5156 44091
rect 1962 43959 1972 44015
rect 2028 43959 2038 44015
rect 1962 43891 2038 43959
rect 1962 43835 1972 43891
rect 2028 43835 2038 43891
rect 1962 43767 2038 43835
rect 1962 43711 1972 43767
rect 2028 43711 2038 43767
rect 1962 43643 2038 43711
rect 1962 43587 1972 43643
rect 2028 43587 2038 43643
rect 1962 43519 2038 43587
rect 1962 43463 1972 43519
rect 2028 43463 2038 43519
rect 1962 43395 2038 43463
rect 1962 43339 1972 43395
rect 2028 43339 2038 43395
rect 1962 43271 2038 43339
rect 1962 43215 1972 43271
rect 2028 43215 2038 43271
rect 1962 43147 2038 43215
rect 1962 43091 1972 43147
rect 2028 43091 2038 43147
rect 1962 43023 2038 43091
rect 1962 42967 1972 43023
rect 2028 42967 2038 43023
rect 1962 42899 2038 42967
rect 1962 42843 1972 42899
rect 2028 42843 2038 42899
rect 1962 42775 2038 42843
rect 1962 42719 1972 42775
rect 2028 42719 2038 42775
rect 1962 42651 2038 42719
rect 1962 42595 1972 42651
rect 2028 42595 2038 42651
rect 1962 42585 2038 42595
rect 4460 44024 4536 44034
rect 5080 44025 5156 44035
rect 5204 45579 5280 45589
rect 5204 45523 5214 45579
rect 5270 45523 5280 45579
rect 5204 45455 5280 45523
rect 6384 45554 6460 45622
rect 6384 45498 6394 45554
rect 6450 45498 6460 45554
rect 5204 45399 5214 45455
rect 5270 45399 5280 45455
rect 5204 45331 5280 45399
rect 5204 45275 5214 45331
rect 5270 45275 5280 45331
rect 5204 45207 5280 45275
rect 5204 45151 5214 45207
rect 5270 45151 5280 45207
rect 5204 45083 5280 45151
rect 5204 45027 5214 45083
rect 5270 45027 5280 45083
rect 5204 44959 5280 45027
rect 5204 44903 5214 44959
rect 5270 44903 5280 44959
rect 5204 44835 5280 44903
rect 5204 44779 5214 44835
rect 5270 44779 5280 44835
rect 5204 44711 5280 44779
rect 5204 44655 5214 44711
rect 5270 44655 5280 44711
rect 5204 44587 5280 44655
rect 5204 44531 5214 44587
rect 5270 44531 5280 44587
rect 5204 44463 5280 44531
rect 5204 44407 5214 44463
rect 5270 44407 5280 44463
rect 5204 44339 5280 44407
rect 5204 44283 5214 44339
rect 5270 44283 5280 44339
rect 5204 44215 5280 44283
rect 5204 44159 5214 44215
rect 5270 44159 5280 44215
rect 5204 44091 5280 44159
rect 5204 44035 5214 44091
rect 5270 44035 5280 44091
rect 4460 43968 4470 44024
rect 4526 43968 4536 44024
rect 4460 43900 4536 43968
rect 5204 43967 5280 44035
rect 5204 43911 5214 43967
rect 5270 43911 5280 43967
rect 4460 43844 4470 43900
rect 4526 43844 4536 43900
rect 4460 43776 4536 43844
rect 4460 43720 4470 43776
rect 4526 43720 4536 43776
rect 4460 43652 4536 43720
rect 4460 43596 4470 43652
rect 4526 43596 4536 43652
rect 4460 43528 4536 43596
rect 4460 43472 4470 43528
rect 4526 43472 4536 43528
rect 4460 43404 4536 43472
rect 4460 43348 4470 43404
rect 4526 43348 4536 43404
rect 4460 43280 4536 43348
rect 4460 43224 4470 43280
rect 4526 43224 4536 43280
rect 4460 43156 4536 43224
rect 4460 43100 4470 43156
rect 4526 43100 4536 43156
rect 4460 43032 4536 43100
rect 4460 42976 4470 43032
rect 4526 42976 4536 43032
rect 4460 42908 4536 42976
rect 4460 42852 4470 42908
rect 4526 42852 4536 42908
rect 4460 42784 4536 42852
rect 4460 42728 4470 42784
rect 4526 42728 4536 42784
rect 4460 42660 4536 42728
rect 4460 42604 4470 42660
rect 4526 42604 4536 42660
rect 4460 42536 4536 42604
rect 4460 42480 4470 42536
rect 4526 42480 4536 42536
rect 4460 42412 4536 42480
rect 4460 42356 4470 42412
rect 4526 42356 4536 42412
rect 4460 42346 4536 42356
rect 4584 43900 4660 43910
rect 5204 43901 5280 43911
rect 5328 45455 5404 45465
rect 5328 45399 5338 45455
rect 5394 45399 5404 45455
rect 5328 45331 5404 45399
rect 6384 45430 6460 45498
rect 6384 45374 6394 45430
rect 6450 45374 6460 45430
rect 5328 45275 5338 45331
rect 5394 45275 5404 45331
rect 5328 45207 5404 45275
rect 5328 45151 5338 45207
rect 5394 45151 5404 45207
rect 5328 45083 5404 45151
rect 5328 45027 5338 45083
rect 5394 45027 5404 45083
rect 5328 44959 5404 45027
rect 5328 44903 5338 44959
rect 5394 44903 5404 44959
rect 5328 44835 5404 44903
rect 5328 44779 5338 44835
rect 5394 44779 5404 44835
rect 5328 44711 5404 44779
rect 5328 44655 5338 44711
rect 5394 44655 5404 44711
rect 5328 44587 5404 44655
rect 5328 44531 5338 44587
rect 5394 44531 5404 44587
rect 5328 44463 5404 44531
rect 5328 44407 5338 44463
rect 5394 44407 5404 44463
rect 5328 44339 5404 44407
rect 5328 44283 5338 44339
rect 5394 44283 5404 44339
rect 5328 44215 5404 44283
rect 5328 44159 5338 44215
rect 5394 44159 5404 44215
rect 5328 44091 5404 44159
rect 5328 44035 5338 44091
rect 5394 44035 5404 44091
rect 5328 43967 5404 44035
rect 5328 43911 5338 43967
rect 5394 43911 5404 43967
rect 4584 43844 4594 43900
rect 4650 43844 4660 43900
rect 4584 43776 4660 43844
rect 5328 43843 5404 43911
rect 5328 43787 5338 43843
rect 5394 43787 5404 43843
rect 4584 43720 4594 43776
rect 4650 43720 4660 43776
rect 4584 43652 4660 43720
rect 4584 43596 4594 43652
rect 4650 43596 4660 43652
rect 4584 43528 4660 43596
rect 4584 43472 4594 43528
rect 4650 43472 4660 43528
rect 4584 43404 4660 43472
rect 4584 43348 4594 43404
rect 4650 43348 4660 43404
rect 4584 43280 4660 43348
rect 4584 43224 4594 43280
rect 4650 43224 4660 43280
rect 4584 43156 4660 43224
rect 4584 43100 4594 43156
rect 4650 43100 4660 43156
rect 4584 43032 4660 43100
rect 4584 42976 4594 43032
rect 4650 42976 4660 43032
rect 4584 42908 4660 42976
rect 4584 42852 4594 42908
rect 4650 42852 4660 42908
rect 4584 42784 4660 42852
rect 4584 42728 4594 42784
rect 4650 42728 4660 42784
rect 4584 42660 4660 42728
rect 4584 42604 4594 42660
rect 4650 42604 4660 42660
rect 4584 42536 4660 42604
rect 4584 42480 4594 42536
rect 4650 42480 4660 42536
rect 4584 42412 4660 42480
rect 4584 42356 4594 42412
rect 4650 42356 4660 42412
rect 4584 42288 4660 42356
rect 4584 42232 4594 42288
rect 4650 42232 4660 42288
rect 4584 42222 4660 42232
rect 4708 43776 4784 43786
rect 5328 43777 5404 43787
rect 5452 45331 5528 45341
rect 5452 45275 5462 45331
rect 5518 45275 5528 45331
rect 5452 45207 5528 45275
rect 6384 45306 6460 45374
rect 6384 45250 6394 45306
rect 6450 45250 6460 45306
rect 5452 45151 5462 45207
rect 5518 45151 5528 45207
rect 5452 45083 5528 45151
rect 5452 45027 5462 45083
rect 5518 45027 5528 45083
rect 5452 44959 5528 45027
rect 5452 44903 5462 44959
rect 5518 44903 5528 44959
rect 5452 44835 5528 44903
rect 5452 44779 5462 44835
rect 5518 44779 5528 44835
rect 5452 44711 5528 44779
rect 5452 44655 5462 44711
rect 5518 44655 5528 44711
rect 5452 44587 5528 44655
rect 5452 44531 5462 44587
rect 5518 44531 5528 44587
rect 5452 44463 5528 44531
rect 5452 44407 5462 44463
rect 5518 44407 5528 44463
rect 5452 44339 5528 44407
rect 5452 44283 5462 44339
rect 5518 44283 5528 44339
rect 5452 44215 5528 44283
rect 5452 44159 5462 44215
rect 5518 44159 5528 44215
rect 5452 44091 5528 44159
rect 5452 44035 5462 44091
rect 5518 44035 5528 44091
rect 5452 43967 5528 44035
rect 5452 43911 5462 43967
rect 5518 43911 5528 43967
rect 5452 43843 5528 43911
rect 5452 43787 5462 43843
rect 5518 43787 5528 43843
rect 4708 43720 4718 43776
rect 4774 43720 4784 43776
rect 4708 43652 4784 43720
rect 5452 43719 5528 43787
rect 5452 43663 5462 43719
rect 5518 43663 5528 43719
rect 4708 43596 4718 43652
rect 4774 43596 4784 43652
rect 4708 43528 4784 43596
rect 4708 43472 4718 43528
rect 4774 43472 4784 43528
rect 4708 43404 4784 43472
rect 4708 43348 4718 43404
rect 4774 43348 4784 43404
rect 4708 43280 4784 43348
rect 4708 43224 4718 43280
rect 4774 43224 4784 43280
rect 4708 43156 4784 43224
rect 4708 43100 4718 43156
rect 4774 43100 4784 43156
rect 4708 43032 4784 43100
rect 4708 42976 4718 43032
rect 4774 42976 4784 43032
rect 4708 42908 4784 42976
rect 4708 42852 4718 42908
rect 4774 42852 4784 42908
rect 4708 42784 4784 42852
rect 4708 42728 4718 42784
rect 4774 42728 4784 42784
rect 4708 42660 4784 42728
rect 4708 42604 4718 42660
rect 4774 42604 4784 42660
rect 4708 42536 4784 42604
rect 4708 42480 4718 42536
rect 4774 42480 4784 42536
rect 4708 42412 4784 42480
rect 4708 42356 4718 42412
rect 4774 42356 4784 42412
rect 4708 42288 4784 42356
rect 4708 42232 4718 42288
rect 4774 42232 4784 42288
rect 4708 42164 4784 42232
rect 4708 42108 4718 42164
rect 4774 42108 4784 42164
rect 4708 42098 4784 42108
rect 4832 43652 4908 43662
rect 5452 43653 5528 43663
rect 5576 45207 5652 45217
rect 5576 45151 5586 45207
rect 5642 45151 5652 45207
rect 5576 45083 5652 45151
rect 6384 45182 6460 45250
rect 6384 45126 6394 45182
rect 6450 45126 6460 45182
rect 5576 45027 5586 45083
rect 5642 45027 5652 45083
rect 5576 44959 5652 45027
rect 5576 44903 5586 44959
rect 5642 44903 5652 44959
rect 5576 44835 5652 44903
rect 5576 44779 5586 44835
rect 5642 44779 5652 44835
rect 5576 44711 5652 44779
rect 5576 44655 5586 44711
rect 5642 44655 5652 44711
rect 5576 44587 5652 44655
rect 5576 44531 5586 44587
rect 5642 44531 5652 44587
rect 5576 44463 5652 44531
rect 5576 44407 5586 44463
rect 5642 44407 5652 44463
rect 5576 44339 5652 44407
rect 5576 44283 5586 44339
rect 5642 44283 5652 44339
rect 5576 44215 5652 44283
rect 5576 44159 5586 44215
rect 5642 44159 5652 44215
rect 5576 44091 5652 44159
rect 5576 44035 5586 44091
rect 5642 44035 5652 44091
rect 5576 43967 5652 44035
rect 5576 43911 5586 43967
rect 5642 43911 5652 43967
rect 5576 43843 5652 43911
rect 5576 43787 5586 43843
rect 5642 43787 5652 43843
rect 5576 43719 5652 43787
rect 5576 43663 5586 43719
rect 5642 43663 5652 43719
rect 4832 43596 4842 43652
rect 4898 43596 4908 43652
rect 4832 43528 4908 43596
rect 5576 43595 5652 43663
rect 5576 43539 5586 43595
rect 5642 43539 5652 43595
rect 4832 43472 4842 43528
rect 4898 43472 4908 43528
rect 4832 43404 4908 43472
rect 4832 43348 4842 43404
rect 4898 43348 4908 43404
rect 4832 43280 4908 43348
rect 4832 43224 4842 43280
rect 4898 43224 4908 43280
rect 4832 43156 4908 43224
rect 4832 43100 4842 43156
rect 4898 43100 4908 43156
rect 4832 43032 4908 43100
rect 4832 42976 4842 43032
rect 4898 42976 4908 43032
rect 4832 42908 4908 42976
rect 4832 42852 4842 42908
rect 4898 42852 4908 42908
rect 4832 42784 4908 42852
rect 4832 42728 4842 42784
rect 4898 42728 4908 42784
rect 4832 42660 4908 42728
rect 4832 42604 4842 42660
rect 4898 42604 4908 42660
rect 4832 42536 4908 42604
rect 4832 42480 4842 42536
rect 4898 42480 4908 42536
rect 4832 42412 4908 42480
rect 4832 42356 4842 42412
rect 4898 42356 4908 42412
rect 4832 42288 4908 42356
rect 4832 42232 4842 42288
rect 4898 42232 4908 42288
rect 4832 42164 4908 42232
rect 4832 42108 4842 42164
rect 4898 42108 4908 42164
rect 4832 42040 4908 42108
rect 4832 41984 4842 42040
rect 4898 41984 4908 42040
rect 4832 41974 4908 41984
rect 4956 43528 5032 43538
rect 5576 43529 5652 43539
rect 5700 45083 5776 45093
rect 5700 45027 5710 45083
rect 5766 45027 5776 45083
rect 5700 44959 5776 45027
rect 6384 45058 6460 45126
rect 6384 45002 6394 45058
rect 6450 45002 6460 45058
rect 6384 44992 6460 45002
rect 6508 46546 6584 46556
rect 6508 46490 6518 46546
rect 6574 46490 6584 46546
rect 6508 46422 6584 46490
rect 6508 46366 6518 46422
rect 6574 46366 6584 46422
rect 6508 46298 6584 46366
rect 6508 46242 6518 46298
rect 6574 46242 6584 46298
rect 6508 46174 6584 46242
rect 6508 46118 6518 46174
rect 6574 46118 6584 46174
rect 6508 46050 6584 46118
rect 6508 45994 6518 46050
rect 6574 45994 6584 46050
rect 6508 45926 6584 45994
rect 6508 45870 6518 45926
rect 6574 45870 6584 45926
rect 6508 45802 6584 45870
rect 6508 45746 6518 45802
rect 6574 45746 6584 45802
rect 6508 45678 6584 45746
rect 6508 45622 6518 45678
rect 6574 45622 6584 45678
rect 6508 45554 6584 45622
rect 6508 45498 6518 45554
rect 6574 45498 6584 45554
rect 6508 45430 6584 45498
rect 6508 45374 6518 45430
rect 6574 45374 6584 45430
rect 6508 45306 6584 45374
rect 6508 45250 6518 45306
rect 6574 45250 6584 45306
rect 6508 45182 6584 45250
rect 6508 45126 6518 45182
rect 6574 45126 6584 45182
rect 6508 45058 6584 45126
rect 6508 45002 6518 45058
rect 6574 45002 6584 45058
rect 5700 44903 5710 44959
rect 5766 44903 5776 44959
rect 5700 44835 5776 44903
rect 5700 44779 5710 44835
rect 5766 44779 5776 44835
rect 5700 44711 5776 44779
rect 5700 44655 5710 44711
rect 5766 44655 5776 44711
rect 5700 44587 5776 44655
rect 5700 44531 5710 44587
rect 5766 44531 5776 44587
rect 5700 44463 5776 44531
rect 5700 44407 5710 44463
rect 5766 44407 5776 44463
rect 5700 44339 5776 44407
rect 5700 44283 5710 44339
rect 5766 44283 5776 44339
rect 5700 44215 5776 44283
rect 5700 44159 5710 44215
rect 5766 44159 5776 44215
rect 5700 44091 5776 44159
rect 5700 44035 5710 44091
rect 5766 44035 5776 44091
rect 5700 43967 5776 44035
rect 5700 43911 5710 43967
rect 5766 43911 5776 43967
rect 5700 43843 5776 43911
rect 5700 43787 5710 43843
rect 5766 43787 5776 43843
rect 5700 43719 5776 43787
rect 5700 43663 5710 43719
rect 5766 43663 5776 43719
rect 5700 43595 5776 43663
rect 5700 43539 5710 43595
rect 5766 43539 5776 43595
rect 4956 43472 4966 43528
rect 5022 43472 5032 43528
rect 4956 43404 5032 43472
rect 5700 43471 5776 43539
rect 5700 43415 5710 43471
rect 5766 43415 5776 43471
rect 4956 43348 4966 43404
rect 5022 43348 5032 43404
rect 4956 43280 5032 43348
rect 4956 43224 4966 43280
rect 5022 43224 5032 43280
rect 4956 43156 5032 43224
rect 4956 43100 4966 43156
rect 5022 43100 5032 43156
rect 4956 43032 5032 43100
rect 4956 42976 4966 43032
rect 5022 42976 5032 43032
rect 4956 42908 5032 42976
rect 4956 42852 4966 42908
rect 5022 42852 5032 42908
rect 4956 42784 5032 42852
rect 4956 42728 4966 42784
rect 5022 42728 5032 42784
rect 4956 42660 5032 42728
rect 4956 42604 4966 42660
rect 5022 42604 5032 42660
rect 4956 42536 5032 42604
rect 4956 42480 4966 42536
rect 5022 42480 5032 42536
rect 4956 42412 5032 42480
rect 4956 42356 4966 42412
rect 5022 42356 5032 42412
rect 4956 42288 5032 42356
rect 4956 42232 4966 42288
rect 5022 42232 5032 42288
rect 4956 42164 5032 42232
rect 4956 42108 4966 42164
rect 5022 42108 5032 42164
rect 4956 42040 5032 42108
rect 4956 41984 4966 42040
rect 5022 41984 5032 42040
rect 4956 41916 5032 41984
rect 4956 41860 4966 41916
rect 5022 41860 5032 41916
rect 4956 41850 5032 41860
rect 5080 43404 5156 43414
rect 5700 43405 5776 43415
rect 5824 44959 5900 44969
rect 5824 44903 5834 44959
rect 5890 44903 5900 44959
rect 5824 44835 5900 44903
rect 6508 44934 6584 45002
rect 6508 44878 6518 44934
rect 6574 44878 6584 44934
rect 6508 44868 6584 44878
rect 6632 46422 6708 46432
rect 6632 46366 6642 46422
rect 6698 46366 6708 46422
rect 6632 46298 6708 46366
rect 6632 46242 6642 46298
rect 6698 46242 6708 46298
rect 6632 46174 6708 46242
rect 6632 46118 6642 46174
rect 6698 46118 6708 46174
rect 6632 46050 6708 46118
rect 6632 45994 6642 46050
rect 6698 45994 6708 46050
rect 6632 45926 6708 45994
rect 6632 45870 6642 45926
rect 6698 45870 6708 45926
rect 6632 45802 6708 45870
rect 6632 45746 6642 45802
rect 6698 45746 6708 45802
rect 6632 45678 6708 45746
rect 6632 45622 6642 45678
rect 6698 45622 6708 45678
rect 6632 45554 6708 45622
rect 6632 45498 6642 45554
rect 6698 45498 6708 45554
rect 6632 45430 6708 45498
rect 6632 45374 6642 45430
rect 6698 45374 6708 45430
rect 6632 45306 6708 45374
rect 6632 45250 6642 45306
rect 6698 45250 6708 45306
rect 6632 45182 6708 45250
rect 6632 45126 6642 45182
rect 6698 45126 6708 45182
rect 6632 45058 6708 45126
rect 6632 45002 6642 45058
rect 6698 45002 6708 45058
rect 6632 44934 6708 45002
rect 6632 44878 6642 44934
rect 6698 44878 6708 44934
rect 5824 44779 5834 44835
rect 5890 44779 5900 44835
rect 5824 44711 5900 44779
rect 5824 44655 5834 44711
rect 5890 44655 5900 44711
rect 5824 44587 5900 44655
rect 5824 44531 5834 44587
rect 5890 44531 5900 44587
rect 5824 44463 5900 44531
rect 5824 44407 5834 44463
rect 5890 44407 5900 44463
rect 5824 44339 5900 44407
rect 5824 44283 5834 44339
rect 5890 44283 5900 44339
rect 5824 44215 5900 44283
rect 5824 44159 5834 44215
rect 5890 44159 5900 44215
rect 5824 44091 5900 44159
rect 5824 44035 5834 44091
rect 5890 44035 5900 44091
rect 5824 43967 5900 44035
rect 5824 43911 5834 43967
rect 5890 43911 5900 43967
rect 5824 43843 5900 43911
rect 5824 43787 5834 43843
rect 5890 43787 5900 43843
rect 5824 43719 5900 43787
rect 5824 43663 5834 43719
rect 5890 43663 5900 43719
rect 5824 43595 5900 43663
rect 5824 43539 5834 43595
rect 5890 43539 5900 43595
rect 5824 43471 5900 43539
rect 5824 43415 5834 43471
rect 5890 43415 5900 43471
rect 5080 43348 5090 43404
rect 5146 43348 5156 43404
rect 5080 43280 5156 43348
rect 5824 43347 5900 43415
rect 5824 43291 5834 43347
rect 5890 43291 5900 43347
rect 5080 43224 5090 43280
rect 5146 43224 5156 43280
rect 5080 43156 5156 43224
rect 5080 43100 5090 43156
rect 5146 43100 5156 43156
rect 5080 43032 5156 43100
rect 5080 42976 5090 43032
rect 5146 42976 5156 43032
rect 5080 42908 5156 42976
rect 5080 42852 5090 42908
rect 5146 42852 5156 42908
rect 5080 42784 5156 42852
rect 5080 42728 5090 42784
rect 5146 42728 5156 42784
rect 5080 42660 5156 42728
rect 5080 42604 5090 42660
rect 5146 42604 5156 42660
rect 5080 42536 5156 42604
rect 5080 42480 5090 42536
rect 5146 42480 5156 42536
rect 5080 42412 5156 42480
rect 5080 42356 5090 42412
rect 5146 42356 5156 42412
rect 5080 42288 5156 42356
rect 5080 42232 5090 42288
rect 5146 42232 5156 42288
rect 5080 42164 5156 42232
rect 5080 42108 5090 42164
rect 5146 42108 5156 42164
rect 5080 42040 5156 42108
rect 5080 41984 5090 42040
rect 5146 41984 5156 42040
rect 5080 41916 5156 41984
rect 5080 41860 5090 41916
rect 5146 41860 5156 41916
rect 4460 41789 4536 41799
rect 4460 41733 4470 41789
rect 4526 41733 4536 41789
rect 4460 41665 4536 41733
rect 5080 41792 5156 41860
rect 5080 41736 5090 41792
rect 5146 41736 5156 41792
rect 5080 41726 5156 41736
rect 5204 43280 5280 43290
rect 5824 43281 5900 43291
rect 5948 44835 6024 44845
rect 5948 44779 5958 44835
rect 6014 44779 6024 44835
rect 5948 44711 6024 44779
rect 6632 44810 6708 44878
rect 6632 44754 6642 44810
rect 6698 44754 6708 44810
rect 6632 44744 6708 44754
rect 6756 46298 6832 46308
rect 6756 46242 6766 46298
rect 6822 46242 6832 46298
rect 6756 46174 6832 46242
rect 6756 46118 6766 46174
rect 6822 46118 6832 46174
rect 6756 46050 6832 46118
rect 6756 45994 6766 46050
rect 6822 45994 6832 46050
rect 6756 45926 6832 45994
rect 6756 45870 6766 45926
rect 6822 45870 6832 45926
rect 6756 45802 6832 45870
rect 6756 45746 6766 45802
rect 6822 45746 6832 45802
rect 6756 45678 6832 45746
rect 6756 45622 6766 45678
rect 6822 45622 6832 45678
rect 6756 45554 6832 45622
rect 6756 45498 6766 45554
rect 6822 45498 6832 45554
rect 6756 45430 6832 45498
rect 6756 45374 6766 45430
rect 6822 45374 6832 45430
rect 6756 45306 6832 45374
rect 6756 45250 6766 45306
rect 6822 45250 6832 45306
rect 6756 45182 6832 45250
rect 6756 45126 6766 45182
rect 6822 45126 6832 45182
rect 6756 45058 6832 45126
rect 6756 45002 6766 45058
rect 6822 45002 6832 45058
rect 6756 44934 6832 45002
rect 6756 44878 6766 44934
rect 6822 44878 6832 44934
rect 6756 44810 6832 44878
rect 6756 44754 6766 44810
rect 6822 44754 6832 44810
rect 5948 44655 5958 44711
rect 6014 44655 6024 44711
rect 5948 44587 6024 44655
rect 5948 44531 5958 44587
rect 6014 44531 6024 44587
rect 5948 44463 6024 44531
rect 5948 44407 5958 44463
rect 6014 44407 6024 44463
rect 5948 44339 6024 44407
rect 5948 44283 5958 44339
rect 6014 44283 6024 44339
rect 5948 44215 6024 44283
rect 5948 44159 5958 44215
rect 6014 44159 6024 44215
rect 5948 44091 6024 44159
rect 5948 44035 5958 44091
rect 6014 44035 6024 44091
rect 5948 43967 6024 44035
rect 5948 43911 5958 43967
rect 6014 43911 6024 43967
rect 5948 43843 6024 43911
rect 5948 43787 5958 43843
rect 6014 43787 6024 43843
rect 5948 43719 6024 43787
rect 5948 43663 5958 43719
rect 6014 43663 6024 43719
rect 5948 43595 6024 43663
rect 5948 43539 5958 43595
rect 6014 43539 6024 43595
rect 5948 43471 6024 43539
rect 5948 43415 5958 43471
rect 6014 43415 6024 43471
rect 5948 43347 6024 43415
rect 5948 43291 5958 43347
rect 6014 43291 6024 43347
rect 5204 43224 5214 43280
rect 5270 43224 5280 43280
rect 5204 43156 5280 43224
rect 5948 43223 6024 43291
rect 5948 43167 5958 43223
rect 6014 43167 6024 43223
rect 5204 43100 5214 43156
rect 5270 43100 5280 43156
rect 5204 43032 5280 43100
rect 5204 42976 5214 43032
rect 5270 42976 5280 43032
rect 5204 42908 5280 42976
rect 5204 42852 5214 42908
rect 5270 42852 5280 42908
rect 5204 42784 5280 42852
rect 5204 42728 5214 42784
rect 5270 42728 5280 42784
rect 5204 42660 5280 42728
rect 5204 42604 5214 42660
rect 5270 42604 5280 42660
rect 5204 42536 5280 42604
rect 5204 42480 5214 42536
rect 5270 42480 5280 42536
rect 5204 42412 5280 42480
rect 5204 42356 5214 42412
rect 5270 42356 5280 42412
rect 5204 42288 5280 42356
rect 5204 42232 5214 42288
rect 5270 42232 5280 42288
rect 5204 42164 5280 42232
rect 5204 42108 5214 42164
rect 5270 42108 5280 42164
rect 5204 42040 5280 42108
rect 5204 41984 5214 42040
rect 5270 41984 5280 42040
rect 5204 41916 5280 41984
rect 5204 41860 5214 41916
rect 5270 41860 5280 41916
rect 5204 41792 5280 41860
rect 5204 41736 5214 41792
rect 5270 41736 5280 41792
rect 4460 41609 4470 41665
rect 4526 41609 4536 41665
rect 4460 41541 4536 41609
rect 4460 41485 4470 41541
rect 4526 41485 4536 41541
rect 4460 41417 4536 41485
rect 4460 41361 4470 41417
rect 4526 41361 4536 41417
rect 4460 41293 4536 41361
rect 4460 41237 4470 41293
rect 4526 41237 4536 41293
rect 4460 41169 4536 41237
rect 4460 41113 4470 41169
rect 4526 41113 4536 41169
rect 4460 41045 4536 41113
rect 4460 40989 4470 41045
rect 4526 40989 4536 41045
rect 4460 40921 4536 40989
rect 4460 40865 4470 40921
rect 4526 40865 4536 40921
rect 4460 40797 4536 40865
rect 4460 40741 4470 40797
rect 4526 40741 4536 40797
rect 4460 40673 4536 40741
rect 4460 40617 4470 40673
rect 4526 40617 4536 40673
rect 4460 40549 4536 40617
rect 4460 40493 4470 40549
rect 4526 40493 4536 40549
rect 4460 40425 4536 40493
rect 4460 40369 4470 40425
rect 4526 40369 4536 40425
rect 4460 40301 4536 40369
rect 4460 40245 4470 40301
rect 4526 40245 4536 40301
rect 4460 40177 4536 40245
rect 4460 40121 4470 40177
rect 4526 40121 4536 40177
rect 4460 40111 4536 40121
rect 4584 41665 4660 41675
rect 4584 41609 4594 41665
rect 4650 41609 4660 41665
rect 4584 41541 4660 41609
rect 5204 41668 5280 41736
rect 5204 41612 5214 41668
rect 5270 41612 5280 41668
rect 5204 41602 5280 41612
rect 5328 43156 5404 43166
rect 5948 43157 6024 43167
rect 6072 44711 6148 44721
rect 6072 44655 6082 44711
rect 6138 44655 6148 44711
rect 6072 44587 6148 44655
rect 6756 44686 6832 44754
rect 6756 44630 6766 44686
rect 6822 44630 6832 44686
rect 6756 44620 6832 44630
rect 6880 46174 6956 46184
rect 6880 46118 6890 46174
rect 6946 46118 6956 46174
rect 6880 46050 6956 46118
rect 6880 45994 6890 46050
rect 6946 45994 6956 46050
rect 6880 45926 6956 45994
rect 6880 45870 6890 45926
rect 6946 45870 6956 45926
rect 6880 45802 6956 45870
rect 6880 45746 6890 45802
rect 6946 45746 6956 45802
rect 6880 45678 6956 45746
rect 6880 45622 6890 45678
rect 6946 45622 6956 45678
rect 6880 45554 6956 45622
rect 6880 45498 6890 45554
rect 6946 45498 6956 45554
rect 6880 45430 6956 45498
rect 6880 45374 6890 45430
rect 6946 45374 6956 45430
rect 6880 45306 6956 45374
rect 6880 45250 6890 45306
rect 6946 45250 6956 45306
rect 6880 45182 6956 45250
rect 6880 45126 6890 45182
rect 6946 45126 6956 45182
rect 6880 45058 6956 45126
rect 6880 45002 6890 45058
rect 6946 45002 6956 45058
rect 6880 44934 6956 45002
rect 6880 44878 6890 44934
rect 6946 44878 6956 44934
rect 6880 44810 6956 44878
rect 6880 44754 6890 44810
rect 6946 44754 6956 44810
rect 6880 44686 6956 44754
rect 6880 44630 6890 44686
rect 6946 44630 6956 44686
rect 6072 44531 6082 44587
rect 6138 44531 6148 44587
rect 6072 44463 6148 44531
rect 6880 44562 6956 44630
rect 6880 44506 6890 44562
rect 6946 44506 6956 44562
rect 6880 44496 6956 44506
rect 7004 46050 7080 46060
rect 7004 45994 7014 46050
rect 7070 45994 7080 46050
rect 7004 45926 7080 45994
rect 7004 45870 7014 45926
rect 7070 45870 7080 45926
rect 7004 45802 7080 45870
rect 7004 45746 7014 45802
rect 7070 45746 7080 45802
rect 7004 45678 7080 45746
rect 7004 45622 7014 45678
rect 7070 45622 7080 45678
rect 7004 45554 7080 45622
rect 7004 45498 7014 45554
rect 7070 45498 7080 45554
rect 7004 45430 7080 45498
rect 7004 45374 7014 45430
rect 7070 45374 7080 45430
rect 7004 45306 7080 45374
rect 7004 45250 7014 45306
rect 7070 45250 7080 45306
rect 7004 45182 7080 45250
rect 7004 45126 7014 45182
rect 7070 45126 7080 45182
rect 7004 45058 7080 45126
rect 7004 45002 7014 45058
rect 7070 45002 7080 45058
rect 7004 44934 7080 45002
rect 7004 44878 7014 44934
rect 7070 44878 7080 44934
rect 7004 44810 7080 44878
rect 7004 44754 7014 44810
rect 7070 44754 7080 44810
rect 7004 44686 7080 44754
rect 7004 44630 7014 44686
rect 7070 44630 7080 44686
rect 7004 44562 7080 44630
rect 7004 44506 7014 44562
rect 7070 44506 7080 44562
rect 6072 44407 6082 44463
rect 6138 44407 6148 44463
rect 6072 44339 6148 44407
rect 7004 44438 7080 44506
rect 7004 44382 7014 44438
rect 7070 44382 7080 44438
rect 7004 44372 7080 44382
rect 7128 45926 7204 45936
rect 7128 45870 7138 45926
rect 7194 45870 7204 45926
rect 7128 45802 7204 45870
rect 7128 45746 7138 45802
rect 7194 45746 7204 45802
rect 7128 45678 7204 45746
rect 7128 45622 7138 45678
rect 7194 45622 7204 45678
rect 7128 45554 7204 45622
rect 7128 45498 7138 45554
rect 7194 45498 7204 45554
rect 7128 45430 7204 45498
rect 7128 45374 7138 45430
rect 7194 45374 7204 45430
rect 7128 45306 7204 45374
rect 7128 45250 7138 45306
rect 7194 45250 7204 45306
rect 7128 45182 7204 45250
rect 7128 45126 7138 45182
rect 7194 45126 7204 45182
rect 7128 45058 7204 45126
rect 7128 45002 7138 45058
rect 7194 45002 7204 45058
rect 7128 44934 7204 45002
rect 7128 44878 7138 44934
rect 7194 44878 7204 44934
rect 7128 44810 7204 44878
rect 7128 44754 7138 44810
rect 7194 44754 7204 44810
rect 7128 44686 7204 44754
rect 7128 44630 7138 44686
rect 7194 44630 7204 44686
rect 7128 44562 7204 44630
rect 7128 44506 7138 44562
rect 7194 44506 7204 44562
rect 7128 44438 7204 44506
rect 7128 44382 7138 44438
rect 7194 44382 7204 44438
rect 6072 44283 6082 44339
rect 6138 44283 6148 44339
rect 6072 44215 6148 44283
rect 7128 44314 7204 44382
rect 7128 44258 7138 44314
rect 7194 44258 7204 44314
rect 7128 44248 7204 44258
rect 7252 45802 7328 45812
rect 7252 45746 7262 45802
rect 7318 45746 7328 45802
rect 7252 45678 7328 45746
rect 7252 45622 7262 45678
rect 7318 45622 7328 45678
rect 7252 45554 7328 45622
rect 7252 45498 7262 45554
rect 7318 45498 7328 45554
rect 7252 45430 7328 45498
rect 7252 45374 7262 45430
rect 7318 45374 7328 45430
rect 7252 45306 7328 45374
rect 7252 45250 7262 45306
rect 7318 45250 7328 45306
rect 7252 45182 7328 45250
rect 7252 45126 7262 45182
rect 7318 45126 7328 45182
rect 7252 45058 7328 45126
rect 7252 45002 7262 45058
rect 7318 45002 7328 45058
rect 7252 44934 7328 45002
rect 7252 44878 7262 44934
rect 7318 44878 7328 44934
rect 7252 44810 7328 44878
rect 7252 44754 7262 44810
rect 7318 44754 7328 44810
rect 7252 44686 7328 44754
rect 7252 44630 7262 44686
rect 7318 44630 7328 44686
rect 7252 44562 7328 44630
rect 7252 44506 7262 44562
rect 7318 44506 7328 44562
rect 7252 44438 7328 44506
rect 7252 44382 7262 44438
rect 7318 44382 7328 44438
rect 7252 44314 7328 44382
rect 7252 44258 7262 44314
rect 7318 44258 7328 44314
rect 6072 44159 6082 44215
rect 6138 44159 6148 44215
rect 6072 44091 6148 44159
rect 7252 44190 7328 44258
rect 7252 44134 7262 44190
rect 7318 44134 7328 44190
rect 7252 44124 7328 44134
rect 8741 44544 10553 44554
rect 8741 44488 8751 44544
rect 8807 44488 8875 44544
rect 8931 44488 8999 44544
rect 9055 44488 9123 44544
rect 9179 44488 9247 44544
rect 9303 44488 9371 44544
rect 9427 44488 9495 44544
rect 9551 44488 9619 44544
rect 9675 44488 9743 44544
rect 9799 44488 9867 44544
rect 9923 44488 9991 44544
rect 10047 44488 10115 44544
rect 10171 44488 10239 44544
rect 10295 44488 10363 44544
rect 10419 44488 10487 44544
rect 10543 44488 10553 44544
rect 8741 44420 10553 44488
rect 8741 44364 8751 44420
rect 8807 44364 8875 44420
rect 8931 44364 8999 44420
rect 9055 44364 9123 44420
rect 9179 44364 9247 44420
rect 9303 44364 9371 44420
rect 9427 44364 9495 44420
rect 9551 44364 9619 44420
rect 9675 44364 9743 44420
rect 9799 44364 9867 44420
rect 9923 44364 9991 44420
rect 10047 44364 10115 44420
rect 10171 44364 10239 44420
rect 10295 44364 10363 44420
rect 10419 44364 10487 44420
rect 10543 44364 10553 44420
rect 8741 44296 10553 44364
rect 8741 44240 8751 44296
rect 8807 44240 8875 44296
rect 8931 44240 8999 44296
rect 9055 44240 9123 44296
rect 9179 44240 9247 44296
rect 9303 44240 9371 44296
rect 9427 44240 9495 44296
rect 9551 44240 9619 44296
rect 9675 44240 9743 44296
rect 9799 44240 9867 44296
rect 9923 44240 9991 44296
rect 10047 44240 10115 44296
rect 10171 44240 10239 44296
rect 10295 44240 10363 44296
rect 10419 44240 10487 44296
rect 10543 44240 10553 44296
rect 8741 44172 10553 44240
rect 6072 44035 6082 44091
rect 6138 44035 6148 44091
rect 6072 43967 6148 44035
rect 6072 43911 6082 43967
rect 6138 43911 6148 43967
rect 6072 43843 6148 43911
rect 6072 43787 6082 43843
rect 6138 43787 6148 43843
rect 6072 43719 6148 43787
rect 6072 43663 6082 43719
rect 6138 43663 6148 43719
rect 6072 43595 6148 43663
rect 6072 43539 6082 43595
rect 6138 43539 6148 43595
rect 6072 43471 6148 43539
rect 6072 43415 6082 43471
rect 6138 43415 6148 43471
rect 6072 43347 6148 43415
rect 6072 43291 6082 43347
rect 6138 43291 6148 43347
rect 6072 43223 6148 43291
rect 8741 44116 8751 44172
rect 8807 44116 8875 44172
rect 8931 44116 8999 44172
rect 9055 44116 9123 44172
rect 9179 44116 9247 44172
rect 9303 44116 9371 44172
rect 9427 44116 9495 44172
rect 9551 44116 9619 44172
rect 9675 44116 9743 44172
rect 9799 44116 9867 44172
rect 9923 44116 9991 44172
rect 10047 44116 10115 44172
rect 10171 44116 10239 44172
rect 10295 44116 10363 44172
rect 10419 44116 10487 44172
rect 10543 44116 10553 44172
rect 8741 44048 10553 44116
rect 8741 43992 8751 44048
rect 8807 43992 8875 44048
rect 8931 43992 8999 44048
rect 9055 43992 9123 44048
rect 9179 43992 9247 44048
rect 9303 43992 9371 44048
rect 9427 43992 9495 44048
rect 9551 43992 9619 44048
rect 9675 43992 9743 44048
rect 9799 43992 9867 44048
rect 9923 43992 9991 44048
rect 10047 43992 10115 44048
rect 10171 43992 10239 44048
rect 10295 43992 10363 44048
rect 10419 43992 10487 44048
rect 10543 43992 10553 44048
rect 8741 43924 10553 43992
rect 8741 43868 8751 43924
rect 8807 43868 8875 43924
rect 8931 43868 8999 43924
rect 9055 43868 9123 43924
rect 9179 43868 9247 43924
rect 9303 43868 9371 43924
rect 9427 43868 9495 43924
rect 9551 43868 9619 43924
rect 9675 43868 9743 43924
rect 9799 43868 9867 43924
rect 9923 43868 9991 43924
rect 10047 43868 10115 43924
rect 10171 43868 10239 43924
rect 10295 43868 10363 43924
rect 10419 43868 10487 43924
rect 10543 43868 10553 43924
rect 8741 43800 10553 43868
rect 8741 43744 8751 43800
rect 8807 43744 8875 43800
rect 8931 43744 8999 43800
rect 9055 43744 9123 43800
rect 9179 43744 9247 43800
rect 9303 43744 9371 43800
rect 9427 43744 9495 43800
rect 9551 43744 9619 43800
rect 9675 43744 9743 43800
rect 9799 43744 9867 43800
rect 9923 43744 9991 43800
rect 10047 43744 10115 43800
rect 10171 43744 10239 43800
rect 10295 43744 10363 43800
rect 10419 43744 10487 43800
rect 10543 43744 10553 43800
rect 8741 43676 10553 43744
rect 8741 43620 8751 43676
rect 8807 43620 8875 43676
rect 8931 43620 8999 43676
rect 9055 43620 9123 43676
rect 9179 43620 9247 43676
rect 9303 43620 9371 43676
rect 9427 43620 9495 43676
rect 9551 43620 9619 43676
rect 9675 43620 9743 43676
rect 9799 43620 9867 43676
rect 9923 43620 9991 43676
rect 10047 43620 10115 43676
rect 10171 43620 10239 43676
rect 10295 43620 10363 43676
rect 10419 43620 10487 43676
rect 10543 43620 10553 43676
rect 8741 43552 10553 43620
rect 8741 43496 8751 43552
rect 8807 43496 8875 43552
rect 8931 43496 8999 43552
rect 9055 43496 9123 43552
rect 9179 43496 9247 43552
rect 9303 43496 9371 43552
rect 9427 43496 9495 43552
rect 9551 43496 9619 43552
rect 9675 43496 9743 43552
rect 9799 43496 9867 43552
rect 9923 43496 9991 43552
rect 10047 43496 10115 43552
rect 10171 43496 10239 43552
rect 10295 43496 10363 43552
rect 10419 43496 10487 43552
rect 10543 43496 10553 43552
rect 8741 43428 10553 43496
rect 8741 43372 8751 43428
rect 8807 43372 8875 43428
rect 8931 43372 8999 43428
rect 9055 43372 9123 43428
rect 9179 43372 9247 43428
rect 9303 43372 9371 43428
rect 9427 43372 9495 43428
rect 9551 43372 9619 43428
rect 9675 43372 9743 43428
rect 9799 43372 9867 43428
rect 9923 43372 9991 43428
rect 10047 43372 10115 43428
rect 10171 43372 10239 43428
rect 10295 43372 10363 43428
rect 10419 43372 10487 43428
rect 10543 43372 10553 43428
rect 8741 43304 10553 43372
rect 8741 43248 8751 43304
rect 8807 43248 8875 43304
rect 8931 43248 8999 43304
rect 9055 43248 9123 43304
rect 9179 43248 9247 43304
rect 9303 43248 9371 43304
rect 9427 43248 9495 43304
rect 9551 43248 9619 43304
rect 9675 43248 9743 43304
rect 9799 43248 9867 43304
rect 9923 43248 9991 43304
rect 10047 43248 10115 43304
rect 10171 43248 10239 43304
rect 10295 43248 10363 43304
rect 10419 43248 10487 43304
rect 10543 43248 10553 43304
rect 8741 43238 10553 43248
rect 12842 44544 13910 44554
rect 12842 44488 12852 44544
rect 12908 44488 12976 44544
rect 13032 44488 13100 44544
rect 13156 44488 13224 44544
rect 13280 44488 13348 44544
rect 13404 44488 13472 44544
rect 13528 44488 13596 44544
rect 13652 44488 13720 44544
rect 13776 44488 13844 44544
rect 13900 44488 13910 44544
rect 12842 44420 13910 44488
rect 12842 44364 12852 44420
rect 12908 44364 12976 44420
rect 13032 44364 13100 44420
rect 13156 44364 13224 44420
rect 13280 44364 13348 44420
rect 13404 44364 13472 44420
rect 13528 44364 13596 44420
rect 13652 44364 13720 44420
rect 13776 44364 13844 44420
rect 13900 44364 13910 44420
rect 12842 44296 13910 44364
rect 12842 44240 12852 44296
rect 12908 44240 12976 44296
rect 13032 44240 13100 44296
rect 13156 44240 13224 44296
rect 13280 44240 13348 44296
rect 13404 44240 13472 44296
rect 13528 44240 13596 44296
rect 13652 44240 13720 44296
rect 13776 44240 13844 44296
rect 13900 44240 13910 44296
rect 12842 44172 13910 44240
rect 12842 44116 12852 44172
rect 12908 44116 12976 44172
rect 13032 44116 13100 44172
rect 13156 44116 13224 44172
rect 13280 44116 13348 44172
rect 13404 44116 13472 44172
rect 13528 44116 13596 44172
rect 13652 44116 13720 44172
rect 13776 44116 13844 44172
rect 13900 44116 13910 44172
rect 12842 44048 13910 44116
rect 12842 43992 12852 44048
rect 12908 43992 12976 44048
rect 13032 43992 13100 44048
rect 13156 43992 13224 44048
rect 13280 43992 13348 44048
rect 13404 43992 13472 44048
rect 13528 43992 13596 44048
rect 13652 43992 13720 44048
rect 13776 43992 13844 44048
rect 13900 43992 13910 44048
rect 12842 43924 13910 43992
rect 12842 43868 12852 43924
rect 12908 43868 12976 43924
rect 13032 43868 13100 43924
rect 13156 43868 13224 43924
rect 13280 43868 13348 43924
rect 13404 43868 13472 43924
rect 13528 43868 13596 43924
rect 13652 43868 13720 43924
rect 13776 43868 13844 43924
rect 13900 43868 13910 43924
rect 12842 43800 13910 43868
rect 12842 43744 12852 43800
rect 12908 43744 12976 43800
rect 13032 43744 13100 43800
rect 13156 43744 13224 43800
rect 13280 43744 13348 43800
rect 13404 43744 13472 43800
rect 13528 43744 13596 43800
rect 13652 43744 13720 43800
rect 13776 43744 13844 43800
rect 13900 43744 13910 43800
rect 12842 43676 13910 43744
rect 12842 43620 12852 43676
rect 12908 43620 12976 43676
rect 13032 43620 13100 43676
rect 13156 43620 13224 43676
rect 13280 43620 13348 43676
rect 13404 43620 13472 43676
rect 13528 43620 13596 43676
rect 13652 43620 13720 43676
rect 13776 43620 13844 43676
rect 13900 43620 13910 43676
rect 12842 43552 13910 43620
rect 12842 43496 12852 43552
rect 12908 43496 12976 43552
rect 13032 43496 13100 43552
rect 13156 43496 13224 43552
rect 13280 43496 13348 43552
rect 13404 43496 13472 43552
rect 13528 43496 13596 43552
rect 13652 43496 13720 43552
rect 13776 43496 13844 43552
rect 13900 43496 13910 43552
rect 12842 43428 13910 43496
rect 12842 43372 12852 43428
rect 12908 43372 12976 43428
rect 13032 43372 13100 43428
rect 13156 43372 13224 43428
rect 13280 43372 13348 43428
rect 13404 43372 13472 43428
rect 13528 43372 13596 43428
rect 13652 43372 13720 43428
rect 13776 43372 13844 43428
rect 13900 43372 13910 43428
rect 12842 43304 13910 43372
rect 12842 43248 12852 43304
rect 12908 43248 12976 43304
rect 13032 43248 13100 43304
rect 13156 43248 13224 43304
rect 13280 43248 13348 43304
rect 13404 43248 13472 43304
rect 13528 43248 13596 43304
rect 13652 43248 13720 43304
rect 13776 43248 13844 43304
rect 13900 43248 13910 43304
rect 12842 43238 13910 43248
rect 6072 43167 6082 43223
rect 6138 43167 6148 43223
rect 5328 43100 5338 43156
rect 5394 43100 5404 43156
rect 5328 43032 5404 43100
rect 6072 43099 6148 43167
rect 6072 43043 6082 43099
rect 6138 43043 6148 43099
rect 5328 42976 5338 43032
rect 5394 42976 5404 43032
rect 5328 42908 5404 42976
rect 5328 42852 5338 42908
rect 5394 42852 5404 42908
rect 5328 42784 5404 42852
rect 5328 42728 5338 42784
rect 5394 42728 5404 42784
rect 5328 42660 5404 42728
rect 5328 42604 5338 42660
rect 5394 42604 5404 42660
rect 5328 42536 5404 42604
rect 5328 42480 5338 42536
rect 5394 42480 5404 42536
rect 5328 42412 5404 42480
rect 5328 42356 5338 42412
rect 5394 42356 5404 42412
rect 5328 42288 5404 42356
rect 5328 42232 5338 42288
rect 5394 42232 5404 42288
rect 5328 42164 5404 42232
rect 5328 42108 5338 42164
rect 5394 42108 5404 42164
rect 5328 42040 5404 42108
rect 5328 41984 5338 42040
rect 5394 41984 5404 42040
rect 5328 41916 5404 41984
rect 5328 41860 5338 41916
rect 5394 41860 5404 41916
rect 5328 41792 5404 41860
rect 5328 41736 5338 41792
rect 5394 41736 5404 41792
rect 5328 41668 5404 41736
rect 5328 41612 5338 41668
rect 5394 41612 5404 41668
rect 4584 41485 4594 41541
rect 4650 41485 4660 41541
rect 4584 41417 4660 41485
rect 4584 41361 4594 41417
rect 4650 41361 4660 41417
rect 4584 41293 4660 41361
rect 4584 41237 4594 41293
rect 4650 41237 4660 41293
rect 4584 41169 4660 41237
rect 4584 41113 4594 41169
rect 4650 41113 4660 41169
rect 4584 41045 4660 41113
rect 4584 40989 4594 41045
rect 4650 40989 4660 41045
rect 4584 40921 4660 40989
rect 4584 40865 4594 40921
rect 4650 40865 4660 40921
rect 4584 40797 4660 40865
rect 4584 40741 4594 40797
rect 4650 40741 4660 40797
rect 4584 40673 4660 40741
rect 4584 40617 4594 40673
rect 4650 40617 4660 40673
rect 4584 40549 4660 40617
rect 4584 40493 4594 40549
rect 4650 40493 4660 40549
rect 4584 40425 4660 40493
rect 4584 40369 4594 40425
rect 4650 40369 4660 40425
rect 4584 40301 4660 40369
rect 4584 40245 4594 40301
rect 4650 40245 4660 40301
rect 4584 40177 4660 40245
rect 4584 40121 4594 40177
rect 4650 40121 4660 40177
rect 4584 40053 4660 40121
rect 4584 39997 4594 40053
rect 4650 39997 4660 40053
rect 4584 39987 4660 39997
rect 4708 41541 4784 41551
rect 4708 41485 4718 41541
rect 4774 41485 4784 41541
rect 4708 41417 4784 41485
rect 5328 41544 5404 41612
rect 5328 41488 5338 41544
rect 5394 41488 5404 41544
rect 5328 41478 5404 41488
rect 5452 43032 5528 43042
rect 6072 43033 6148 43043
rect 5452 42976 5462 43032
rect 5518 42976 5528 43032
rect 5452 42908 5528 42976
rect 7552 42944 8620 42954
rect 5452 42852 5462 42908
rect 5518 42852 5528 42908
rect 5452 42784 5528 42852
rect 5452 42728 5462 42784
rect 5518 42728 5528 42784
rect 5452 42660 5528 42728
rect 5452 42604 5462 42660
rect 5518 42604 5528 42660
rect 5452 42536 5528 42604
rect 5452 42480 5462 42536
rect 5518 42480 5528 42536
rect 5452 42412 5528 42480
rect 5452 42356 5462 42412
rect 5518 42356 5528 42412
rect 5452 42288 5528 42356
rect 5452 42232 5462 42288
rect 5518 42232 5528 42288
rect 5452 42164 5528 42232
rect 5452 42108 5462 42164
rect 5518 42108 5528 42164
rect 5452 42040 5528 42108
rect 5452 41984 5462 42040
rect 5518 41984 5528 42040
rect 5452 41916 5528 41984
rect 5452 41860 5462 41916
rect 5518 41860 5528 41916
rect 5452 41792 5528 41860
rect 5452 41736 5462 41792
rect 5518 41736 5528 41792
rect 5452 41668 5528 41736
rect 5452 41612 5462 41668
rect 5518 41612 5528 41668
rect 5452 41544 5528 41612
rect 5452 41488 5462 41544
rect 5518 41488 5528 41544
rect 4708 41361 4718 41417
rect 4774 41361 4784 41417
rect 4708 41293 4784 41361
rect 4708 41237 4718 41293
rect 4774 41237 4784 41293
rect 4708 41169 4784 41237
rect 4708 41113 4718 41169
rect 4774 41113 4784 41169
rect 4708 41045 4784 41113
rect 4708 40989 4718 41045
rect 4774 40989 4784 41045
rect 4708 40921 4784 40989
rect 4708 40865 4718 40921
rect 4774 40865 4784 40921
rect 4708 40797 4784 40865
rect 4708 40741 4718 40797
rect 4774 40741 4784 40797
rect 4708 40673 4784 40741
rect 4708 40617 4718 40673
rect 4774 40617 4784 40673
rect 4708 40549 4784 40617
rect 4708 40493 4718 40549
rect 4774 40493 4784 40549
rect 4708 40425 4784 40493
rect 4708 40369 4718 40425
rect 4774 40369 4784 40425
rect 4708 40301 4784 40369
rect 4708 40245 4718 40301
rect 4774 40245 4784 40301
rect 4708 40177 4784 40245
rect 4708 40121 4718 40177
rect 4774 40121 4784 40177
rect 4708 40053 4784 40121
rect 4708 39997 4718 40053
rect 4774 39997 4784 40053
rect 4708 39929 4784 39997
rect 4708 39873 4718 39929
rect 4774 39873 4784 39929
rect 4708 39863 4784 39873
rect 4832 41417 4908 41427
rect 4832 41361 4842 41417
rect 4898 41361 4908 41417
rect 4832 41293 4908 41361
rect 5452 41420 5528 41488
rect 5452 41364 5462 41420
rect 5518 41364 5528 41420
rect 5452 41354 5528 41364
rect 5576 42908 5652 42918
rect 5576 42852 5586 42908
rect 5642 42852 5652 42908
rect 5576 42784 5652 42852
rect 7552 42888 7562 42944
rect 7618 42888 7686 42944
rect 7742 42888 7810 42944
rect 7866 42888 7934 42944
rect 7990 42888 8058 42944
rect 8114 42888 8182 42944
rect 8238 42888 8306 42944
rect 8362 42888 8430 42944
rect 8486 42888 8554 42944
rect 8610 42888 8620 42944
rect 7552 42820 8620 42888
rect 5576 42728 5586 42784
rect 5642 42728 5652 42784
rect 5576 42660 5652 42728
rect 5576 42604 5586 42660
rect 5642 42604 5652 42660
rect 5576 42536 5652 42604
rect 5576 42480 5586 42536
rect 5642 42480 5652 42536
rect 5576 42412 5652 42480
rect 5576 42356 5586 42412
rect 5642 42356 5652 42412
rect 5576 42288 5652 42356
rect 5576 42232 5586 42288
rect 5642 42232 5652 42288
rect 5576 42164 5652 42232
rect 5576 42108 5586 42164
rect 5642 42108 5652 42164
rect 5576 42040 5652 42108
rect 5576 41984 5586 42040
rect 5642 41984 5652 42040
rect 5576 41916 5652 41984
rect 5576 41860 5586 41916
rect 5642 41860 5652 41916
rect 5576 41792 5652 41860
rect 5576 41736 5586 41792
rect 5642 41736 5652 41792
rect 5576 41668 5652 41736
rect 5576 41612 5586 41668
rect 5642 41612 5652 41668
rect 5576 41544 5652 41612
rect 5576 41488 5586 41544
rect 5642 41488 5652 41544
rect 5576 41420 5652 41488
rect 5576 41364 5586 41420
rect 5642 41364 5652 41420
rect 4832 41237 4842 41293
rect 4898 41237 4908 41293
rect 4832 41169 4908 41237
rect 4832 41113 4842 41169
rect 4898 41113 4908 41169
rect 4832 41045 4908 41113
rect 4832 40989 4842 41045
rect 4898 40989 4908 41045
rect 4832 40921 4908 40989
rect 4832 40865 4842 40921
rect 4898 40865 4908 40921
rect 4832 40797 4908 40865
rect 4832 40741 4842 40797
rect 4898 40741 4908 40797
rect 4832 40673 4908 40741
rect 4832 40617 4842 40673
rect 4898 40617 4908 40673
rect 4832 40549 4908 40617
rect 4832 40493 4842 40549
rect 4898 40493 4908 40549
rect 4832 40425 4908 40493
rect 4832 40369 4842 40425
rect 4898 40369 4908 40425
rect 4832 40301 4908 40369
rect 4832 40245 4842 40301
rect 4898 40245 4908 40301
rect 4832 40177 4908 40245
rect 4832 40121 4842 40177
rect 4898 40121 4908 40177
rect 4832 40053 4908 40121
rect 4832 39997 4842 40053
rect 4898 39997 4908 40053
rect 4832 39929 4908 39997
rect 4832 39873 4842 39929
rect 4898 39873 4908 39929
rect 4832 39805 4908 39873
rect 4832 39749 4842 39805
rect 4898 39749 4908 39805
rect 4832 39739 4908 39749
rect 4956 41293 5032 41303
rect 4956 41237 4966 41293
rect 5022 41237 5032 41293
rect 4956 41169 5032 41237
rect 5576 41296 5652 41364
rect 5576 41240 5586 41296
rect 5642 41240 5652 41296
rect 5576 41230 5652 41240
rect 5700 42784 5776 42794
rect 5700 42728 5710 42784
rect 5766 42728 5776 42784
rect 5700 42660 5776 42728
rect 7552 42764 7562 42820
rect 7618 42764 7686 42820
rect 7742 42764 7810 42820
rect 7866 42764 7934 42820
rect 7990 42764 8058 42820
rect 8114 42764 8182 42820
rect 8238 42764 8306 42820
rect 8362 42764 8430 42820
rect 8486 42764 8554 42820
rect 8610 42764 8620 42820
rect 7552 42696 8620 42764
rect 5700 42604 5710 42660
rect 5766 42604 5776 42660
rect 5700 42536 5776 42604
rect 5700 42480 5710 42536
rect 5766 42480 5776 42536
rect 5700 42412 5776 42480
rect 5700 42356 5710 42412
rect 5766 42356 5776 42412
rect 5700 42288 5776 42356
rect 5700 42232 5710 42288
rect 5766 42232 5776 42288
rect 5700 42164 5776 42232
rect 5700 42108 5710 42164
rect 5766 42108 5776 42164
rect 5700 42040 5776 42108
rect 5700 41984 5710 42040
rect 5766 41984 5776 42040
rect 5700 41916 5776 41984
rect 5700 41860 5710 41916
rect 5766 41860 5776 41916
rect 5700 41792 5776 41860
rect 5700 41736 5710 41792
rect 5766 41736 5776 41792
rect 5700 41668 5776 41736
rect 5700 41612 5710 41668
rect 5766 41612 5776 41668
rect 5700 41544 5776 41612
rect 5700 41488 5710 41544
rect 5766 41488 5776 41544
rect 5700 41420 5776 41488
rect 5700 41364 5710 41420
rect 5766 41364 5776 41420
rect 5700 41296 5776 41364
rect 5700 41240 5710 41296
rect 5766 41240 5776 41296
rect 4956 41113 4966 41169
rect 5022 41113 5032 41169
rect 4956 41045 5032 41113
rect 4956 40989 4966 41045
rect 5022 40989 5032 41045
rect 4956 40921 5032 40989
rect 4956 40865 4966 40921
rect 5022 40865 5032 40921
rect 4956 40797 5032 40865
rect 4956 40741 4966 40797
rect 5022 40741 5032 40797
rect 4956 40673 5032 40741
rect 4956 40617 4966 40673
rect 5022 40617 5032 40673
rect 4956 40549 5032 40617
rect 4956 40493 4966 40549
rect 5022 40493 5032 40549
rect 4956 40425 5032 40493
rect 4956 40369 4966 40425
rect 5022 40369 5032 40425
rect 4956 40301 5032 40369
rect 4956 40245 4966 40301
rect 5022 40245 5032 40301
rect 4956 40177 5032 40245
rect 4956 40121 4966 40177
rect 5022 40121 5032 40177
rect 4956 40053 5032 40121
rect 4956 39997 4966 40053
rect 5022 39997 5032 40053
rect 4956 39929 5032 39997
rect 4956 39873 4966 39929
rect 5022 39873 5032 39929
rect 4956 39805 5032 39873
rect 4956 39749 4966 39805
rect 5022 39749 5032 39805
rect 4956 39681 5032 39749
rect 4956 39625 4966 39681
rect 5022 39625 5032 39681
rect 4956 39615 5032 39625
rect 5080 41169 5156 41179
rect 5080 41113 5090 41169
rect 5146 41113 5156 41169
rect 5080 41045 5156 41113
rect 5700 41172 5776 41240
rect 5700 41116 5710 41172
rect 5766 41116 5776 41172
rect 5700 41106 5776 41116
rect 5824 42660 5900 42670
rect 5824 42604 5834 42660
rect 5890 42604 5900 42660
rect 5824 42536 5900 42604
rect 7552 42640 7562 42696
rect 7618 42640 7686 42696
rect 7742 42640 7810 42696
rect 7866 42640 7934 42696
rect 7990 42640 8058 42696
rect 8114 42640 8182 42696
rect 8238 42640 8306 42696
rect 8362 42640 8430 42696
rect 8486 42640 8554 42696
rect 8610 42640 8620 42696
rect 7552 42572 8620 42640
rect 5824 42480 5834 42536
rect 5890 42480 5900 42536
rect 5824 42412 5900 42480
rect 5824 42356 5834 42412
rect 5890 42356 5900 42412
rect 5824 42288 5900 42356
rect 5824 42232 5834 42288
rect 5890 42232 5900 42288
rect 5824 42164 5900 42232
rect 5824 42108 5834 42164
rect 5890 42108 5900 42164
rect 5824 42040 5900 42108
rect 5824 41984 5834 42040
rect 5890 41984 5900 42040
rect 5824 41916 5900 41984
rect 5824 41860 5834 41916
rect 5890 41860 5900 41916
rect 5824 41792 5900 41860
rect 5824 41736 5834 41792
rect 5890 41736 5900 41792
rect 5824 41668 5900 41736
rect 5824 41612 5834 41668
rect 5890 41612 5900 41668
rect 5824 41544 5900 41612
rect 5824 41488 5834 41544
rect 5890 41488 5900 41544
rect 5824 41420 5900 41488
rect 5824 41364 5834 41420
rect 5890 41364 5900 41420
rect 5824 41296 5900 41364
rect 5824 41240 5834 41296
rect 5890 41240 5900 41296
rect 5824 41172 5900 41240
rect 5824 41116 5834 41172
rect 5890 41116 5900 41172
rect 5080 40989 5090 41045
rect 5146 40989 5156 41045
rect 5080 40921 5156 40989
rect 5080 40865 5090 40921
rect 5146 40865 5156 40921
rect 5080 40797 5156 40865
rect 5080 40741 5090 40797
rect 5146 40741 5156 40797
rect 5080 40673 5156 40741
rect 5080 40617 5090 40673
rect 5146 40617 5156 40673
rect 5080 40549 5156 40617
rect 5080 40493 5090 40549
rect 5146 40493 5156 40549
rect 5080 40425 5156 40493
rect 5080 40369 5090 40425
rect 5146 40369 5156 40425
rect 5080 40301 5156 40369
rect 5080 40245 5090 40301
rect 5146 40245 5156 40301
rect 5080 40177 5156 40245
rect 5080 40121 5090 40177
rect 5146 40121 5156 40177
rect 5080 40053 5156 40121
rect 5080 39997 5090 40053
rect 5146 39997 5156 40053
rect 5080 39929 5156 39997
rect 5080 39873 5090 39929
rect 5146 39873 5156 39929
rect 5080 39805 5156 39873
rect 5080 39749 5090 39805
rect 5146 39749 5156 39805
rect 5080 39681 5156 39749
rect 5080 39625 5090 39681
rect 5146 39625 5156 39681
rect 5080 39557 5156 39625
rect 5080 39501 5090 39557
rect 5146 39501 5156 39557
rect 5080 39491 5156 39501
rect 5204 41045 5280 41055
rect 5204 40989 5214 41045
rect 5270 40989 5280 41045
rect 5204 40921 5280 40989
rect 5824 41048 5900 41116
rect 5824 40992 5834 41048
rect 5890 40992 5900 41048
rect 5824 40982 5900 40992
rect 5948 42536 6024 42546
rect 5948 42480 5958 42536
rect 6014 42480 6024 42536
rect 5948 42412 6024 42480
rect 7552 42516 7562 42572
rect 7618 42516 7686 42572
rect 7742 42516 7810 42572
rect 7866 42516 7934 42572
rect 7990 42516 8058 42572
rect 8114 42516 8182 42572
rect 8238 42516 8306 42572
rect 8362 42516 8430 42572
rect 8486 42516 8554 42572
rect 8610 42516 8620 42572
rect 7552 42448 8620 42516
rect 5948 42356 5958 42412
rect 6014 42356 6024 42412
rect 5948 42288 6024 42356
rect 5948 42232 5958 42288
rect 6014 42232 6024 42288
rect 5948 42164 6024 42232
rect 5948 42108 5958 42164
rect 6014 42108 6024 42164
rect 5948 42040 6024 42108
rect 5948 41984 5958 42040
rect 6014 41984 6024 42040
rect 5948 41916 6024 41984
rect 5948 41860 5958 41916
rect 6014 41860 6024 41916
rect 5948 41792 6024 41860
rect 5948 41736 5958 41792
rect 6014 41736 6024 41792
rect 5948 41668 6024 41736
rect 5948 41612 5958 41668
rect 6014 41612 6024 41668
rect 5948 41544 6024 41612
rect 5948 41488 5958 41544
rect 6014 41488 6024 41544
rect 5948 41420 6024 41488
rect 5948 41364 5958 41420
rect 6014 41364 6024 41420
rect 5948 41296 6024 41364
rect 5948 41240 5958 41296
rect 6014 41240 6024 41296
rect 5948 41172 6024 41240
rect 5948 41116 5958 41172
rect 6014 41116 6024 41172
rect 5948 41048 6024 41116
rect 5948 40992 5958 41048
rect 6014 40992 6024 41048
rect 5204 40865 5214 40921
rect 5270 40865 5280 40921
rect 5204 40797 5280 40865
rect 5204 40741 5214 40797
rect 5270 40741 5280 40797
rect 5204 40673 5280 40741
rect 5204 40617 5214 40673
rect 5270 40617 5280 40673
rect 5204 40549 5280 40617
rect 5204 40493 5214 40549
rect 5270 40493 5280 40549
rect 5204 40425 5280 40493
rect 5204 40369 5214 40425
rect 5270 40369 5280 40425
rect 5204 40301 5280 40369
rect 5204 40245 5214 40301
rect 5270 40245 5280 40301
rect 5204 40177 5280 40245
rect 5204 40121 5214 40177
rect 5270 40121 5280 40177
rect 5204 40053 5280 40121
rect 5204 39997 5214 40053
rect 5270 39997 5280 40053
rect 5204 39929 5280 39997
rect 5204 39873 5214 39929
rect 5270 39873 5280 39929
rect 5204 39805 5280 39873
rect 5204 39749 5214 39805
rect 5270 39749 5280 39805
rect 5204 39681 5280 39749
rect 5204 39625 5214 39681
rect 5270 39625 5280 39681
rect 5204 39557 5280 39625
rect 5204 39501 5214 39557
rect 5270 39501 5280 39557
rect 5204 39433 5280 39501
rect 5204 39377 5214 39433
rect 5270 39377 5280 39433
rect 5204 39367 5280 39377
rect 5328 40921 5404 40931
rect 5328 40865 5338 40921
rect 5394 40865 5404 40921
rect 5328 40797 5404 40865
rect 5948 40924 6024 40992
rect 5948 40868 5958 40924
rect 6014 40868 6024 40924
rect 5948 40858 6024 40868
rect 6072 42412 6148 42422
rect 6072 42356 6082 42412
rect 6138 42356 6148 42412
rect 6072 42288 6148 42356
rect 6072 42232 6082 42288
rect 6138 42232 6148 42288
rect 6072 42164 6148 42232
rect 6072 42108 6082 42164
rect 6138 42108 6148 42164
rect 6072 42040 6148 42108
rect 6072 41984 6082 42040
rect 6138 41984 6148 42040
rect 6072 41916 6148 41984
rect 6072 41860 6082 41916
rect 6138 41860 6148 41916
rect 6072 41792 6148 41860
rect 6072 41736 6082 41792
rect 6138 41736 6148 41792
rect 6072 41668 6148 41736
rect 6072 41612 6082 41668
rect 6138 41612 6148 41668
rect 7552 42392 7562 42448
rect 7618 42392 7686 42448
rect 7742 42392 7810 42448
rect 7866 42392 7934 42448
rect 7990 42392 8058 42448
rect 8114 42392 8182 42448
rect 8238 42392 8306 42448
rect 8362 42392 8430 42448
rect 8486 42392 8554 42448
rect 8610 42392 8620 42448
rect 7552 42324 8620 42392
rect 7552 42268 7562 42324
rect 7618 42268 7686 42324
rect 7742 42268 7810 42324
rect 7866 42268 7934 42324
rect 7990 42268 8058 42324
rect 8114 42268 8182 42324
rect 8238 42268 8306 42324
rect 8362 42268 8430 42324
rect 8486 42268 8554 42324
rect 8610 42268 8620 42324
rect 7552 42200 8620 42268
rect 7552 42144 7562 42200
rect 7618 42144 7686 42200
rect 7742 42144 7810 42200
rect 7866 42144 7934 42200
rect 7990 42144 8058 42200
rect 8114 42144 8182 42200
rect 8238 42144 8306 42200
rect 8362 42144 8430 42200
rect 8486 42144 8554 42200
rect 8610 42144 8620 42200
rect 7552 42076 8620 42144
rect 7552 42020 7562 42076
rect 7618 42020 7686 42076
rect 7742 42020 7810 42076
rect 7866 42020 7934 42076
rect 7990 42020 8058 42076
rect 8114 42020 8182 42076
rect 8238 42020 8306 42076
rect 8362 42020 8430 42076
rect 8486 42020 8554 42076
rect 8610 42020 8620 42076
rect 7552 41952 8620 42020
rect 7552 41896 7562 41952
rect 7618 41896 7686 41952
rect 7742 41896 7810 41952
rect 7866 41896 7934 41952
rect 7990 41896 8058 41952
rect 8114 41896 8182 41952
rect 8238 41896 8306 41952
rect 8362 41896 8430 41952
rect 8486 41896 8554 41952
rect 8610 41896 8620 41952
rect 7552 41828 8620 41896
rect 7552 41772 7562 41828
rect 7618 41772 7686 41828
rect 7742 41772 7810 41828
rect 7866 41772 7934 41828
rect 7990 41772 8058 41828
rect 8114 41772 8182 41828
rect 8238 41772 8306 41828
rect 8362 41772 8430 41828
rect 8486 41772 8554 41828
rect 8610 41772 8620 41828
rect 7552 41704 8620 41772
rect 7552 41648 7562 41704
rect 7618 41648 7686 41704
rect 7742 41648 7810 41704
rect 7866 41648 7934 41704
rect 7990 41648 8058 41704
rect 8114 41648 8182 41704
rect 8238 41648 8306 41704
rect 8362 41648 8430 41704
rect 8486 41648 8554 41704
rect 8610 41648 8620 41704
rect 7552 41638 8620 41648
rect 10669 42944 12481 42954
rect 10669 42888 10679 42944
rect 10735 42888 10803 42944
rect 10859 42888 10927 42944
rect 10983 42888 11051 42944
rect 11107 42888 11175 42944
rect 11231 42888 11299 42944
rect 11355 42888 11423 42944
rect 11479 42888 11547 42944
rect 11603 42888 11671 42944
rect 11727 42888 11795 42944
rect 11851 42888 11919 42944
rect 11975 42888 12043 42944
rect 12099 42888 12167 42944
rect 12223 42888 12291 42944
rect 12347 42888 12415 42944
rect 12471 42888 12481 42944
rect 10669 42820 12481 42888
rect 10669 42764 10679 42820
rect 10735 42764 10803 42820
rect 10859 42764 10927 42820
rect 10983 42764 11051 42820
rect 11107 42764 11175 42820
rect 11231 42764 11299 42820
rect 11355 42764 11423 42820
rect 11479 42764 11547 42820
rect 11603 42764 11671 42820
rect 11727 42764 11795 42820
rect 11851 42764 11919 42820
rect 11975 42764 12043 42820
rect 12099 42764 12167 42820
rect 12223 42764 12291 42820
rect 12347 42764 12415 42820
rect 12471 42764 12481 42820
rect 10669 42696 12481 42764
rect 10669 42640 10679 42696
rect 10735 42640 10803 42696
rect 10859 42640 10927 42696
rect 10983 42640 11051 42696
rect 11107 42640 11175 42696
rect 11231 42640 11299 42696
rect 11355 42640 11423 42696
rect 11479 42640 11547 42696
rect 11603 42640 11671 42696
rect 11727 42640 11795 42696
rect 11851 42640 11919 42696
rect 11975 42640 12043 42696
rect 12099 42640 12167 42696
rect 12223 42640 12291 42696
rect 12347 42640 12415 42696
rect 12471 42640 12481 42696
rect 10669 42572 12481 42640
rect 10669 42516 10679 42572
rect 10735 42516 10803 42572
rect 10859 42516 10927 42572
rect 10983 42516 11051 42572
rect 11107 42516 11175 42572
rect 11231 42516 11299 42572
rect 11355 42516 11423 42572
rect 11479 42516 11547 42572
rect 11603 42516 11671 42572
rect 11727 42516 11795 42572
rect 11851 42516 11919 42572
rect 11975 42516 12043 42572
rect 12099 42516 12167 42572
rect 12223 42516 12291 42572
rect 12347 42516 12415 42572
rect 12471 42516 12481 42572
rect 10669 42448 12481 42516
rect 10669 42392 10679 42448
rect 10735 42392 10803 42448
rect 10859 42392 10927 42448
rect 10983 42392 11051 42448
rect 11107 42392 11175 42448
rect 11231 42392 11299 42448
rect 11355 42392 11423 42448
rect 11479 42392 11547 42448
rect 11603 42392 11671 42448
rect 11727 42392 11795 42448
rect 11851 42392 11919 42448
rect 11975 42392 12043 42448
rect 12099 42392 12167 42448
rect 12223 42392 12291 42448
rect 12347 42392 12415 42448
rect 12471 42392 12481 42448
rect 10669 42324 12481 42392
rect 10669 42268 10679 42324
rect 10735 42268 10803 42324
rect 10859 42268 10927 42324
rect 10983 42268 11051 42324
rect 11107 42268 11175 42324
rect 11231 42268 11299 42324
rect 11355 42268 11423 42324
rect 11479 42268 11547 42324
rect 11603 42268 11671 42324
rect 11727 42268 11795 42324
rect 11851 42268 11919 42324
rect 11975 42268 12043 42324
rect 12099 42268 12167 42324
rect 12223 42268 12291 42324
rect 12347 42268 12415 42324
rect 12471 42268 12481 42324
rect 10669 42200 12481 42268
rect 10669 42144 10679 42200
rect 10735 42144 10803 42200
rect 10859 42144 10927 42200
rect 10983 42144 11051 42200
rect 11107 42144 11175 42200
rect 11231 42144 11299 42200
rect 11355 42144 11423 42200
rect 11479 42144 11547 42200
rect 11603 42144 11671 42200
rect 11727 42144 11795 42200
rect 11851 42144 11919 42200
rect 11975 42144 12043 42200
rect 12099 42144 12167 42200
rect 12223 42144 12291 42200
rect 12347 42144 12415 42200
rect 12471 42144 12481 42200
rect 10669 42076 12481 42144
rect 10669 42020 10679 42076
rect 10735 42020 10803 42076
rect 10859 42020 10927 42076
rect 10983 42020 11051 42076
rect 11107 42020 11175 42076
rect 11231 42020 11299 42076
rect 11355 42020 11423 42076
rect 11479 42020 11547 42076
rect 11603 42020 11671 42076
rect 11727 42020 11795 42076
rect 11851 42020 11919 42076
rect 11975 42020 12043 42076
rect 12099 42020 12167 42076
rect 12223 42020 12291 42076
rect 12347 42020 12415 42076
rect 12471 42020 12481 42076
rect 10669 41952 12481 42020
rect 10669 41896 10679 41952
rect 10735 41896 10803 41952
rect 10859 41896 10927 41952
rect 10983 41896 11051 41952
rect 11107 41896 11175 41952
rect 11231 41896 11299 41952
rect 11355 41896 11423 41952
rect 11479 41896 11547 41952
rect 11603 41896 11671 41952
rect 11727 41896 11795 41952
rect 11851 41896 11919 41952
rect 11975 41896 12043 41952
rect 12099 41896 12167 41952
rect 12223 41896 12291 41952
rect 12347 41896 12415 41952
rect 12471 41896 12481 41952
rect 10669 41828 12481 41896
rect 10669 41772 10679 41828
rect 10735 41772 10803 41828
rect 10859 41772 10927 41828
rect 10983 41772 11051 41828
rect 11107 41772 11175 41828
rect 11231 41772 11299 41828
rect 11355 41772 11423 41828
rect 11479 41772 11547 41828
rect 11603 41772 11671 41828
rect 11727 41772 11795 41828
rect 11851 41772 11919 41828
rect 11975 41772 12043 41828
rect 12099 41772 12167 41828
rect 12223 41772 12291 41828
rect 12347 41772 12415 41828
rect 12471 41772 12481 41828
rect 10669 41704 12481 41772
rect 10669 41648 10679 41704
rect 10735 41648 10803 41704
rect 10859 41648 10927 41704
rect 10983 41648 11051 41704
rect 11107 41648 11175 41704
rect 11231 41648 11299 41704
rect 11355 41648 11423 41704
rect 11479 41648 11547 41704
rect 11603 41648 11671 41704
rect 11727 41648 11795 41704
rect 11851 41648 11919 41704
rect 11975 41648 12043 41704
rect 12099 41648 12167 41704
rect 12223 41648 12291 41704
rect 12347 41648 12415 41704
rect 12471 41648 12481 41704
rect 10669 41638 12481 41648
rect 6072 41544 6148 41612
rect 6072 41488 6082 41544
rect 6138 41488 6148 41544
rect 6072 41420 6148 41488
rect 6072 41364 6082 41420
rect 6138 41364 6148 41420
rect 6072 41296 6148 41364
rect 6072 41240 6082 41296
rect 6138 41240 6148 41296
rect 6072 41172 6148 41240
rect 6072 41116 6082 41172
rect 6138 41116 6148 41172
rect 6072 41048 6148 41116
rect 6072 40992 6082 41048
rect 6138 40992 6148 41048
rect 6072 40924 6148 40992
rect 6072 40868 6082 40924
rect 6138 40868 6148 40924
rect 5328 40741 5338 40797
rect 5394 40741 5404 40797
rect 5328 40673 5404 40741
rect 5328 40617 5338 40673
rect 5394 40617 5404 40673
rect 5328 40549 5404 40617
rect 5328 40493 5338 40549
rect 5394 40493 5404 40549
rect 5328 40425 5404 40493
rect 5328 40369 5338 40425
rect 5394 40369 5404 40425
rect 5328 40301 5404 40369
rect 5328 40245 5338 40301
rect 5394 40245 5404 40301
rect 5328 40177 5404 40245
rect 5328 40121 5338 40177
rect 5394 40121 5404 40177
rect 5328 40053 5404 40121
rect 5328 39997 5338 40053
rect 5394 39997 5404 40053
rect 5328 39929 5404 39997
rect 5328 39873 5338 39929
rect 5394 39873 5404 39929
rect 5328 39805 5404 39873
rect 5328 39749 5338 39805
rect 5394 39749 5404 39805
rect 5328 39681 5404 39749
rect 5328 39625 5338 39681
rect 5394 39625 5404 39681
rect 5328 39557 5404 39625
rect 5328 39501 5338 39557
rect 5394 39501 5404 39557
rect 5328 39433 5404 39501
rect 5328 39377 5338 39433
rect 5394 39377 5404 39433
rect 5328 39309 5404 39377
rect 5328 39253 5338 39309
rect 5394 39253 5404 39309
rect 5328 39243 5404 39253
rect 5452 40797 5528 40807
rect 5452 40741 5462 40797
rect 5518 40741 5528 40797
rect 5452 40673 5528 40741
rect 6072 40800 6148 40868
rect 6072 40744 6082 40800
rect 6138 40744 6148 40800
rect 6072 40734 6148 40744
rect 7552 41344 8620 41354
rect 7552 41288 7562 41344
rect 7618 41288 7686 41344
rect 7742 41288 7810 41344
rect 7866 41288 7934 41344
rect 7990 41288 8058 41344
rect 8114 41288 8182 41344
rect 8238 41288 8306 41344
rect 8362 41288 8430 41344
rect 8486 41288 8554 41344
rect 8610 41288 8620 41344
rect 7552 41220 8620 41288
rect 7552 41164 7562 41220
rect 7618 41164 7686 41220
rect 7742 41164 7810 41220
rect 7866 41164 7934 41220
rect 7990 41164 8058 41220
rect 8114 41164 8182 41220
rect 8238 41164 8306 41220
rect 8362 41164 8430 41220
rect 8486 41164 8554 41220
rect 8610 41164 8620 41220
rect 7552 41096 8620 41164
rect 7552 41040 7562 41096
rect 7618 41040 7686 41096
rect 7742 41040 7810 41096
rect 7866 41040 7934 41096
rect 7990 41040 8058 41096
rect 8114 41040 8182 41096
rect 8238 41040 8306 41096
rect 8362 41040 8430 41096
rect 8486 41040 8554 41096
rect 8610 41040 8620 41096
rect 7552 40972 8620 41040
rect 7552 40916 7562 40972
rect 7618 40916 7686 40972
rect 7742 40916 7810 40972
rect 7866 40916 7934 40972
rect 7990 40916 8058 40972
rect 8114 40916 8182 40972
rect 8238 40916 8306 40972
rect 8362 40916 8430 40972
rect 8486 40916 8554 40972
rect 8610 40916 8620 40972
rect 7552 40848 8620 40916
rect 7552 40792 7562 40848
rect 7618 40792 7686 40848
rect 7742 40792 7810 40848
rect 7866 40792 7934 40848
rect 7990 40792 8058 40848
rect 8114 40792 8182 40848
rect 8238 40792 8306 40848
rect 8362 40792 8430 40848
rect 8486 40792 8554 40848
rect 8610 40792 8620 40848
rect 7552 40724 8620 40792
rect 5452 40617 5462 40673
rect 5518 40617 5528 40673
rect 5452 40549 5528 40617
rect 5452 40493 5462 40549
rect 5518 40493 5528 40549
rect 5452 40425 5528 40493
rect 5452 40369 5462 40425
rect 5518 40369 5528 40425
rect 5452 40301 5528 40369
rect 5452 40245 5462 40301
rect 5518 40245 5528 40301
rect 5452 40177 5528 40245
rect 5452 40121 5462 40177
rect 5518 40121 5528 40177
rect 5452 40053 5528 40121
rect 5452 39997 5462 40053
rect 5518 39997 5528 40053
rect 5452 39929 5528 39997
rect 5452 39873 5462 39929
rect 5518 39873 5528 39929
rect 5452 39805 5528 39873
rect 5452 39749 5462 39805
rect 5518 39749 5528 39805
rect 5452 39681 5528 39749
rect 5452 39625 5462 39681
rect 5518 39625 5528 39681
rect 5452 39557 5528 39625
rect 5452 39501 5462 39557
rect 5518 39501 5528 39557
rect 5452 39433 5528 39501
rect 5452 39377 5462 39433
rect 5518 39377 5528 39433
rect 5452 39309 5528 39377
rect 5452 39253 5462 39309
rect 5518 39253 5528 39309
rect 5452 39185 5528 39253
rect 5452 39129 5462 39185
rect 5518 39129 5528 39185
rect 5452 39119 5528 39129
rect 5576 40673 5652 40683
rect 5576 40617 5586 40673
rect 5642 40617 5652 40673
rect 5576 40549 5652 40617
rect 7552 40668 7562 40724
rect 7618 40668 7686 40724
rect 7742 40668 7810 40724
rect 7866 40668 7934 40724
rect 7990 40668 8058 40724
rect 8114 40668 8182 40724
rect 8238 40668 8306 40724
rect 8362 40668 8430 40724
rect 8486 40668 8554 40724
rect 8610 40668 8620 40724
rect 7552 40600 8620 40668
rect 5576 40493 5586 40549
rect 5642 40493 5652 40549
rect 5576 40425 5652 40493
rect 5576 40369 5586 40425
rect 5642 40369 5652 40425
rect 5576 40301 5652 40369
rect 5576 40245 5586 40301
rect 5642 40245 5652 40301
rect 5576 40177 5652 40245
rect 5576 40121 5586 40177
rect 5642 40121 5652 40177
rect 5576 40053 5652 40121
rect 5576 39997 5586 40053
rect 5642 39997 5652 40053
rect 5576 39929 5652 39997
rect 5576 39873 5586 39929
rect 5642 39873 5652 39929
rect 5576 39805 5652 39873
rect 5576 39749 5586 39805
rect 5642 39749 5652 39805
rect 5576 39681 5652 39749
rect 5576 39625 5586 39681
rect 5642 39625 5652 39681
rect 5576 39557 5652 39625
rect 5576 39501 5586 39557
rect 5642 39501 5652 39557
rect 5576 39433 5652 39501
rect 5576 39377 5586 39433
rect 5642 39377 5652 39433
rect 5576 39309 5652 39377
rect 5576 39253 5586 39309
rect 5642 39253 5652 39309
rect 5576 39185 5652 39253
rect 5576 39129 5586 39185
rect 5642 39129 5652 39185
rect 5576 39061 5652 39129
rect 5576 39005 5586 39061
rect 5642 39005 5652 39061
rect 5576 38995 5652 39005
rect 5700 40549 5776 40559
rect 5700 40493 5710 40549
rect 5766 40493 5776 40549
rect 5700 40425 5776 40493
rect 7552 40544 7562 40600
rect 7618 40544 7686 40600
rect 7742 40544 7810 40600
rect 7866 40544 7934 40600
rect 7990 40544 8058 40600
rect 8114 40544 8182 40600
rect 8238 40544 8306 40600
rect 8362 40544 8430 40600
rect 8486 40544 8554 40600
rect 8610 40544 8620 40600
rect 7552 40476 8620 40544
rect 5700 40369 5710 40425
rect 5766 40369 5776 40425
rect 5700 40301 5776 40369
rect 5700 40245 5710 40301
rect 5766 40245 5776 40301
rect 5700 40177 5776 40245
rect 5700 40121 5710 40177
rect 5766 40121 5776 40177
rect 5700 40053 5776 40121
rect 5700 39997 5710 40053
rect 5766 39997 5776 40053
rect 5700 39929 5776 39997
rect 5700 39873 5710 39929
rect 5766 39873 5776 39929
rect 5700 39805 5776 39873
rect 5700 39749 5710 39805
rect 5766 39749 5776 39805
rect 5700 39681 5776 39749
rect 5700 39625 5710 39681
rect 5766 39625 5776 39681
rect 5700 39557 5776 39625
rect 5700 39501 5710 39557
rect 5766 39501 5776 39557
rect 5700 39433 5776 39501
rect 5700 39377 5710 39433
rect 5766 39377 5776 39433
rect 5700 39309 5776 39377
rect 5700 39253 5710 39309
rect 5766 39253 5776 39309
rect 5700 39185 5776 39253
rect 5700 39129 5710 39185
rect 5766 39129 5776 39185
rect 5700 39061 5776 39129
rect 5700 39005 5710 39061
rect 5766 39005 5776 39061
rect 5700 38937 5776 39005
rect 5700 38881 5710 38937
rect 5766 38881 5776 38937
rect 5700 38871 5776 38881
rect 5824 40425 5900 40435
rect 5824 40369 5834 40425
rect 5890 40369 5900 40425
rect 5824 40301 5900 40369
rect 7552 40420 7562 40476
rect 7618 40420 7686 40476
rect 7742 40420 7810 40476
rect 7866 40420 7934 40476
rect 7990 40420 8058 40476
rect 8114 40420 8182 40476
rect 8238 40420 8306 40476
rect 8362 40420 8430 40476
rect 8486 40420 8554 40476
rect 8610 40420 8620 40476
rect 7552 40352 8620 40420
rect 5824 40245 5834 40301
rect 5890 40245 5900 40301
rect 5824 40177 5900 40245
rect 5824 40121 5834 40177
rect 5890 40121 5900 40177
rect 5824 40053 5900 40121
rect 5824 39997 5834 40053
rect 5890 39997 5900 40053
rect 5824 39929 5900 39997
rect 5824 39873 5834 39929
rect 5890 39873 5900 39929
rect 5824 39805 5900 39873
rect 5824 39749 5834 39805
rect 5890 39749 5900 39805
rect 5824 39681 5900 39749
rect 5824 39625 5834 39681
rect 5890 39625 5900 39681
rect 5824 39557 5900 39625
rect 5824 39501 5834 39557
rect 5890 39501 5900 39557
rect 5824 39433 5900 39501
rect 5824 39377 5834 39433
rect 5890 39377 5900 39433
rect 5824 39309 5900 39377
rect 5824 39253 5834 39309
rect 5890 39253 5900 39309
rect 5824 39185 5900 39253
rect 5824 39129 5834 39185
rect 5890 39129 5900 39185
rect 5824 39061 5900 39129
rect 5824 39005 5834 39061
rect 5890 39005 5900 39061
rect 5824 38937 5900 39005
rect 5824 38881 5834 38937
rect 5890 38881 5900 38937
rect 5824 38813 5900 38881
rect 5824 38757 5834 38813
rect 5890 38757 5900 38813
rect 5824 38747 5900 38757
rect 5948 40301 6024 40311
rect 5948 40245 5958 40301
rect 6014 40245 6024 40301
rect 5948 40177 6024 40245
rect 7552 40296 7562 40352
rect 7618 40296 7686 40352
rect 7742 40296 7810 40352
rect 7866 40296 7934 40352
rect 7990 40296 8058 40352
rect 8114 40296 8182 40352
rect 8238 40296 8306 40352
rect 8362 40296 8430 40352
rect 8486 40296 8554 40352
rect 8610 40296 8620 40352
rect 7552 40228 8620 40296
rect 5948 40121 5958 40177
rect 6014 40121 6024 40177
rect 5948 40053 6024 40121
rect 5948 39997 5958 40053
rect 6014 39997 6024 40053
rect 5948 39929 6024 39997
rect 5948 39873 5958 39929
rect 6014 39873 6024 39929
rect 5948 39805 6024 39873
rect 5948 39749 5958 39805
rect 6014 39749 6024 39805
rect 5948 39681 6024 39749
rect 5948 39625 5958 39681
rect 6014 39625 6024 39681
rect 5948 39557 6024 39625
rect 5948 39501 5958 39557
rect 6014 39501 6024 39557
rect 5948 39433 6024 39501
rect 5948 39377 5958 39433
rect 6014 39377 6024 39433
rect 5948 39309 6024 39377
rect 5948 39253 5958 39309
rect 6014 39253 6024 39309
rect 5948 39185 6024 39253
rect 5948 39129 5958 39185
rect 6014 39129 6024 39185
rect 5948 39061 6024 39129
rect 5948 39005 5958 39061
rect 6014 39005 6024 39061
rect 5948 38937 6024 39005
rect 5948 38881 5958 38937
rect 6014 38881 6024 38937
rect 5948 38813 6024 38881
rect 5948 38757 5958 38813
rect 6014 38757 6024 38813
rect 5948 38689 6024 38757
rect 5948 38633 5958 38689
rect 6014 38633 6024 38689
rect 5948 38623 6024 38633
rect 6072 40177 6148 40187
rect 6072 40121 6082 40177
rect 6138 40121 6148 40177
rect 6072 40053 6148 40121
rect 6072 39997 6082 40053
rect 6138 39997 6148 40053
rect 7552 40172 7562 40228
rect 7618 40172 7686 40228
rect 7742 40172 7810 40228
rect 7866 40172 7934 40228
rect 7990 40172 8058 40228
rect 8114 40172 8182 40228
rect 8238 40172 8306 40228
rect 8362 40172 8430 40228
rect 8486 40172 8554 40228
rect 8610 40172 8620 40228
rect 7552 40104 8620 40172
rect 7552 40048 7562 40104
rect 7618 40048 7686 40104
rect 7742 40048 7810 40104
rect 7866 40048 7934 40104
rect 7990 40048 8058 40104
rect 8114 40048 8182 40104
rect 8238 40048 8306 40104
rect 8362 40048 8430 40104
rect 8486 40048 8554 40104
rect 8610 40048 8620 40104
rect 7552 40038 8620 40048
rect 10669 41344 12481 41354
rect 10669 41288 10679 41344
rect 10735 41288 10803 41344
rect 10859 41288 10927 41344
rect 10983 41288 11051 41344
rect 11107 41288 11175 41344
rect 11231 41288 11299 41344
rect 11355 41288 11423 41344
rect 11479 41288 11547 41344
rect 11603 41288 11671 41344
rect 11727 41288 11795 41344
rect 11851 41288 11919 41344
rect 11975 41288 12043 41344
rect 12099 41288 12167 41344
rect 12223 41288 12291 41344
rect 12347 41288 12415 41344
rect 12471 41288 12481 41344
rect 10669 41220 12481 41288
rect 10669 41164 10679 41220
rect 10735 41164 10803 41220
rect 10859 41164 10927 41220
rect 10983 41164 11051 41220
rect 11107 41164 11175 41220
rect 11231 41164 11299 41220
rect 11355 41164 11423 41220
rect 11479 41164 11547 41220
rect 11603 41164 11671 41220
rect 11727 41164 11795 41220
rect 11851 41164 11919 41220
rect 11975 41164 12043 41220
rect 12099 41164 12167 41220
rect 12223 41164 12291 41220
rect 12347 41164 12415 41220
rect 12471 41164 12481 41220
rect 10669 41096 12481 41164
rect 10669 41040 10679 41096
rect 10735 41040 10803 41096
rect 10859 41040 10927 41096
rect 10983 41040 11051 41096
rect 11107 41040 11175 41096
rect 11231 41040 11299 41096
rect 11355 41040 11423 41096
rect 11479 41040 11547 41096
rect 11603 41040 11671 41096
rect 11727 41040 11795 41096
rect 11851 41040 11919 41096
rect 11975 41040 12043 41096
rect 12099 41040 12167 41096
rect 12223 41040 12291 41096
rect 12347 41040 12415 41096
rect 12471 41040 12481 41096
rect 10669 40972 12481 41040
rect 10669 40916 10679 40972
rect 10735 40916 10803 40972
rect 10859 40916 10927 40972
rect 10983 40916 11051 40972
rect 11107 40916 11175 40972
rect 11231 40916 11299 40972
rect 11355 40916 11423 40972
rect 11479 40916 11547 40972
rect 11603 40916 11671 40972
rect 11727 40916 11795 40972
rect 11851 40916 11919 40972
rect 11975 40916 12043 40972
rect 12099 40916 12167 40972
rect 12223 40916 12291 40972
rect 12347 40916 12415 40972
rect 12471 40916 12481 40972
rect 10669 40848 12481 40916
rect 10669 40792 10679 40848
rect 10735 40792 10803 40848
rect 10859 40792 10927 40848
rect 10983 40792 11051 40848
rect 11107 40792 11175 40848
rect 11231 40792 11299 40848
rect 11355 40792 11423 40848
rect 11479 40792 11547 40848
rect 11603 40792 11671 40848
rect 11727 40792 11795 40848
rect 11851 40792 11919 40848
rect 11975 40792 12043 40848
rect 12099 40792 12167 40848
rect 12223 40792 12291 40848
rect 12347 40792 12415 40848
rect 12471 40792 12481 40848
rect 10669 40724 12481 40792
rect 10669 40668 10679 40724
rect 10735 40668 10803 40724
rect 10859 40668 10927 40724
rect 10983 40668 11051 40724
rect 11107 40668 11175 40724
rect 11231 40668 11299 40724
rect 11355 40668 11423 40724
rect 11479 40668 11547 40724
rect 11603 40668 11671 40724
rect 11727 40668 11795 40724
rect 11851 40668 11919 40724
rect 11975 40668 12043 40724
rect 12099 40668 12167 40724
rect 12223 40668 12291 40724
rect 12347 40668 12415 40724
rect 12471 40668 12481 40724
rect 10669 40600 12481 40668
rect 10669 40544 10679 40600
rect 10735 40544 10803 40600
rect 10859 40544 10927 40600
rect 10983 40544 11051 40600
rect 11107 40544 11175 40600
rect 11231 40544 11299 40600
rect 11355 40544 11423 40600
rect 11479 40544 11547 40600
rect 11603 40544 11671 40600
rect 11727 40544 11795 40600
rect 11851 40544 11919 40600
rect 11975 40544 12043 40600
rect 12099 40544 12167 40600
rect 12223 40544 12291 40600
rect 12347 40544 12415 40600
rect 12471 40544 12481 40600
rect 10669 40476 12481 40544
rect 10669 40420 10679 40476
rect 10735 40420 10803 40476
rect 10859 40420 10927 40476
rect 10983 40420 11051 40476
rect 11107 40420 11175 40476
rect 11231 40420 11299 40476
rect 11355 40420 11423 40476
rect 11479 40420 11547 40476
rect 11603 40420 11671 40476
rect 11727 40420 11795 40476
rect 11851 40420 11919 40476
rect 11975 40420 12043 40476
rect 12099 40420 12167 40476
rect 12223 40420 12291 40476
rect 12347 40420 12415 40476
rect 12471 40420 12481 40476
rect 10669 40352 12481 40420
rect 10669 40296 10679 40352
rect 10735 40296 10803 40352
rect 10859 40296 10927 40352
rect 10983 40296 11051 40352
rect 11107 40296 11175 40352
rect 11231 40296 11299 40352
rect 11355 40296 11423 40352
rect 11479 40296 11547 40352
rect 11603 40296 11671 40352
rect 11727 40296 11795 40352
rect 11851 40296 11919 40352
rect 11975 40296 12043 40352
rect 12099 40296 12167 40352
rect 12223 40296 12291 40352
rect 12347 40296 12415 40352
rect 12471 40296 12481 40352
rect 10669 40228 12481 40296
rect 10669 40172 10679 40228
rect 10735 40172 10803 40228
rect 10859 40172 10927 40228
rect 10983 40172 11051 40228
rect 11107 40172 11175 40228
rect 11231 40172 11299 40228
rect 11355 40172 11423 40228
rect 11479 40172 11547 40228
rect 11603 40172 11671 40228
rect 11727 40172 11795 40228
rect 11851 40172 11919 40228
rect 11975 40172 12043 40228
rect 12099 40172 12167 40228
rect 12223 40172 12291 40228
rect 12347 40172 12415 40228
rect 12471 40172 12481 40228
rect 10669 40104 12481 40172
rect 10669 40048 10679 40104
rect 10735 40048 10803 40104
rect 10859 40048 10927 40104
rect 10983 40048 11051 40104
rect 11107 40048 11175 40104
rect 11231 40048 11299 40104
rect 11355 40048 11423 40104
rect 11479 40048 11547 40104
rect 11603 40048 11671 40104
rect 11727 40048 11795 40104
rect 11851 40048 11919 40104
rect 11975 40048 12043 40104
rect 12099 40048 12167 40104
rect 12223 40048 12291 40104
rect 12347 40048 12415 40104
rect 12471 40048 12481 40104
rect 10669 40038 12481 40048
rect 6072 39929 6148 39997
rect 6072 39873 6082 39929
rect 6138 39873 6148 39929
rect 6072 39805 6148 39873
rect 6072 39749 6082 39805
rect 6138 39749 6148 39805
rect 6072 39681 6148 39749
rect 6072 39625 6082 39681
rect 6138 39625 6148 39681
rect 6072 39557 6148 39625
rect 6072 39501 6082 39557
rect 6138 39501 6148 39557
rect 6072 39433 6148 39501
rect 6072 39377 6082 39433
rect 6138 39377 6148 39433
rect 6072 39309 6148 39377
rect 6072 39253 6082 39309
rect 6138 39253 6148 39309
rect 6072 39185 6148 39253
rect 6072 39129 6082 39185
rect 6138 39129 6148 39185
rect 6072 39061 6148 39129
rect 6072 39005 6082 39061
rect 6138 39005 6148 39061
rect 6072 38937 6148 39005
rect 6072 38881 6082 38937
rect 6138 38881 6148 38937
rect 6072 38813 6148 38881
rect 6072 38757 6082 38813
rect 6138 38757 6148 38813
rect 6072 38689 6148 38757
rect 6072 38633 6082 38689
rect 6138 38633 6148 38689
rect 6072 38565 6148 38633
rect 6072 38509 6082 38565
rect 6138 38509 6148 38565
rect 6072 38499 6148 38509
rect 7552 39744 8620 39754
rect 7552 39688 7562 39744
rect 7618 39688 7686 39744
rect 7742 39688 7810 39744
rect 7866 39688 7934 39744
rect 7990 39688 8058 39744
rect 8114 39688 8182 39744
rect 8238 39688 8306 39744
rect 8362 39688 8430 39744
rect 8486 39688 8554 39744
rect 8610 39688 8620 39744
rect 7552 39620 8620 39688
rect 7552 39564 7562 39620
rect 7618 39564 7686 39620
rect 7742 39564 7810 39620
rect 7866 39564 7934 39620
rect 7990 39564 8058 39620
rect 8114 39564 8182 39620
rect 8238 39564 8306 39620
rect 8362 39564 8430 39620
rect 8486 39564 8554 39620
rect 8610 39564 8620 39620
rect 7552 39496 8620 39564
rect 7552 39440 7562 39496
rect 7618 39440 7686 39496
rect 7742 39440 7810 39496
rect 7866 39440 7934 39496
rect 7990 39440 8058 39496
rect 8114 39440 8182 39496
rect 8238 39440 8306 39496
rect 8362 39440 8430 39496
rect 8486 39440 8554 39496
rect 8610 39440 8620 39496
rect 7552 39372 8620 39440
rect 7552 39316 7562 39372
rect 7618 39316 7686 39372
rect 7742 39316 7810 39372
rect 7866 39316 7934 39372
rect 7990 39316 8058 39372
rect 8114 39316 8182 39372
rect 8238 39316 8306 39372
rect 8362 39316 8430 39372
rect 8486 39316 8554 39372
rect 8610 39316 8620 39372
rect 7552 39248 8620 39316
rect 7552 39192 7562 39248
rect 7618 39192 7686 39248
rect 7742 39192 7810 39248
rect 7866 39192 7934 39248
rect 7990 39192 8058 39248
rect 8114 39192 8182 39248
rect 8238 39192 8306 39248
rect 8362 39192 8430 39248
rect 8486 39192 8554 39248
rect 8610 39192 8620 39248
rect 7552 39124 8620 39192
rect 7552 39068 7562 39124
rect 7618 39068 7686 39124
rect 7742 39068 7810 39124
rect 7866 39068 7934 39124
rect 7990 39068 8058 39124
rect 8114 39068 8182 39124
rect 8238 39068 8306 39124
rect 8362 39068 8430 39124
rect 8486 39068 8554 39124
rect 8610 39068 8620 39124
rect 7552 39000 8620 39068
rect 7552 38944 7562 39000
rect 7618 38944 7686 39000
rect 7742 38944 7810 39000
rect 7866 38944 7934 39000
rect 7990 38944 8058 39000
rect 8114 38944 8182 39000
rect 8238 38944 8306 39000
rect 8362 38944 8430 39000
rect 8486 38944 8554 39000
rect 8610 38944 8620 39000
rect 7552 38876 8620 38944
rect 7552 38820 7562 38876
rect 7618 38820 7686 38876
rect 7742 38820 7810 38876
rect 7866 38820 7934 38876
rect 7990 38820 8058 38876
rect 8114 38820 8182 38876
rect 8238 38820 8306 38876
rect 8362 38820 8430 38876
rect 8486 38820 8554 38876
rect 8610 38820 8620 38876
rect 7552 38752 8620 38820
rect 7552 38696 7562 38752
rect 7618 38696 7686 38752
rect 7742 38696 7810 38752
rect 7866 38696 7934 38752
rect 7990 38696 8058 38752
rect 8114 38696 8182 38752
rect 8238 38696 8306 38752
rect 8362 38696 8430 38752
rect 8486 38696 8554 38752
rect 8610 38696 8620 38752
rect 7552 38628 8620 38696
rect 7552 38572 7562 38628
rect 7618 38572 7686 38628
rect 7742 38572 7810 38628
rect 7866 38572 7934 38628
rect 7990 38572 8058 38628
rect 8114 38572 8182 38628
rect 8238 38572 8306 38628
rect 8362 38572 8430 38628
rect 8486 38572 8554 38628
rect 8610 38572 8620 38628
rect 7552 38504 8620 38572
rect 7552 38448 7562 38504
rect 7618 38448 7686 38504
rect 7742 38448 7810 38504
rect 7866 38448 7934 38504
rect 7990 38448 8058 38504
rect 8114 38448 8182 38504
rect 8238 38448 8306 38504
rect 8362 38448 8430 38504
rect 8486 38448 8554 38504
rect 8610 38448 8620 38504
rect 7552 38438 8620 38448
rect 10669 39744 12481 39754
rect 10669 39688 10679 39744
rect 10735 39688 10803 39744
rect 10859 39688 10927 39744
rect 10983 39688 11051 39744
rect 11107 39688 11175 39744
rect 11231 39688 11299 39744
rect 11355 39688 11423 39744
rect 11479 39688 11547 39744
rect 11603 39688 11671 39744
rect 11727 39688 11795 39744
rect 11851 39688 11919 39744
rect 11975 39688 12043 39744
rect 12099 39688 12167 39744
rect 12223 39688 12291 39744
rect 12347 39688 12415 39744
rect 12471 39688 12481 39744
rect 10669 39620 12481 39688
rect 10669 39564 10679 39620
rect 10735 39564 10803 39620
rect 10859 39564 10927 39620
rect 10983 39564 11051 39620
rect 11107 39564 11175 39620
rect 11231 39564 11299 39620
rect 11355 39564 11423 39620
rect 11479 39564 11547 39620
rect 11603 39564 11671 39620
rect 11727 39564 11795 39620
rect 11851 39564 11919 39620
rect 11975 39564 12043 39620
rect 12099 39564 12167 39620
rect 12223 39564 12291 39620
rect 12347 39564 12415 39620
rect 12471 39564 12481 39620
rect 10669 39496 12481 39564
rect 10669 39440 10679 39496
rect 10735 39440 10803 39496
rect 10859 39440 10927 39496
rect 10983 39440 11051 39496
rect 11107 39440 11175 39496
rect 11231 39440 11299 39496
rect 11355 39440 11423 39496
rect 11479 39440 11547 39496
rect 11603 39440 11671 39496
rect 11727 39440 11795 39496
rect 11851 39440 11919 39496
rect 11975 39440 12043 39496
rect 12099 39440 12167 39496
rect 12223 39440 12291 39496
rect 12347 39440 12415 39496
rect 12471 39440 12481 39496
rect 10669 39372 12481 39440
rect 10669 39316 10679 39372
rect 10735 39316 10803 39372
rect 10859 39316 10927 39372
rect 10983 39316 11051 39372
rect 11107 39316 11175 39372
rect 11231 39316 11299 39372
rect 11355 39316 11423 39372
rect 11479 39316 11547 39372
rect 11603 39316 11671 39372
rect 11727 39316 11795 39372
rect 11851 39316 11919 39372
rect 11975 39316 12043 39372
rect 12099 39316 12167 39372
rect 12223 39316 12291 39372
rect 12347 39316 12415 39372
rect 12471 39316 12481 39372
rect 10669 39248 12481 39316
rect 10669 39192 10679 39248
rect 10735 39192 10803 39248
rect 10859 39192 10927 39248
rect 10983 39192 11051 39248
rect 11107 39192 11175 39248
rect 11231 39192 11299 39248
rect 11355 39192 11423 39248
rect 11479 39192 11547 39248
rect 11603 39192 11671 39248
rect 11727 39192 11795 39248
rect 11851 39192 11919 39248
rect 11975 39192 12043 39248
rect 12099 39192 12167 39248
rect 12223 39192 12291 39248
rect 12347 39192 12415 39248
rect 12471 39192 12481 39248
rect 10669 39124 12481 39192
rect 10669 39068 10679 39124
rect 10735 39068 10803 39124
rect 10859 39068 10927 39124
rect 10983 39068 11051 39124
rect 11107 39068 11175 39124
rect 11231 39068 11299 39124
rect 11355 39068 11423 39124
rect 11479 39068 11547 39124
rect 11603 39068 11671 39124
rect 11727 39068 11795 39124
rect 11851 39068 11919 39124
rect 11975 39068 12043 39124
rect 12099 39068 12167 39124
rect 12223 39068 12291 39124
rect 12347 39068 12415 39124
rect 12471 39068 12481 39124
rect 10669 39000 12481 39068
rect 10669 38944 10679 39000
rect 10735 38944 10803 39000
rect 10859 38944 10927 39000
rect 10983 38944 11051 39000
rect 11107 38944 11175 39000
rect 11231 38944 11299 39000
rect 11355 38944 11423 39000
rect 11479 38944 11547 39000
rect 11603 38944 11671 39000
rect 11727 38944 11795 39000
rect 11851 38944 11919 39000
rect 11975 38944 12043 39000
rect 12099 38944 12167 39000
rect 12223 38944 12291 39000
rect 12347 38944 12415 39000
rect 12471 38944 12481 39000
rect 10669 38876 12481 38944
rect 10669 38820 10679 38876
rect 10735 38820 10803 38876
rect 10859 38820 10927 38876
rect 10983 38820 11051 38876
rect 11107 38820 11175 38876
rect 11231 38820 11299 38876
rect 11355 38820 11423 38876
rect 11479 38820 11547 38876
rect 11603 38820 11671 38876
rect 11727 38820 11795 38876
rect 11851 38820 11919 38876
rect 11975 38820 12043 38876
rect 12099 38820 12167 38876
rect 12223 38820 12291 38876
rect 12347 38820 12415 38876
rect 12471 38820 12481 38876
rect 10669 38752 12481 38820
rect 10669 38696 10679 38752
rect 10735 38696 10803 38752
rect 10859 38696 10927 38752
rect 10983 38696 11051 38752
rect 11107 38696 11175 38752
rect 11231 38696 11299 38752
rect 11355 38696 11423 38752
rect 11479 38696 11547 38752
rect 11603 38696 11671 38752
rect 11727 38696 11795 38752
rect 11851 38696 11919 38752
rect 11975 38696 12043 38752
rect 12099 38696 12167 38752
rect 12223 38696 12291 38752
rect 12347 38696 12415 38752
rect 12471 38696 12481 38752
rect 10669 38628 12481 38696
rect 10669 38572 10679 38628
rect 10735 38572 10803 38628
rect 10859 38572 10927 38628
rect 10983 38572 11051 38628
rect 11107 38572 11175 38628
rect 11231 38572 11299 38628
rect 11355 38572 11423 38628
rect 11479 38572 11547 38628
rect 11603 38572 11671 38628
rect 11727 38572 11795 38628
rect 11851 38572 11919 38628
rect 11975 38572 12043 38628
rect 12099 38572 12167 38628
rect 12223 38572 12291 38628
rect 12347 38572 12415 38628
rect 12471 38572 12481 38628
rect 10669 38504 12481 38572
rect 10669 38448 10679 38504
rect 10735 38448 10803 38504
rect 10859 38448 10927 38504
rect 10983 38448 11051 38504
rect 11107 38448 11175 38504
rect 11231 38448 11299 38504
rect 11355 38448 11423 38504
rect 11479 38448 11547 38504
rect 11603 38448 11671 38504
rect 11727 38448 11795 38504
rect 11851 38448 11919 38504
rect 11975 38448 12043 38504
rect 12099 38448 12167 38504
rect 12223 38448 12291 38504
rect 12347 38448 12415 38504
rect 12471 38448 12481 38504
rect 10669 38438 12481 38448
rect 2517 37000 2593 37010
rect 2517 36944 2527 37000
rect 2583 36944 2593 37000
rect 2517 36876 2593 36944
rect 2517 36820 2527 36876
rect 2583 36820 2593 36876
rect 2517 36752 2593 36820
rect 2517 36696 2527 36752
rect 2583 36696 2593 36752
rect 2517 36628 2593 36696
rect 2517 36572 2527 36628
rect 2583 36572 2593 36628
rect 2517 36504 2593 36572
rect 2517 36448 2527 36504
rect 2583 36448 2593 36504
rect 2517 36380 2593 36448
rect 2517 36324 2527 36380
rect 2583 36324 2593 36380
rect 2517 36256 2593 36324
rect 2517 36200 2527 36256
rect 2583 36200 2593 36256
rect 2517 36132 2593 36200
rect 2517 36076 2527 36132
rect 2583 36076 2593 36132
rect 2517 36008 2593 36076
rect 2517 35952 2527 36008
rect 2583 35952 2593 36008
rect 2517 35884 2593 35952
rect 2517 35828 2527 35884
rect 2583 35828 2593 35884
rect 2517 35760 2593 35828
rect 2517 35704 2527 35760
rect 2583 35704 2593 35760
rect 2517 35636 2593 35704
rect 2517 35580 2527 35636
rect 2583 35580 2593 35636
rect 2517 35512 2593 35580
rect 2517 35456 2527 35512
rect 2583 35456 2593 35512
rect 2517 35388 2593 35456
rect 2517 35332 2527 35388
rect 2583 35332 2593 35388
rect 2517 35264 2593 35332
rect 2517 35208 2527 35264
rect 2583 35208 2593 35264
rect 2517 35140 2593 35208
rect 2517 35084 2527 35140
rect 2583 35084 2593 35140
rect 2517 35016 2593 35084
rect 2517 34960 2527 35016
rect 2583 34960 2593 35016
rect 2517 34892 2593 34960
rect 2517 34836 2527 34892
rect 2583 34836 2593 34892
rect 2517 34768 2593 34836
rect 2517 34712 2527 34768
rect 2583 34712 2593 34768
rect 2517 34644 2593 34712
rect 2517 34588 2527 34644
rect 2583 34588 2593 34644
rect 2517 34520 2593 34588
rect 2517 34464 2527 34520
rect 2583 34464 2593 34520
rect 2517 34396 2593 34464
rect 2517 34340 2527 34396
rect 2583 34340 2593 34396
rect 2517 34272 2593 34340
rect 2517 34216 2527 34272
rect 2583 34216 2593 34272
rect 2517 34148 2593 34216
rect 2517 34092 2527 34148
rect 2583 34092 2593 34148
rect 2517 34024 2593 34092
rect 2517 33968 2527 34024
rect 2583 33968 2593 34024
rect 2517 33900 2593 33968
rect 2517 33844 2527 33900
rect 2583 33844 2593 33900
rect 2517 33776 2593 33844
rect 1145 33766 1221 33776
rect 1145 33710 1155 33766
rect 1211 33710 1221 33766
rect 1145 33642 1221 33710
rect 2517 33720 2527 33776
rect 2583 33720 2593 33776
rect 2517 33652 2593 33720
rect 1145 33586 1155 33642
rect 1211 33586 1221 33642
rect 1145 33518 1221 33586
rect 1145 33462 1155 33518
rect 1211 33462 1221 33518
rect 1145 33394 1221 33462
rect 1145 33338 1155 33394
rect 1211 33338 1221 33394
rect 1145 33270 1221 33338
rect 1145 33214 1155 33270
rect 1211 33214 1221 33270
rect 1145 33146 1221 33214
rect 1145 33090 1155 33146
rect 1211 33090 1221 33146
rect 1145 33022 1221 33090
rect 1145 32966 1155 33022
rect 1211 32966 1221 33022
rect 1145 32898 1221 32966
rect 1145 32842 1155 32898
rect 1211 32842 1221 32898
rect 1145 32774 1221 32842
rect 1145 32718 1155 32774
rect 1211 32718 1221 32774
rect 1145 32650 1221 32718
rect 1145 32594 1155 32650
rect 1211 32594 1221 32650
rect 1145 32526 1221 32594
rect 1145 32470 1155 32526
rect 1211 32470 1221 32526
rect 1145 32402 1221 32470
rect 1145 32346 1155 32402
rect 1211 32346 1221 32402
rect 1145 32278 1221 32346
rect 1145 32222 1155 32278
rect 1211 32222 1221 32278
rect 1145 32154 1221 32222
rect 1145 32098 1155 32154
rect 1211 32098 1221 32154
rect 1145 32030 1221 32098
rect 1145 31974 1155 32030
rect 1211 31974 1221 32030
rect 1145 31906 1221 31974
rect 1145 31850 1155 31906
rect 1211 31850 1221 31906
rect 1145 31782 1221 31850
rect 1145 31726 1155 31782
rect 1211 31726 1221 31782
rect 1145 31658 1221 31726
rect 1145 31602 1155 31658
rect 1211 31602 1221 31658
rect 1145 31534 1221 31602
rect 1145 31478 1155 31534
rect 1211 31478 1221 31534
rect 1145 31410 1221 31478
rect 1145 31354 1155 31410
rect 1211 31354 1221 31410
rect 1145 31286 1221 31354
rect 1145 31230 1155 31286
rect 1211 31230 1221 31286
rect 1145 31162 1221 31230
rect 1145 31106 1155 31162
rect 1211 31106 1221 31162
rect 1145 31038 1221 31106
rect 1145 30982 1155 31038
rect 1211 30982 1221 31038
rect 1145 30914 1221 30982
rect 1145 30858 1155 30914
rect 1211 30858 1221 30914
rect 1145 30790 1221 30858
rect 1145 30734 1155 30790
rect 1211 30734 1221 30790
rect 1145 30666 1221 30734
rect 1145 30610 1155 30666
rect 1211 30610 1221 30666
rect 1145 30542 1221 30610
rect 1145 30486 1155 30542
rect 1211 30486 1221 30542
rect 1145 30418 1221 30486
rect 1145 30362 1155 30418
rect 1211 30362 1221 30418
rect 1145 30294 1221 30362
rect 1145 30238 1155 30294
rect 1211 30238 1221 30294
rect 1145 30170 1221 30238
rect 1145 30114 1155 30170
rect 1211 30114 1221 30170
rect 1145 30046 1221 30114
rect 1145 29990 1155 30046
rect 1211 29990 1221 30046
rect 1145 29922 1221 29990
rect 1145 29866 1155 29922
rect 1211 29866 1221 29922
rect 1145 29798 1221 29866
rect 1145 29742 1155 29798
rect 1211 29742 1221 29798
rect 1145 29732 1221 29742
rect 1269 33642 1345 33652
rect 1269 33586 1279 33642
rect 1335 33586 1345 33642
rect 1269 33518 1345 33586
rect 2517 33596 2527 33652
rect 2583 33596 2593 33652
rect 2517 33528 2593 33596
rect 1269 33462 1279 33518
rect 1335 33462 1345 33518
rect 1269 33394 1345 33462
rect 1269 33338 1279 33394
rect 1335 33338 1345 33394
rect 1269 33270 1345 33338
rect 1269 33214 1279 33270
rect 1335 33214 1345 33270
rect 1269 33146 1345 33214
rect 1269 33090 1279 33146
rect 1335 33090 1345 33146
rect 1269 33022 1345 33090
rect 1269 32966 1279 33022
rect 1335 32966 1345 33022
rect 1269 32898 1345 32966
rect 1269 32842 1279 32898
rect 1335 32842 1345 32898
rect 1269 32774 1345 32842
rect 1269 32718 1279 32774
rect 1335 32718 1345 32774
rect 1269 32650 1345 32718
rect 1269 32594 1279 32650
rect 1335 32594 1345 32650
rect 1269 32526 1345 32594
rect 1269 32470 1279 32526
rect 1335 32470 1345 32526
rect 1269 32402 1345 32470
rect 1269 32346 1279 32402
rect 1335 32346 1345 32402
rect 1269 32278 1345 32346
rect 1269 32222 1279 32278
rect 1335 32222 1345 32278
rect 1269 32154 1345 32222
rect 1269 32098 1279 32154
rect 1335 32098 1345 32154
rect 1269 32030 1345 32098
rect 1269 31974 1279 32030
rect 1335 31974 1345 32030
rect 1269 31906 1345 31974
rect 1269 31850 1279 31906
rect 1335 31850 1345 31906
rect 1269 31782 1345 31850
rect 1269 31726 1279 31782
rect 1335 31726 1345 31782
rect 1269 31658 1345 31726
rect 1269 31602 1279 31658
rect 1335 31602 1345 31658
rect 1269 31534 1345 31602
rect 1269 31478 1279 31534
rect 1335 31478 1345 31534
rect 1269 31410 1345 31478
rect 1269 31354 1279 31410
rect 1335 31354 1345 31410
rect 1269 31286 1345 31354
rect 1269 31230 1279 31286
rect 1335 31230 1345 31286
rect 1269 31162 1345 31230
rect 1269 31106 1279 31162
rect 1335 31106 1345 31162
rect 1269 31038 1345 31106
rect 1269 30982 1279 31038
rect 1335 30982 1345 31038
rect 1269 30914 1345 30982
rect 1269 30858 1279 30914
rect 1335 30858 1345 30914
rect 1269 30790 1345 30858
rect 1269 30734 1279 30790
rect 1335 30734 1345 30790
rect 1269 30666 1345 30734
rect 1269 30610 1279 30666
rect 1335 30610 1345 30666
rect 1269 30542 1345 30610
rect 1269 30486 1279 30542
rect 1335 30486 1345 30542
rect 1269 30418 1345 30486
rect 1269 30362 1279 30418
rect 1335 30362 1345 30418
rect 1269 30294 1345 30362
rect 1269 30238 1279 30294
rect 1335 30238 1345 30294
rect 1269 30170 1345 30238
rect 1269 30114 1279 30170
rect 1335 30114 1345 30170
rect 1269 30046 1345 30114
rect 1269 29990 1279 30046
rect 1335 29990 1345 30046
rect 1269 29922 1345 29990
rect 1269 29866 1279 29922
rect 1335 29866 1345 29922
rect 1269 29798 1345 29866
rect 1269 29742 1279 29798
rect 1335 29742 1345 29798
rect 1269 29674 1345 29742
rect 1269 29618 1279 29674
rect 1335 29618 1345 29674
rect 1269 29608 1345 29618
rect 1393 33518 1469 33528
rect 1393 33462 1403 33518
rect 1459 33462 1469 33518
rect 1393 33394 1469 33462
rect 2517 33472 2527 33528
rect 2583 33472 2593 33528
rect 2517 33404 2593 33472
rect 1393 33338 1403 33394
rect 1459 33338 1469 33394
rect 1393 33270 1469 33338
rect 1393 33214 1403 33270
rect 1459 33214 1469 33270
rect 1393 33146 1469 33214
rect 1393 33090 1403 33146
rect 1459 33090 1469 33146
rect 1393 33022 1469 33090
rect 1393 32966 1403 33022
rect 1459 32966 1469 33022
rect 1393 32898 1469 32966
rect 1393 32842 1403 32898
rect 1459 32842 1469 32898
rect 1393 32774 1469 32842
rect 1393 32718 1403 32774
rect 1459 32718 1469 32774
rect 1393 32650 1469 32718
rect 1393 32594 1403 32650
rect 1459 32594 1469 32650
rect 1393 32526 1469 32594
rect 1393 32470 1403 32526
rect 1459 32470 1469 32526
rect 1393 32402 1469 32470
rect 1393 32346 1403 32402
rect 1459 32346 1469 32402
rect 1393 32278 1469 32346
rect 1393 32222 1403 32278
rect 1459 32222 1469 32278
rect 1393 32154 1469 32222
rect 1393 32098 1403 32154
rect 1459 32098 1469 32154
rect 1393 32030 1469 32098
rect 1393 31974 1403 32030
rect 1459 31974 1469 32030
rect 1393 31906 1469 31974
rect 1393 31850 1403 31906
rect 1459 31850 1469 31906
rect 1393 31782 1469 31850
rect 1393 31726 1403 31782
rect 1459 31726 1469 31782
rect 1393 31658 1469 31726
rect 1393 31602 1403 31658
rect 1459 31602 1469 31658
rect 1393 31534 1469 31602
rect 1393 31478 1403 31534
rect 1459 31478 1469 31534
rect 1393 31410 1469 31478
rect 1393 31354 1403 31410
rect 1459 31354 1469 31410
rect 1393 31286 1469 31354
rect 1393 31230 1403 31286
rect 1459 31230 1469 31286
rect 1393 31162 1469 31230
rect 1393 31106 1403 31162
rect 1459 31106 1469 31162
rect 1393 31038 1469 31106
rect 1393 30982 1403 31038
rect 1459 30982 1469 31038
rect 1393 30914 1469 30982
rect 1393 30858 1403 30914
rect 1459 30858 1469 30914
rect 1393 30790 1469 30858
rect 1393 30734 1403 30790
rect 1459 30734 1469 30790
rect 1393 30666 1469 30734
rect 1393 30610 1403 30666
rect 1459 30610 1469 30666
rect 1393 30542 1469 30610
rect 1393 30486 1403 30542
rect 1459 30486 1469 30542
rect 1393 30418 1469 30486
rect 1393 30362 1403 30418
rect 1459 30362 1469 30418
rect 1393 30294 1469 30362
rect 1393 30238 1403 30294
rect 1459 30238 1469 30294
rect 1393 30170 1469 30238
rect 1393 30114 1403 30170
rect 1459 30114 1469 30170
rect 1393 30046 1469 30114
rect 1393 29990 1403 30046
rect 1459 29990 1469 30046
rect 1393 29922 1469 29990
rect 1393 29866 1403 29922
rect 1459 29866 1469 29922
rect 1393 29798 1469 29866
rect 1393 29742 1403 29798
rect 1459 29742 1469 29798
rect 1393 29674 1469 29742
rect 1393 29618 1403 29674
rect 1459 29618 1469 29674
rect 1393 29550 1469 29618
rect 1393 29494 1403 29550
rect 1459 29494 1469 29550
rect 1393 29484 1469 29494
rect 1517 33394 1593 33404
rect 1517 33338 1527 33394
rect 1583 33338 1593 33394
rect 1517 33270 1593 33338
rect 2517 33348 2527 33404
rect 2583 33348 2593 33404
rect 2517 33280 2593 33348
rect 1517 33214 1527 33270
rect 1583 33214 1593 33270
rect 1517 33146 1593 33214
rect 1517 33090 1527 33146
rect 1583 33090 1593 33146
rect 1517 33022 1593 33090
rect 1517 32966 1527 33022
rect 1583 32966 1593 33022
rect 1517 32898 1593 32966
rect 1517 32842 1527 32898
rect 1583 32842 1593 32898
rect 1517 32774 1593 32842
rect 1517 32718 1527 32774
rect 1583 32718 1593 32774
rect 1517 32650 1593 32718
rect 1517 32594 1527 32650
rect 1583 32594 1593 32650
rect 1517 32526 1593 32594
rect 1517 32470 1527 32526
rect 1583 32470 1593 32526
rect 1517 32402 1593 32470
rect 1517 32346 1527 32402
rect 1583 32346 1593 32402
rect 1517 32278 1593 32346
rect 1517 32222 1527 32278
rect 1583 32222 1593 32278
rect 1517 32154 1593 32222
rect 1517 32098 1527 32154
rect 1583 32098 1593 32154
rect 1517 32030 1593 32098
rect 1517 31974 1527 32030
rect 1583 31974 1593 32030
rect 1517 31906 1593 31974
rect 1517 31850 1527 31906
rect 1583 31850 1593 31906
rect 1517 31782 1593 31850
rect 1517 31726 1527 31782
rect 1583 31726 1593 31782
rect 1517 31658 1593 31726
rect 1517 31602 1527 31658
rect 1583 31602 1593 31658
rect 1517 31534 1593 31602
rect 1517 31478 1527 31534
rect 1583 31478 1593 31534
rect 1517 31410 1593 31478
rect 1517 31354 1527 31410
rect 1583 31354 1593 31410
rect 1517 31286 1593 31354
rect 1517 31230 1527 31286
rect 1583 31230 1593 31286
rect 1517 31162 1593 31230
rect 1517 31106 1527 31162
rect 1583 31106 1593 31162
rect 1517 31038 1593 31106
rect 1517 30982 1527 31038
rect 1583 30982 1593 31038
rect 1517 30914 1593 30982
rect 1517 30858 1527 30914
rect 1583 30858 1593 30914
rect 1517 30790 1593 30858
rect 1517 30734 1527 30790
rect 1583 30734 1593 30790
rect 1517 30666 1593 30734
rect 1517 30610 1527 30666
rect 1583 30610 1593 30666
rect 1517 30542 1593 30610
rect 1517 30486 1527 30542
rect 1583 30486 1593 30542
rect 1517 30418 1593 30486
rect 1517 30362 1527 30418
rect 1583 30362 1593 30418
rect 1517 30294 1593 30362
rect 1517 30238 1527 30294
rect 1583 30238 1593 30294
rect 1517 30170 1593 30238
rect 1517 30114 1527 30170
rect 1583 30114 1593 30170
rect 1517 30046 1593 30114
rect 1517 29990 1527 30046
rect 1583 29990 1593 30046
rect 1517 29922 1593 29990
rect 1517 29866 1527 29922
rect 1583 29866 1593 29922
rect 1517 29798 1593 29866
rect 1517 29742 1527 29798
rect 1583 29742 1593 29798
rect 1517 29674 1593 29742
rect 1517 29618 1527 29674
rect 1583 29618 1593 29674
rect 1517 29550 1593 29618
rect 1517 29494 1527 29550
rect 1583 29494 1593 29550
rect 1517 29426 1593 29494
rect 1517 29370 1527 29426
rect 1583 29370 1593 29426
rect 1517 29360 1593 29370
rect 1641 33270 1717 33280
rect 1641 33214 1651 33270
rect 1707 33214 1717 33270
rect 1641 33146 1717 33214
rect 2517 33224 2527 33280
rect 2583 33224 2593 33280
rect 2517 33156 2593 33224
rect 1641 33090 1651 33146
rect 1707 33090 1717 33146
rect 1641 33022 1717 33090
rect 1641 32966 1651 33022
rect 1707 32966 1717 33022
rect 1641 32898 1717 32966
rect 1641 32842 1651 32898
rect 1707 32842 1717 32898
rect 1641 32774 1717 32842
rect 1641 32718 1651 32774
rect 1707 32718 1717 32774
rect 1641 32650 1717 32718
rect 1641 32594 1651 32650
rect 1707 32594 1717 32650
rect 1641 32526 1717 32594
rect 1641 32470 1651 32526
rect 1707 32470 1717 32526
rect 1641 32402 1717 32470
rect 1641 32346 1651 32402
rect 1707 32346 1717 32402
rect 1641 32278 1717 32346
rect 1641 32222 1651 32278
rect 1707 32222 1717 32278
rect 1641 32154 1717 32222
rect 1641 32098 1651 32154
rect 1707 32098 1717 32154
rect 1641 32030 1717 32098
rect 1641 31974 1651 32030
rect 1707 31974 1717 32030
rect 1641 31906 1717 31974
rect 1641 31850 1651 31906
rect 1707 31850 1717 31906
rect 1641 31782 1717 31850
rect 1641 31726 1651 31782
rect 1707 31726 1717 31782
rect 1641 31658 1717 31726
rect 1641 31602 1651 31658
rect 1707 31602 1717 31658
rect 1641 31534 1717 31602
rect 1641 31478 1651 31534
rect 1707 31478 1717 31534
rect 1641 31410 1717 31478
rect 1641 31354 1651 31410
rect 1707 31354 1717 31410
rect 1641 31286 1717 31354
rect 1641 31230 1651 31286
rect 1707 31230 1717 31286
rect 1641 31162 1717 31230
rect 1641 31106 1651 31162
rect 1707 31106 1717 31162
rect 1641 31038 1717 31106
rect 1641 30982 1651 31038
rect 1707 30982 1717 31038
rect 1641 30914 1717 30982
rect 1641 30858 1651 30914
rect 1707 30858 1717 30914
rect 1641 30790 1717 30858
rect 1641 30734 1651 30790
rect 1707 30734 1717 30790
rect 1641 30666 1717 30734
rect 1641 30610 1651 30666
rect 1707 30610 1717 30666
rect 1641 30542 1717 30610
rect 1641 30486 1651 30542
rect 1707 30486 1717 30542
rect 1641 30418 1717 30486
rect 1641 30362 1651 30418
rect 1707 30362 1717 30418
rect 1641 30294 1717 30362
rect 1641 30238 1651 30294
rect 1707 30238 1717 30294
rect 1641 30170 1717 30238
rect 1641 30114 1651 30170
rect 1707 30114 1717 30170
rect 1641 30046 1717 30114
rect 1641 29990 1651 30046
rect 1707 29990 1717 30046
rect 1641 29922 1717 29990
rect 1641 29866 1651 29922
rect 1707 29866 1717 29922
rect 1641 29798 1717 29866
rect 1641 29742 1651 29798
rect 1707 29742 1717 29798
rect 1641 29674 1717 29742
rect 1641 29618 1651 29674
rect 1707 29618 1717 29674
rect 1641 29550 1717 29618
rect 1641 29494 1651 29550
rect 1707 29494 1717 29550
rect 1641 29426 1717 29494
rect 1641 29370 1651 29426
rect 1707 29370 1717 29426
rect 1117 29307 1193 29317
rect 1117 29251 1127 29307
rect 1183 29251 1193 29307
rect 1117 29183 1193 29251
rect 1641 29302 1717 29370
rect 1641 29246 1651 29302
rect 1707 29246 1717 29302
rect 1641 29236 1717 29246
rect 1765 33146 1841 33156
rect 1765 33090 1775 33146
rect 1831 33090 1841 33146
rect 1765 33022 1841 33090
rect 2517 33100 2527 33156
rect 2583 33100 2593 33156
rect 2517 33032 2593 33100
rect 1765 32966 1775 33022
rect 1831 32966 1841 33022
rect 1765 32898 1841 32966
rect 1765 32842 1775 32898
rect 1831 32842 1841 32898
rect 1765 32774 1841 32842
rect 1765 32718 1775 32774
rect 1831 32718 1841 32774
rect 1765 32650 1841 32718
rect 1765 32594 1775 32650
rect 1831 32594 1841 32650
rect 1765 32526 1841 32594
rect 1765 32470 1775 32526
rect 1831 32470 1841 32526
rect 1765 32402 1841 32470
rect 1765 32346 1775 32402
rect 1831 32346 1841 32402
rect 1765 32278 1841 32346
rect 1765 32222 1775 32278
rect 1831 32222 1841 32278
rect 1765 32154 1841 32222
rect 1765 32098 1775 32154
rect 1831 32098 1841 32154
rect 1765 32030 1841 32098
rect 1765 31974 1775 32030
rect 1831 31974 1841 32030
rect 1765 31906 1841 31974
rect 1765 31850 1775 31906
rect 1831 31850 1841 31906
rect 1765 31782 1841 31850
rect 1765 31726 1775 31782
rect 1831 31726 1841 31782
rect 1765 31658 1841 31726
rect 1765 31602 1775 31658
rect 1831 31602 1841 31658
rect 1765 31534 1841 31602
rect 1765 31478 1775 31534
rect 1831 31478 1841 31534
rect 1765 31410 1841 31478
rect 1765 31354 1775 31410
rect 1831 31354 1841 31410
rect 1765 31286 1841 31354
rect 1765 31230 1775 31286
rect 1831 31230 1841 31286
rect 1765 31162 1841 31230
rect 1765 31106 1775 31162
rect 1831 31106 1841 31162
rect 1765 31038 1841 31106
rect 1765 30982 1775 31038
rect 1831 30982 1841 31038
rect 1765 30914 1841 30982
rect 1765 30858 1775 30914
rect 1831 30858 1841 30914
rect 1765 30790 1841 30858
rect 1765 30734 1775 30790
rect 1831 30734 1841 30790
rect 1765 30666 1841 30734
rect 1765 30610 1775 30666
rect 1831 30610 1841 30666
rect 1765 30542 1841 30610
rect 1765 30486 1775 30542
rect 1831 30486 1841 30542
rect 1765 30418 1841 30486
rect 1765 30362 1775 30418
rect 1831 30362 1841 30418
rect 1765 30294 1841 30362
rect 1765 30238 1775 30294
rect 1831 30238 1841 30294
rect 1765 30170 1841 30238
rect 1765 30114 1775 30170
rect 1831 30114 1841 30170
rect 1765 30046 1841 30114
rect 1765 29990 1775 30046
rect 1831 29990 1841 30046
rect 1765 29922 1841 29990
rect 1765 29866 1775 29922
rect 1831 29866 1841 29922
rect 1765 29798 1841 29866
rect 1765 29742 1775 29798
rect 1831 29742 1841 29798
rect 1765 29674 1841 29742
rect 1765 29618 1775 29674
rect 1831 29618 1841 29674
rect 1765 29550 1841 29618
rect 1765 29494 1775 29550
rect 1831 29494 1841 29550
rect 1765 29426 1841 29494
rect 1765 29370 1775 29426
rect 1831 29370 1841 29426
rect 1765 29302 1841 29370
rect 1765 29246 1775 29302
rect 1831 29246 1841 29302
rect 1117 29127 1127 29183
rect 1183 29127 1193 29183
rect 1117 29059 1193 29127
rect 1117 29003 1127 29059
rect 1183 29003 1193 29059
rect 1117 28935 1193 29003
rect 1117 28879 1127 28935
rect 1183 28879 1193 28935
rect 1117 28811 1193 28879
rect 1117 28755 1127 28811
rect 1183 28755 1193 28811
rect 1117 28687 1193 28755
rect 1117 28631 1127 28687
rect 1183 28631 1193 28687
rect 1117 28563 1193 28631
rect 1117 28507 1127 28563
rect 1183 28507 1193 28563
rect 1117 28439 1193 28507
rect 1117 28383 1127 28439
rect 1183 28383 1193 28439
rect 1117 28315 1193 28383
rect 1117 28259 1127 28315
rect 1183 28259 1193 28315
rect 1117 28191 1193 28259
rect 1117 28135 1127 28191
rect 1183 28135 1193 28191
rect 1117 28067 1193 28135
rect 1117 28011 1127 28067
rect 1183 28011 1193 28067
rect 1117 27943 1193 28011
rect 1117 27887 1127 27943
rect 1183 27887 1193 27943
rect 1117 27819 1193 27887
rect 1117 27763 1127 27819
rect 1183 27763 1193 27819
rect 1117 27695 1193 27763
rect 1117 27639 1127 27695
rect 1183 27639 1193 27695
rect 1117 27571 1193 27639
rect 1117 27515 1127 27571
rect 1183 27515 1193 27571
rect 1117 27505 1193 27515
rect 1241 29183 1317 29193
rect 1241 29127 1251 29183
rect 1307 29127 1317 29183
rect 1241 29059 1317 29127
rect 1765 29178 1841 29246
rect 1765 29122 1775 29178
rect 1831 29122 1841 29178
rect 1765 29112 1841 29122
rect 1889 33022 1965 33032
rect 1889 32966 1899 33022
rect 1955 32966 1965 33022
rect 2517 32976 2527 33032
rect 2583 32976 2593 33032
rect 2517 32966 2593 32976
rect 2641 36876 2717 36886
rect 2641 36820 2651 36876
rect 2707 36820 2717 36876
rect 2641 36752 2717 36820
rect 2641 36696 2651 36752
rect 2707 36696 2717 36752
rect 2641 36628 2717 36696
rect 2641 36572 2651 36628
rect 2707 36572 2717 36628
rect 2641 36504 2717 36572
rect 2641 36448 2651 36504
rect 2707 36448 2717 36504
rect 2641 36380 2717 36448
rect 2641 36324 2651 36380
rect 2707 36324 2717 36380
rect 2641 36256 2717 36324
rect 2641 36200 2651 36256
rect 2707 36200 2717 36256
rect 2641 36132 2717 36200
rect 2641 36076 2651 36132
rect 2707 36076 2717 36132
rect 2641 36008 2717 36076
rect 2641 35952 2651 36008
rect 2707 35952 2717 36008
rect 2641 35884 2717 35952
rect 2641 35828 2651 35884
rect 2707 35828 2717 35884
rect 2641 35760 2717 35828
rect 2641 35704 2651 35760
rect 2707 35704 2717 35760
rect 2641 35636 2717 35704
rect 2641 35580 2651 35636
rect 2707 35580 2717 35636
rect 2641 35512 2717 35580
rect 2641 35456 2651 35512
rect 2707 35456 2717 35512
rect 2641 35388 2717 35456
rect 2641 35332 2651 35388
rect 2707 35332 2717 35388
rect 2641 35264 2717 35332
rect 2641 35208 2651 35264
rect 2707 35208 2717 35264
rect 2641 35140 2717 35208
rect 2641 35084 2651 35140
rect 2707 35084 2717 35140
rect 2641 35016 2717 35084
rect 2641 34960 2651 35016
rect 2707 34960 2717 35016
rect 2641 34892 2717 34960
rect 2641 34836 2651 34892
rect 2707 34836 2717 34892
rect 2641 34768 2717 34836
rect 2641 34712 2651 34768
rect 2707 34712 2717 34768
rect 2641 34644 2717 34712
rect 2641 34588 2651 34644
rect 2707 34588 2717 34644
rect 2641 34520 2717 34588
rect 2641 34464 2651 34520
rect 2707 34464 2717 34520
rect 2641 34396 2717 34464
rect 2641 34340 2651 34396
rect 2707 34340 2717 34396
rect 2641 34272 2717 34340
rect 2641 34216 2651 34272
rect 2707 34216 2717 34272
rect 2641 34148 2717 34216
rect 2641 34092 2651 34148
rect 2707 34092 2717 34148
rect 2641 34024 2717 34092
rect 2641 33968 2651 34024
rect 2707 33968 2717 34024
rect 2641 33900 2717 33968
rect 2641 33844 2651 33900
rect 2707 33844 2717 33900
rect 2641 33776 2717 33844
rect 2641 33720 2651 33776
rect 2707 33720 2717 33776
rect 2641 33652 2717 33720
rect 2641 33596 2651 33652
rect 2707 33596 2717 33652
rect 2641 33528 2717 33596
rect 2641 33472 2651 33528
rect 2707 33472 2717 33528
rect 2641 33404 2717 33472
rect 2641 33348 2651 33404
rect 2707 33348 2717 33404
rect 2641 33280 2717 33348
rect 2641 33224 2651 33280
rect 2707 33224 2717 33280
rect 2641 33156 2717 33224
rect 2641 33100 2651 33156
rect 2707 33100 2717 33156
rect 2641 33032 2717 33100
rect 2641 32976 2651 33032
rect 2707 32976 2717 33032
rect 1889 32898 1965 32966
rect 2641 32908 2717 32976
rect 1889 32842 1899 32898
rect 1955 32842 1965 32898
rect 1889 32774 1965 32842
rect 1889 32718 1899 32774
rect 1955 32718 1965 32774
rect 1889 32650 1965 32718
rect 1889 32594 1899 32650
rect 1955 32594 1965 32650
rect 1889 32526 1965 32594
rect 1889 32470 1899 32526
rect 1955 32470 1965 32526
rect 1889 32402 1965 32470
rect 1889 32346 1899 32402
rect 1955 32346 1965 32402
rect 1889 32278 1965 32346
rect 1889 32222 1899 32278
rect 1955 32222 1965 32278
rect 1889 32154 1965 32222
rect 1889 32098 1899 32154
rect 1955 32098 1965 32154
rect 1889 32030 1965 32098
rect 1889 31974 1899 32030
rect 1955 31974 1965 32030
rect 1889 31906 1965 31974
rect 1889 31850 1899 31906
rect 1955 31850 1965 31906
rect 1889 31782 1965 31850
rect 1889 31726 1899 31782
rect 1955 31726 1965 31782
rect 1889 31658 1965 31726
rect 1889 31602 1899 31658
rect 1955 31602 1965 31658
rect 1889 31534 1965 31602
rect 1889 31478 1899 31534
rect 1955 31478 1965 31534
rect 1889 31410 1965 31478
rect 1889 31354 1899 31410
rect 1955 31354 1965 31410
rect 1889 31286 1965 31354
rect 1889 31230 1899 31286
rect 1955 31230 1965 31286
rect 1889 31162 1965 31230
rect 1889 31106 1899 31162
rect 1955 31106 1965 31162
rect 1889 31038 1965 31106
rect 1889 30982 1899 31038
rect 1955 30982 1965 31038
rect 1889 30914 1965 30982
rect 1889 30858 1899 30914
rect 1955 30858 1965 30914
rect 1889 30790 1965 30858
rect 1889 30734 1899 30790
rect 1955 30734 1965 30790
rect 1889 30666 1965 30734
rect 1889 30610 1899 30666
rect 1955 30610 1965 30666
rect 1889 30542 1965 30610
rect 1889 30486 1899 30542
rect 1955 30486 1965 30542
rect 1889 30418 1965 30486
rect 1889 30362 1899 30418
rect 1955 30362 1965 30418
rect 1889 30294 1965 30362
rect 1889 30238 1899 30294
rect 1955 30238 1965 30294
rect 1889 30170 1965 30238
rect 1889 30114 1899 30170
rect 1955 30114 1965 30170
rect 1889 30046 1965 30114
rect 1889 29990 1899 30046
rect 1955 29990 1965 30046
rect 1889 29922 1965 29990
rect 1889 29866 1899 29922
rect 1955 29866 1965 29922
rect 1889 29798 1965 29866
rect 1889 29742 1899 29798
rect 1955 29742 1965 29798
rect 1889 29674 1965 29742
rect 1889 29618 1899 29674
rect 1955 29618 1965 29674
rect 1889 29550 1965 29618
rect 1889 29494 1899 29550
rect 1955 29494 1965 29550
rect 1889 29426 1965 29494
rect 1889 29370 1899 29426
rect 1955 29370 1965 29426
rect 1889 29302 1965 29370
rect 1889 29246 1899 29302
rect 1955 29246 1965 29302
rect 1889 29178 1965 29246
rect 1889 29122 1899 29178
rect 1955 29122 1965 29178
rect 1241 29003 1251 29059
rect 1307 29003 1317 29059
rect 1241 28935 1317 29003
rect 1241 28879 1251 28935
rect 1307 28879 1317 28935
rect 1241 28811 1317 28879
rect 1241 28755 1251 28811
rect 1307 28755 1317 28811
rect 1241 28687 1317 28755
rect 1241 28631 1251 28687
rect 1307 28631 1317 28687
rect 1241 28563 1317 28631
rect 1241 28507 1251 28563
rect 1307 28507 1317 28563
rect 1241 28439 1317 28507
rect 1241 28383 1251 28439
rect 1307 28383 1317 28439
rect 1241 28315 1317 28383
rect 1241 28259 1251 28315
rect 1307 28259 1317 28315
rect 1241 28191 1317 28259
rect 1241 28135 1251 28191
rect 1307 28135 1317 28191
rect 1241 28067 1317 28135
rect 1241 28011 1251 28067
rect 1307 28011 1317 28067
rect 1241 27943 1317 28011
rect 1241 27887 1251 27943
rect 1307 27887 1317 27943
rect 1241 27819 1317 27887
rect 1241 27763 1251 27819
rect 1307 27763 1317 27819
rect 1241 27695 1317 27763
rect 1241 27639 1251 27695
rect 1307 27639 1317 27695
rect 1241 27571 1317 27639
rect 1241 27515 1251 27571
rect 1307 27515 1317 27571
rect 1241 27447 1317 27515
rect 1241 27391 1251 27447
rect 1307 27391 1317 27447
rect 1241 27381 1317 27391
rect 1365 29059 1441 29069
rect 1365 29003 1375 29059
rect 1431 29003 1441 29059
rect 1365 28935 1441 29003
rect 1889 29054 1965 29122
rect 1889 28998 1899 29054
rect 1955 28998 1965 29054
rect 1889 28988 1965 28998
rect 2013 32898 2089 32908
rect 2013 32842 2023 32898
rect 2079 32842 2089 32898
rect 2641 32852 2651 32908
rect 2707 32852 2717 32908
rect 2641 32842 2717 32852
rect 2765 36752 2841 36762
rect 2765 36696 2775 36752
rect 2831 36696 2841 36752
rect 2765 36628 2841 36696
rect 2765 36572 2775 36628
rect 2831 36572 2841 36628
rect 2765 36504 2841 36572
rect 2765 36448 2775 36504
rect 2831 36448 2841 36504
rect 2765 36380 2841 36448
rect 2765 36324 2775 36380
rect 2831 36324 2841 36380
rect 2765 36256 2841 36324
rect 2765 36200 2775 36256
rect 2831 36200 2841 36256
rect 2765 36132 2841 36200
rect 2765 36076 2775 36132
rect 2831 36076 2841 36132
rect 2765 36008 2841 36076
rect 2765 35952 2775 36008
rect 2831 35952 2841 36008
rect 2765 35884 2841 35952
rect 2765 35828 2775 35884
rect 2831 35828 2841 35884
rect 2765 35760 2841 35828
rect 2765 35704 2775 35760
rect 2831 35704 2841 35760
rect 2765 35636 2841 35704
rect 2765 35580 2775 35636
rect 2831 35580 2841 35636
rect 2765 35512 2841 35580
rect 2765 35456 2775 35512
rect 2831 35456 2841 35512
rect 2765 35388 2841 35456
rect 2765 35332 2775 35388
rect 2831 35332 2841 35388
rect 2765 35264 2841 35332
rect 2765 35208 2775 35264
rect 2831 35208 2841 35264
rect 2765 35140 2841 35208
rect 2765 35084 2775 35140
rect 2831 35084 2841 35140
rect 2765 35016 2841 35084
rect 2765 34960 2775 35016
rect 2831 34960 2841 35016
rect 2765 34892 2841 34960
rect 2765 34836 2775 34892
rect 2831 34836 2841 34892
rect 2765 34768 2841 34836
rect 2765 34712 2775 34768
rect 2831 34712 2841 34768
rect 2765 34644 2841 34712
rect 2765 34588 2775 34644
rect 2831 34588 2841 34644
rect 2765 34520 2841 34588
rect 2765 34464 2775 34520
rect 2831 34464 2841 34520
rect 2765 34396 2841 34464
rect 2765 34340 2775 34396
rect 2831 34340 2841 34396
rect 2765 34272 2841 34340
rect 2765 34216 2775 34272
rect 2831 34216 2841 34272
rect 2765 34148 2841 34216
rect 2765 34092 2775 34148
rect 2831 34092 2841 34148
rect 2765 34024 2841 34092
rect 2765 33968 2775 34024
rect 2831 33968 2841 34024
rect 2765 33900 2841 33968
rect 2765 33844 2775 33900
rect 2831 33844 2841 33900
rect 2765 33776 2841 33844
rect 2765 33720 2775 33776
rect 2831 33720 2841 33776
rect 2765 33652 2841 33720
rect 2765 33596 2775 33652
rect 2831 33596 2841 33652
rect 2765 33528 2841 33596
rect 2765 33472 2775 33528
rect 2831 33472 2841 33528
rect 2765 33404 2841 33472
rect 2765 33348 2775 33404
rect 2831 33348 2841 33404
rect 2765 33280 2841 33348
rect 2765 33224 2775 33280
rect 2831 33224 2841 33280
rect 2765 33156 2841 33224
rect 2765 33100 2775 33156
rect 2831 33100 2841 33156
rect 2765 33032 2841 33100
rect 2765 32976 2775 33032
rect 2831 32976 2841 33032
rect 2765 32908 2841 32976
rect 2765 32852 2775 32908
rect 2831 32852 2841 32908
rect 2013 32774 2089 32842
rect 2013 32718 2023 32774
rect 2079 32718 2089 32774
rect 2765 32784 2841 32852
rect 2765 32728 2775 32784
rect 2831 32728 2841 32784
rect 2765 32718 2841 32728
rect 2889 36628 2965 36638
rect 2889 36572 2899 36628
rect 2955 36572 2965 36628
rect 2889 36504 2965 36572
rect 14757 36572 14833 36582
rect 2889 36448 2899 36504
rect 2955 36448 2965 36504
rect 2889 36380 2965 36448
rect 2889 36324 2899 36380
rect 2955 36324 2965 36380
rect 2889 36256 2965 36324
rect 2889 36200 2899 36256
rect 2955 36200 2965 36256
rect 2889 36132 2965 36200
rect 2889 36076 2899 36132
rect 2955 36076 2965 36132
rect 2889 36008 2965 36076
rect 2889 35952 2899 36008
rect 2955 35952 2965 36008
rect 2889 35884 2965 35952
rect 2889 35828 2899 35884
rect 2955 35828 2965 35884
rect 2889 35760 2965 35828
rect 2889 35704 2899 35760
rect 2955 35704 2965 35760
rect 2889 35636 2965 35704
rect 2889 35580 2899 35636
rect 2955 35580 2965 35636
rect 2889 35512 2965 35580
rect 2889 35456 2899 35512
rect 2955 35456 2965 35512
rect 2889 35388 2965 35456
rect 2889 35332 2899 35388
rect 2955 35332 2965 35388
rect 2889 35264 2965 35332
rect 2889 35208 2899 35264
rect 2955 35208 2965 35264
rect 2889 35140 2965 35208
rect 2889 35084 2899 35140
rect 2955 35084 2965 35140
rect 2889 35016 2965 35084
rect 2889 34960 2899 35016
rect 2955 34960 2965 35016
rect 2889 34892 2965 34960
rect 2889 34836 2899 34892
rect 2955 34836 2965 34892
rect 2889 34768 2965 34836
rect 2889 34712 2899 34768
rect 2955 34712 2965 34768
rect 2889 34644 2965 34712
rect 2889 34588 2899 34644
rect 2955 34588 2965 34644
rect 2889 34520 2965 34588
rect 2889 34464 2899 34520
rect 2955 34464 2965 34520
rect 2889 34396 2965 34464
rect 2889 34340 2899 34396
rect 2955 34340 2965 34396
rect 2889 34272 2965 34340
rect 2889 34216 2899 34272
rect 2955 34216 2965 34272
rect 2889 34148 2965 34216
rect 2889 34092 2899 34148
rect 2955 34092 2965 34148
rect 2889 34024 2965 34092
rect 2889 33968 2899 34024
rect 2955 33968 2965 34024
rect 2889 33900 2965 33968
rect 2889 33844 2899 33900
rect 2955 33844 2965 33900
rect 2889 33776 2965 33844
rect 2889 33720 2899 33776
rect 2955 33720 2965 33776
rect 2889 33652 2965 33720
rect 2889 33596 2899 33652
rect 2955 33596 2965 33652
rect 2889 33528 2965 33596
rect 2889 33472 2899 33528
rect 2955 33472 2965 33528
rect 2889 33404 2965 33472
rect 2889 33348 2899 33404
rect 2955 33348 2965 33404
rect 2889 33280 2965 33348
rect 2889 33224 2899 33280
rect 2955 33224 2965 33280
rect 2889 33156 2965 33224
rect 2889 33100 2899 33156
rect 2955 33100 2965 33156
rect 2889 33032 2965 33100
rect 2889 32976 2899 33032
rect 2955 32976 2965 33032
rect 2889 32908 2965 32976
rect 2889 32852 2899 32908
rect 2955 32852 2965 32908
rect 2889 32784 2965 32852
rect 2889 32728 2899 32784
rect 2955 32728 2965 32784
rect 2013 32650 2089 32718
rect 2013 32594 2023 32650
rect 2079 32594 2089 32650
rect 2889 32660 2965 32728
rect 2889 32604 2899 32660
rect 2955 32604 2965 32660
rect 2889 32594 2965 32604
rect 3013 36504 3089 36514
rect 3013 36448 3023 36504
rect 3079 36448 3089 36504
rect 3013 36380 3089 36448
rect 3013 36324 3023 36380
rect 3079 36324 3089 36380
rect 3013 36256 3089 36324
rect 3013 36200 3023 36256
rect 3079 36200 3089 36256
rect 3013 36132 3089 36200
rect 3013 36076 3023 36132
rect 3079 36076 3089 36132
rect 3013 36008 3089 36076
rect 3013 35952 3023 36008
rect 3079 35952 3089 36008
rect 3013 35884 3089 35952
rect 3013 35828 3023 35884
rect 3079 35828 3089 35884
rect 3013 35760 3089 35828
rect 3013 35704 3023 35760
rect 3079 35704 3089 35760
rect 3013 35636 3089 35704
rect 3013 35580 3023 35636
rect 3079 35580 3089 35636
rect 3013 35512 3089 35580
rect 3013 35456 3023 35512
rect 3079 35456 3089 35512
rect 3013 35388 3089 35456
rect 3013 35332 3023 35388
rect 3079 35332 3089 35388
rect 3013 35264 3089 35332
rect 3013 35208 3023 35264
rect 3079 35208 3089 35264
rect 3013 35140 3089 35208
rect 3013 35084 3023 35140
rect 3079 35084 3089 35140
rect 3013 35016 3089 35084
rect 3013 34960 3023 35016
rect 3079 34960 3089 35016
rect 3013 34892 3089 34960
rect 3013 34836 3023 34892
rect 3079 34836 3089 34892
rect 3013 34768 3089 34836
rect 3013 34712 3023 34768
rect 3079 34712 3089 34768
rect 3013 34644 3089 34712
rect 3013 34588 3023 34644
rect 3079 34588 3089 34644
rect 3013 34520 3089 34588
rect 3013 34464 3023 34520
rect 3079 34464 3089 34520
rect 3013 34396 3089 34464
rect 3013 34340 3023 34396
rect 3079 34340 3089 34396
rect 3013 34272 3089 34340
rect 3013 34216 3023 34272
rect 3079 34216 3089 34272
rect 3013 34148 3089 34216
rect 3013 34092 3023 34148
rect 3079 34092 3089 34148
rect 3013 34024 3089 34092
rect 3013 33968 3023 34024
rect 3079 33968 3089 34024
rect 3013 33900 3089 33968
rect 3013 33844 3023 33900
rect 3079 33844 3089 33900
rect 3013 33776 3089 33844
rect 3013 33720 3023 33776
rect 3079 33720 3089 33776
rect 3013 33652 3089 33720
rect 3013 33596 3023 33652
rect 3079 33596 3089 33652
rect 3013 33528 3089 33596
rect 3013 33472 3023 33528
rect 3079 33472 3089 33528
rect 3013 33404 3089 33472
rect 3013 33348 3023 33404
rect 3079 33348 3089 33404
rect 3013 33280 3089 33348
rect 3013 33224 3023 33280
rect 3079 33224 3089 33280
rect 3013 33156 3089 33224
rect 3013 33100 3023 33156
rect 3079 33100 3089 33156
rect 3013 33032 3089 33100
rect 3013 32976 3023 33032
rect 3079 32976 3089 33032
rect 3013 32908 3089 32976
rect 3013 32852 3023 32908
rect 3079 32852 3089 32908
rect 3013 32784 3089 32852
rect 3013 32728 3023 32784
rect 3079 32728 3089 32784
rect 3013 32660 3089 32728
rect 3013 32604 3023 32660
rect 3079 32604 3089 32660
rect 2013 32526 2089 32594
rect 2013 32470 2023 32526
rect 2079 32470 2089 32526
rect 3013 32536 3089 32604
rect 3013 32480 3023 32536
rect 3079 32480 3089 32536
rect 3013 32470 3089 32480
rect 3137 36380 3213 36390
rect 3137 36324 3147 36380
rect 3203 36324 3213 36380
rect 3137 36256 3213 36324
rect 3137 36200 3147 36256
rect 3203 36200 3213 36256
rect 3137 36132 3213 36200
rect 3137 36076 3147 36132
rect 3203 36076 3213 36132
rect 3137 36008 3213 36076
rect 3137 35952 3147 36008
rect 3203 35952 3213 36008
rect 3137 35884 3213 35952
rect 3137 35828 3147 35884
rect 3203 35828 3213 35884
rect 3137 35760 3213 35828
rect 3137 35704 3147 35760
rect 3203 35704 3213 35760
rect 3137 35636 3213 35704
rect 3137 35580 3147 35636
rect 3203 35580 3213 35636
rect 3137 35512 3213 35580
rect 3137 35456 3147 35512
rect 3203 35456 3213 35512
rect 3137 35388 3213 35456
rect 3137 35332 3147 35388
rect 3203 35332 3213 35388
rect 3137 35264 3213 35332
rect 3137 35208 3147 35264
rect 3203 35208 3213 35264
rect 3137 35140 3213 35208
rect 3137 35084 3147 35140
rect 3203 35084 3213 35140
rect 3137 35016 3213 35084
rect 3137 34960 3147 35016
rect 3203 34960 3213 35016
rect 3137 34892 3213 34960
rect 3137 34836 3147 34892
rect 3203 34836 3213 34892
rect 3137 34768 3213 34836
rect 3137 34712 3147 34768
rect 3203 34712 3213 34768
rect 3137 34644 3213 34712
rect 3137 34588 3147 34644
rect 3203 34588 3213 34644
rect 3137 34520 3213 34588
rect 3137 34464 3147 34520
rect 3203 34464 3213 34520
rect 3137 34396 3213 34464
rect 3137 34340 3147 34396
rect 3203 34340 3213 34396
rect 3137 34272 3213 34340
rect 3137 34216 3147 34272
rect 3203 34216 3213 34272
rect 3137 34148 3213 34216
rect 3137 34092 3147 34148
rect 3203 34092 3213 34148
rect 3137 34024 3213 34092
rect 3137 33968 3147 34024
rect 3203 33968 3213 34024
rect 3137 33900 3213 33968
rect 3137 33844 3147 33900
rect 3203 33844 3213 33900
rect 3137 33776 3213 33844
rect 3137 33720 3147 33776
rect 3203 33720 3213 33776
rect 3137 33652 3213 33720
rect 3137 33596 3147 33652
rect 3203 33596 3213 33652
rect 3137 33528 3213 33596
rect 3137 33472 3147 33528
rect 3203 33472 3213 33528
rect 3137 33404 3213 33472
rect 3137 33348 3147 33404
rect 3203 33348 3213 33404
rect 3137 33280 3213 33348
rect 3137 33224 3147 33280
rect 3203 33224 3213 33280
rect 3137 33156 3213 33224
rect 3137 33100 3147 33156
rect 3203 33100 3213 33156
rect 3137 33032 3213 33100
rect 3137 32976 3147 33032
rect 3203 32976 3213 33032
rect 3137 32908 3213 32976
rect 3137 32852 3147 32908
rect 3203 32852 3213 32908
rect 3137 32784 3213 32852
rect 3137 32728 3147 32784
rect 3203 32728 3213 32784
rect 3137 32660 3213 32728
rect 3137 32604 3147 32660
rect 3203 32604 3213 32660
rect 3137 32536 3213 32604
rect 3137 32480 3147 32536
rect 3203 32480 3213 32536
rect 2013 32402 2089 32470
rect 2013 32346 2023 32402
rect 2079 32346 2089 32402
rect 3137 32412 3213 32480
rect 3137 32356 3147 32412
rect 3203 32356 3213 32412
rect 3137 32346 3213 32356
rect 3261 36256 3337 36266
rect 3261 36200 3271 36256
rect 3327 36200 3337 36256
rect 3261 36132 3337 36200
rect 3261 36076 3271 36132
rect 3327 36076 3337 36132
rect 3261 36008 3337 36076
rect 3261 35952 3271 36008
rect 3327 35952 3337 36008
rect 3261 35884 3337 35952
rect 3261 35828 3271 35884
rect 3327 35828 3337 35884
rect 3261 35760 3337 35828
rect 3261 35704 3271 35760
rect 3327 35704 3337 35760
rect 3261 35636 3337 35704
rect 3261 35580 3271 35636
rect 3327 35580 3337 35636
rect 3261 35512 3337 35580
rect 3261 35456 3271 35512
rect 3327 35456 3337 35512
rect 3261 35388 3337 35456
rect 3261 35332 3271 35388
rect 3327 35332 3337 35388
rect 3261 35264 3337 35332
rect 3261 35208 3271 35264
rect 3327 35208 3337 35264
rect 3261 35140 3337 35208
rect 3261 35084 3271 35140
rect 3327 35084 3337 35140
rect 3261 35016 3337 35084
rect 3261 34960 3271 35016
rect 3327 34960 3337 35016
rect 3261 34892 3337 34960
rect 3261 34836 3271 34892
rect 3327 34836 3337 34892
rect 3261 34768 3337 34836
rect 3261 34712 3271 34768
rect 3327 34712 3337 34768
rect 3261 34644 3337 34712
rect 3261 34588 3271 34644
rect 3327 34588 3337 34644
rect 3261 34520 3337 34588
rect 3261 34464 3271 34520
rect 3327 34464 3337 34520
rect 3261 34396 3337 34464
rect 3261 34340 3271 34396
rect 3327 34340 3337 34396
rect 3261 34272 3337 34340
rect 3261 34216 3271 34272
rect 3327 34216 3337 34272
rect 3261 34148 3337 34216
rect 3261 34092 3271 34148
rect 3327 34092 3337 34148
rect 3261 34024 3337 34092
rect 3261 33968 3271 34024
rect 3327 33968 3337 34024
rect 3261 33900 3337 33968
rect 3261 33844 3271 33900
rect 3327 33844 3337 33900
rect 3261 33776 3337 33844
rect 3261 33720 3271 33776
rect 3327 33720 3337 33776
rect 3261 33652 3337 33720
rect 3261 33596 3271 33652
rect 3327 33596 3337 33652
rect 3261 33528 3337 33596
rect 3261 33472 3271 33528
rect 3327 33472 3337 33528
rect 3261 33404 3337 33472
rect 3261 33348 3271 33404
rect 3327 33348 3337 33404
rect 3261 33280 3337 33348
rect 3261 33224 3271 33280
rect 3327 33224 3337 33280
rect 3261 33156 3337 33224
rect 3261 33100 3271 33156
rect 3327 33100 3337 33156
rect 3261 33032 3337 33100
rect 3261 32976 3271 33032
rect 3327 32976 3337 33032
rect 3261 32908 3337 32976
rect 3261 32852 3271 32908
rect 3327 32852 3337 32908
rect 3261 32784 3337 32852
rect 3261 32728 3271 32784
rect 3327 32728 3337 32784
rect 3261 32660 3337 32728
rect 3261 32604 3271 32660
rect 3327 32604 3337 32660
rect 3261 32536 3337 32604
rect 3261 32480 3271 32536
rect 3327 32480 3337 32536
rect 3261 32412 3337 32480
rect 3261 32356 3271 32412
rect 3327 32356 3337 32412
rect 2013 32278 2089 32346
rect 2013 32222 2023 32278
rect 2079 32222 2089 32278
rect 3261 32288 3337 32356
rect 3261 32232 3271 32288
rect 3327 32232 3337 32288
rect 3261 32222 3337 32232
rect 3385 36132 3461 36142
rect 3385 36076 3395 36132
rect 3451 36076 3461 36132
rect 3385 36008 3461 36076
rect 3385 35952 3395 36008
rect 3451 35952 3461 36008
rect 3385 35884 3461 35952
rect 3385 35828 3395 35884
rect 3451 35828 3461 35884
rect 3385 35760 3461 35828
rect 3385 35704 3395 35760
rect 3451 35704 3461 35760
rect 3385 35636 3461 35704
rect 3385 35580 3395 35636
rect 3451 35580 3461 35636
rect 3385 35512 3461 35580
rect 3385 35456 3395 35512
rect 3451 35456 3461 35512
rect 3385 35388 3461 35456
rect 3385 35332 3395 35388
rect 3451 35332 3461 35388
rect 3385 35264 3461 35332
rect 3385 35208 3395 35264
rect 3451 35208 3461 35264
rect 3385 35140 3461 35208
rect 3385 35084 3395 35140
rect 3451 35084 3461 35140
rect 3385 35016 3461 35084
rect 3385 34960 3395 35016
rect 3451 34960 3461 35016
rect 3385 34892 3461 34960
rect 3385 34836 3395 34892
rect 3451 34836 3461 34892
rect 3385 34768 3461 34836
rect 3385 34712 3395 34768
rect 3451 34712 3461 34768
rect 3385 34644 3461 34712
rect 3385 34588 3395 34644
rect 3451 34588 3461 34644
rect 3385 34520 3461 34588
rect 3385 34464 3395 34520
rect 3451 34464 3461 34520
rect 3385 34396 3461 34464
rect 3385 34340 3395 34396
rect 3451 34340 3461 34396
rect 3385 34272 3461 34340
rect 3385 34216 3395 34272
rect 3451 34216 3461 34272
rect 3385 34148 3461 34216
rect 3385 34092 3395 34148
rect 3451 34092 3461 34148
rect 3385 34024 3461 34092
rect 3385 33968 3395 34024
rect 3451 33968 3461 34024
rect 3385 33900 3461 33968
rect 3385 33844 3395 33900
rect 3451 33844 3461 33900
rect 3385 33776 3461 33844
rect 3385 33720 3395 33776
rect 3451 33720 3461 33776
rect 3385 33652 3461 33720
rect 3385 33596 3395 33652
rect 3451 33596 3461 33652
rect 3385 33528 3461 33596
rect 3385 33472 3395 33528
rect 3451 33472 3461 33528
rect 3385 33404 3461 33472
rect 3385 33348 3395 33404
rect 3451 33348 3461 33404
rect 3385 33280 3461 33348
rect 3385 33224 3395 33280
rect 3451 33224 3461 33280
rect 3385 33156 3461 33224
rect 3385 33100 3395 33156
rect 3451 33100 3461 33156
rect 3385 33032 3461 33100
rect 3385 32976 3395 33032
rect 3451 32976 3461 33032
rect 3385 32908 3461 32976
rect 3385 32852 3395 32908
rect 3451 32852 3461 32908
rect 3385 32784 3461 32852
rect 3385 32728 3395 32784
rect 3451 32728 3461 32784
rect 3385 32660 3461 32728
rect 3385 32604 3395 32660
rect 3451 32604 3461 32660
rect 3385 32536 3461 32604
rect 3385 32480 3395 32536
rect 3451 32480 3461 32536
rect 3385 32412 3461 32480
rect 3385 32356 3395 32412
rect 3451 32356 3461 32412
rect 3385 32288 3461 32356
rect 3385 32232 3395 32288
rect 3451 32232 3461 32288
rect 2013 32154 2089 32222
rect 2013 32098 2023 32154
rect 2079 32098 2089 32154
rect 3385 32164 3461 32232
rect 3385 32108 3395 32164
rect 3451 32108 3461 32164
rect 3385 32098 3461 32108
rect 3509 35946 3585 35956
rect 3509 35890 3519 35946
rect 3575 35890 3585 35946
rect 3509 35822 3585 35890
rect 3509 35766 3519 35822
rect 3575 35766 3585 35822
rect 3509 35698 3585 35766
rect 3509 35642 3519 35698
rect 3575 35642 3585 35698
rect 3509 35574 3585 35642
rect 3509 35518 3519 35574
rect 3575 35518 3585 35574
rect 3509 35450 3585 35518
rect 3509 35394 3519 35450
rect 3575 35394 3585 35450
rect 3509 35326 3585 35394
rect 3509 35270 3519 35326
rect 3575 35270 3585 35326
rect 3509 35202 3585 35270
rect 3509 35146 3519 35202
rect 3575 35146 3585 35202
rect 3509 35078 3585 35146
rect 3509 35022 3519 35078
rect 3575 35022 3585 35078
rect 3509 34954 3585 35022
rect 3509 34898 3519 34954
rect 3575 34898 3585 34954
rect 3509 34830 3585 34898
rect 3509 34774 3519 34830
rect 3575 34774 3585 34830
rect 3509 34706 3585 34774
rect 3509 34650 3519 34706
rect 3575 34650 3585 34706
rect 3509 34582 3585 34650
rect 3509 34526 3519 34582
rect 3575 34526 3585 34582
rect 3509 34458 3585 34526
rect 3509 34402 3519 34458
rect 3575 34402 3585 34458
rect 3509 34334 3585 34402
rect 3509 34278 3519 34334
rect 3575 34278 3585 34334
rect 3509 34210 3585 34278
rect 3509 34154 3519 34210
rect 3575 34154 3585 34210
rect 3509 34086 3585 34154
rect 3509 34030 3519 34086
rect 3575 34030 3585 34086
rect 3509 33962 3585 34030
rect 3509 33906 3519 33962
rect 3575 33906 3585 33962
rect 3509 33838 3585 33906
rect 3509 33782 3519 33838
rect 3575 33782 3585 33838
rect 3509 33714 3585 33782
rect 3509 33658 3519 33714
rect 3575 33658 3585 33714
rect 3509 33590 3585 33658
rect 3509 33534 3519 33590
rect 3575 33534 3585 33590
rect 3509 33466 3585 33534
rect 3509 33410 3519 33466
rect 3575 33410 3585 33466
rect 3509 33342 3585 33410
rect 3509 33286 3519 33342
rect 3575 33286 3585 33342
rect 3509 33218 3585 33286
rect 3509 33162 3519 33218
rect 3575 33162 3585 33218
rect 3509 33094 3585 33162
rect 3509 33038 3519 33094
rect 3575 33038 3585 33094
rect 3509 32970 3585 33038
rect 3509 32914 3519 32970
rect 3575 32914 3585 32970
rect 3509 32846 3585 32914
rect 3509 32790 3519 32846
rect 3575 32790 3585 32846
rect 3509 32722 3585 32790
rect 3509 32666 3519 32722
rect 3575 32666 3585 32722
rect 3509 32598 3585 32666
rect 3509 32542 3519 32598
rect 3575 32542 3585 32598
rect 3509 32474 3585 32542
rect 3509 32418 3519 32474
rect 3575 32418 3585 32474
rect 3509 32350 3585 32418
rect 3509 32294 3519 32350
rect 3575 32294 3585 32350
rect 3509 32226 3585 32294
rect 3509 32170 3519 32226
rect 3575 32170 3585 32226
rect 3509 32102 3585 32170
rect 2013 32030 2089 32098
rect 3509 32046 3519 32102
rect 3575 32046 3585 32102
rect 3509 32036 3585 32046
rect 3633 35813 3709 35823
rect 3633 35757 3643 35813
rect 3699 35757 3709 35813
rect 3633 35689 3709 35757
rect 3633 35633 3643 35689
rect 3699 35633 3709 35689
rect 3633 35565 3709 35633
rect 3633 35509 3643 35565
rect 3699 35509 3709 35565
rect 3633 35441 3709 35509
rect 3633 35385 3643 35441
rect 3699 35385 3709 35441
rect 3633 35317 3709 35385
rect 3633 35261 3643 35317
rect 3699 35261 3709 35317
rect 3633 35193 3709 35261
rect 3633 35137 3643 35193
rect 3699 35137 3709 35193
rect 3633 35069 3709 35137
rect 3633 35013 3643 35069
rect 3699 35013 3709 35069
rect 3633 34945 3709 35013
rect 3633 34889 3643 34945
rect 3699 34889 3709 34945
rect 3633 34821 3709 34889
rect 3633 34765 3643 34821
rect 3699 34765 3709 34821
rect 3633 34697 3709 34765
rect 3633 34641 3643 34697
rect 3699 34641 3709 34697
rect 3633 34573 3709 34641
rect 3633 34517 3643 34573
rect 3699 34517 3709 34573
rect 3633 34449 3709 34517
rect 3633 34393 3643 34449
rect 3699 34393 3709 34449
rect 3633 34325 3709 34393
rect 3633 34269 3643 34325
rect 3699 34269 3709 34325
rect 3633 34201 3709 34269
rect 3633 34145 3643 34201
rect 3699 34145 3709 34201
rect 3633 34077 3709 34145
rect 3633 34021 3643 34077
rect 3699 34021 3709 34077
rect 3633 33953 3709 34021
rect 3633 33897 3643 33953
rect 3699 33897 3709 33953
rect 3633 33829 3709 33897
rect 3633 33773 3643 33829
rect 3699 33773 3709 33829
rect 3633 33705 3709 33773
rect 3633 33649 3643 33705
rect 3699 33649 3709 33705
rect 3633 33581 3709 33649
rect 3633 33525 3643 33581
rect 3699 33525 3709 33581
rect 3633 33457 3709 33525
rect 3633 33401 3643 33457
rect 3699 33401 3709 33457
rect 3633 33333 3709 33401
rect 3633 33277 3643 33333
rect 3699 33277 3709 33333
rect 3633 33209 3709 33277
rect 3633 33153 3643 33209
rect 3699 33153 3709 33209
rect 3633 33085 3709 33153
rect 3633 33029 3643 33085
rect 3699 33029 3709 33085
rect 3633 32961 3709 33029
rect 3633 32905 3643 32961
rect 3699 32905 3709 32961
rect 3633 32837 3709 32905
rect 3633 32781 3643 32837
rect 3699 32781 3709 32837
rect 3633 32713 3709 32781
rect 3633 32657 3643 32713
rect 3699 32657 3709 32713
rect 3633 32589 3709 32657
rect 3633 32533 3643 32589
rect 3699 32533 3709 32589
rect 3633 32465 3709 32533
rect 3633 32409 3643 32465
rect 3699 32409 3709 32465
rect 3633 32341 3709 32409
rect 3633 32285 3643 32341
rect 3699 32285 3709 32341
rect 3633 32217 3709 32285
rect 3633 32161 3643 32217
rect 3699 32161 3709 32217
rect 3633 32093 3709 32161
rect 3633 32037 3643 32093
rect 3699 32037 3709 32093
rect 3757 35710 3833 35720
rect 3757 35654 3767 35710
rect 3823 35654 3833 35710
rect 3757 35586 3833 35654
rect 3757 35530 3767 35586
rect 3823 35530 3833 35586
rect 3757 35462 3833 35530
rect 3757 35406 3767 35462
rect 3823 35406 3833 35462
rect 3757 35338 3833 35406
rect 3757 35282 3767 35338
rect 3823 35282 3833 35338
rect 3757 35214 3833 35282
rect 3757 35158 3767 35214
rect 3823 35158 3833 35214
rect 3757 35090 3833 35158
rect 3757 35034 3767 35090
rect 3823 35034 3833 35090
rect 3757 34966 3833 35034
rect 3757 34910 3767 34966
rect 3823 34910 3833 34966
rect 3757 34842 3833 34910
rect 3757 34786 3767 34842
rect 3823 34786 3833 34842
rect 3757 34718 3833 34786
rect 3757 34662 3767 34718
rect 3823 34662 3833 34718
rect 3757 34594 3833 34662
rect 3757 34538 3767 34594
rect 3823 34538 3833 34594
rect 3757 34470 3833 34538
rect 3757 34414 3767 34470
rect 3823 34414 3833 34470
rect 3757 34346 3833 34414
rect 3757 34290 3767 34346
rect 3823 34290 3833 34346
rect 3757 34222 3833 34290
rect 3757 34166 3767 34222
rect 3823 34166 3833 34222
rect 3757 34098 3833 34166
rect 3757 34042 3767 34098
rect 3823 34042 3833 34098
rect 3757 33974 3833 34042
rect 3757 33918 3767 33974
rect 3823 33918 3833 33974
rect 3757 33850 3833 33918
rect 3757 33794 3767 33850
rect 3823 33794 3833 33850
rect 3757 33726 3833 33794
rect 3757 33670 3767 33726
rect 3823 33670 3833 33726
rect 3757 33602 3833 33670
rect 3757 33546 3767 33602
rect 3823 33546 3833 33602
rect 3757 33478 3833 33546
rect 3757 33422 3767 33478
rect 3823 33422 3833 33478
rect 3757 33354 3833 33422
rect 3757 33298 3767 33354
rect 3823 33298 3833 33354
rect 3757 33230 3833 33298
rect 3757 33174 3767 33230
rect 3823 33174 3833 33230
rect 3757 33106 3833 33174
rect 3757 33050 3767 33106
rect 3823 33050 3833 33106
rect 3757 32982 3833 33050
rect 3757 32926 3767 32982
rect 3823 32926 3833 32982
rect 3757 32858 3833 32926
rect 3757 32802 3767 32858
rect 3823 32802 3833 32858
rect 3757 32734 3833 32802
rect 3757 32678 3767 32734
rect 3823 32678 3833 32734
rect 3757 32610 3833 32678
rect 3757 32554 3767 32610
rect 3823 32554 3833 32610
rect 3757 32486 3833 32554
rect 3757 32430 3767 32486
rect 3823 32430 3833 32486
rect 3757 32362 3833 32430
rect 3757 32306 3767 32362
rect 3823 32306 3833 32362
rect 3757 32238 3833 32306
rect 3757 32182 3767 32238
rect 3823 32182 3833 32238
rect 3757 32114 3833 32182
rect 3757 32058 3767 32114
rect 3823 32058 3833 32114
rect 3881 35606 3957 35616
rect 3881 35550 3891 35606
rect 3947 35550 3957 35606
rect 3881 35482 3957 35550
rect 3881 35426 3891 35482
rect 3947 35426 3957 35482
rect 3881 35358 3957 35426
rect 3881 35302 3891 35358
rect 3947 35302 3957 35358
rect 3881 35234 3957 35302
rect 3881 35178 3891 35234
rect 3947 35178 3957 35234
rect 3881 35110 3957 35178
rect 3881 35054 3891 35110
rect 3947 35054 3957 35110
rect 3881 34986 3957 35054
rect 3881 34930 3891 34986
rect 3947 34930 3957 34986
rect 3881 34862 3957 34930
rect 3881 34806 3891 34862
rect 3947 34806 3957 34862
rect 3881 34738 3957 34806
rect 3881 34682 3891 34738
rect 3947 34682 3957 34738
rect 3881 34614 3957 34682
rect 3881 34558 3891 34614
rect 3947 34558 3957 34614
rect 3881 34490 3957 34558
rect 3881 34434 3891 34490
rect 3947 34434 3957 34490
rect 3881 34366 3957 34434
rect 3881 34310 3891 34366
rect 3947 34310 3957 34366
rect 3881 34242 3957 34310
rect 3881 34186 3891 34242
rect 3947 34186 3957 34242
rect 3881 34118 3957 34186
rect 3881 34062 3891 34118
rect 3947 34062 3957 34118
rect 3881 33994 3957 34062
rect 3881 33938 3891 33994
rect 3947 33938 3957 33994
rect 3881 33870 3957 33938
rect 3881 33814 3891 33870
rect 3947 33814 3957 33870
rect 3881 33746 3957 33814
rect 3881 33690 3891 33746
rect 3947 33690 3957 33746
rect 3881 33622 3957 33690
rect 3881 33566 3891 33622
rect 3947 33566 3957 33622
rect 3881 33498 3957 33566
rect 3881 33442 3891 33498
rect 3947 33442 3957 33498
rect 3881 33374 3957 33442
rect 3881 33318 3891 33374
rect 3947 33318 3957 33374
rect 3881 33250 3957 33318
rect 3881 33194 3891 33250
rect 3947 33194 3957 33250
rect 3881 33126 3957 33194
rect 3881 33070 3891 33126
rect 3947 33070 3957 33126
rect 3881 33002 3957 33070
rect 3881 32946 3891 33002
rect 3947 32946 3957 33002
rect 3881 32878 3957 32946
rect 3881 32822 3891 32878
rect 3947 32822 3957 32878
rect 3881 32754 3957 32822
rect 3881 32698 3891 32754
rect 3947 32698 3957 32754
rect 3881 32630 3957 32698
rect 3881 32574 3891 32630
rect 3947 32574 3957 32630
rect 3881 32506 3957 32574
rect 3881 32450 3891 32506
rect 3947 32450 3957 32506
rect 3881 32382 3957 32450
rect 3881 32326 3891 32382
rect 3947 32326 3957 32382
rect 3881 32258 3957 32326
rect 3881 32202 3891 32258
rect 3947 32202 3957 32258
rect 3881 32134 3957 32202
rect 3881 32078 3891 32134
rect 3947 32078 3957 32134
rect 3881 32068 3957 32078
rect 4005 35535 4081 35545
rect 4005 35479 4015 35535
rect 4071 35479 4081 35535
rect 4005 35411 4081 35479
rect 4005 35355 4015 35411
rect 4071 35355 4081 35411
rect 4005 35287 4081 35355
rect 4005 35231 4015 35287
rect 4071 35231 4081 35287
rect 4005 35163 4081 35231
rect 4005 35107 4015 35163
rect 4071 35107 4081 35163
rect 4005 35039 4081 35107
rect 4005 34983 4015 35039
rect 4071 34983 4081 35039
rect 4005 34915 4081 34983
rect 4005 34859 4015 34915
rect 4071 34859 4081 34915
rect 4005 34791 4081 34859
rect 4005 34735 4015 34791
rect 4071 34735 4081 34791
rect 4005 34667 4081 34735
rect 4005 34611 4015 34667
rect 4071 34611 4081 34667
rect 4005 34543 4081 34611
rect 4005 34487 4015 34543
rect 4071 34487 4081 34543
rect 4005 34419 4081 34487
rect 4005 34363 4015 34419
rect 4071 34363 4081 34419
rect 4005 34295 4081 34363
rect 4005 34239 4015 34295
rect 4071 34239 4081 34295
rect 4005 34171 4081 34239
rect 4005 34115 4015 34171
rect 4071 34115 4081 34171
rect 4005 34047 4081 34115
rect 4005 33991 4015 34047
rect 4071 33991 4081 34047
rect 4005 33923 4081 33991
rect 4005 33867 4015 33923
rect 4071 33867 4081 33923
rect 4005 33799 4081 33867
rect 4005 33743 4015 33799
rect 4071 33743 4081 33799
rect 4005 33675 4081 33743
rect 4005 33619 4015 33675
rect 4071 33619 4081 33675
rect 4005 33551 4081 33619
rect 4005 33495 4015 33551
rect 4071 33495 4081 33551
rect 4005 33427 4081 33495
rect 4005 33371 4015 33427
rect 4071 33371 4081 33427
rect 4005 33303 4081 33371
rect 4005 33247 4015 33303
rect 4071 33247 4081 33303
rect 4005 33179 4081 33247
rect 4005 33123 4015 33179
rect 4071 33123 4081 33179
rect 4005 33055 4081 33123
rect 4005 32999 4015 33055
rect 4071 32999 4081 33055
rect 4005 32931 4081 32999
rect 4005 32875 4015 32931
rect 4071 32875 4081 32931
rect 4005 32807 4081 32875
rect 4005 32751 4015 32807
rect 4071 32751 4081 32807
rect 4005 32683 4081 32751
rect 4005 32627 4015 32683
rect 4071 32627 4081 32683
rect 4005 32559 4081 32627
rect 4005 32503 4015 32559
rect 4071 32503 4081 32559
rect 4005 32435 4081 32503
rect 4005 32379 4015 32435
rect 4071 32379 4081 32435
rect 4005 32311 4081 32379
rect 4005 32255 4015 32311
rect 4071 32255 4081 32311
rect 4005 32187 4081 32255
rect 4005 32131 4015 32187
rect 4071 32131 4081 32187
rect 3757 32048 3833 32058
rect 4005 32063 4081 32131
rect 2013 31974 2023 32030
rect 2079 31974 2089 32030
rect 3633 32027 3709 32037
rect 4005 32007 4015 32063
rect 4071 32007 4081 32063
rect 4005 31997 4081 32007
rect 4129 35417 4205 35427
rect 4129 35361 4139 35417
rect 4195 35361 4205 35417
rect 4129 35293 4205 35361
rect 4129 35237 4139 35293
rect 4195 35237 4205 35293
rect 4129 35169 4205 35237
rect 14757 35220 14767 36572
rect 14823 35220 14833 36572
rect 14757 35210 14833 35220
rect 4129 35113 4139 35169
rect 4195 35113 4205 35169
rect 4129 35045 4205 35113
rect 4129 34989 4139 35045
rect 4195 34989 4205 35045
rect 4129 34921 4205 34989
rect 4129 34865 4139 34921
rect 4195 34865 4205 34921
rect 4129 34797 4205 34865
rect 4129 34741 4139 34797
rect 4195 34741 4205 34797
rect 4129 34673 4205 34741
rect 4129 34617 4139 34673
rect 4195 34617 4205 34673
rect 4129 34549 4205 34617
rect 4129 34493 4139 34549
rect 4195 34493 4205 34549
rect 4129 34425 4205 34493
rect 4129 34369 4139 34425
rect 4195 34369 4205 34425
rect 4129 34301 4205 34369
rect 4129 34245 4139 34301
rect 4195 34245 4205 34301
rect 4129 34177 4205 34245
rect 4129 34121 4139 34177
rect 4195 34121 4205 34177
rect 4129 34053 4205 34121
rect 4129 33997 4139 34053
rect 4195 33997 4205 34053
rect 4129 33929 4205 33997
rect 4129 33873 4139 33929
rect 4195 33873 4205 33929
rect 4129 33805 4205 33873
rect 4129 33749 4139 33805
rect 4195 33749 4205 33805
rect 4129 33681 4205 33749
rect 4129 33625 4139 33681
rect 4195 33625 4205 33681
rect 4129 33557 4205 33625
rect 4129 33501 4139 33557
rect 4195 33501 4205 33557
rect 4129 33433 4205 33501
rect 4129 33377 4139 33433
rect 4195 33377 4205 33433
rect 4129 33309 4205 33377
rect 4129 33253 4139 33309
rect 4195 33253 4205 33309
rect 4129 33185 4205 33253
rect 4129 33129 4139 33185
rect 4195 33129 4205 33185
rect 4129 33061 4205 33129
rect 4129 33005 4139 33061
rect 4195 33005 4205 33061
rect 4129 32937 4205 33005
rect 4129 32881 4139 32937
rect 4195 32881 4205 32937
rect 4129 32813 4205 32881
rect 4129 32757 4139 32813
rect 4195 32757 4205 32813
rect 4129 32689 4205 32757
rect 4129 32633 4139 32689
rect 4195 32633 4205 32689
rect 4129 32565 4205 32633
rect 4129 32509 4139 32565
rect 4195 32509 4205 32565
rect 4129 32441 4205 32509
rect 4129 32385 4139 32441
rect 4195 32385 4205 32441
rect 4129 32317 4205 32385
rect 4129 32261 4139 32317
rect 4195 32261 4205 32317
rect 4129 32193 4205 32261
rect 4129 32137 4139 32193
rect 4195 32137 4205 32193
rect 4129 32069 4205 32137
rect 4129 32013 4139 32069
rect 4195 32013 4205 32069
rect 6358 34950 7426 34960
rect 6358 34894 6368 34950
rect 6424 34894 6492 34950
rect 6548 34894 6616 34950
rect 6672 34894 6740 34950
rect 6796 34894 6864 34950
rect 6920 34894 6988 34950
rect 7044 34894 7112 34950
rect 7168 34894 7236 34950
rect 7292 34894 7360 34950
rect 7416 34894 7426 34950
rect 6358 34826 7426 34894
rect 6358 34770 6368 34826
rect 6424 34770 6492 34826
rect 6548 34770 6616 34826
rect 6672 34770 6740 34826
rect 6796 34770 6864 34826
rect 6920 34770 6988 34826
rect 7044 34770 7112 34826
rect 7168 34770 7236 34826
rect 7292 34770 7360 34826
rect 7416 34770 7426 34826
rect 6358 34702 7426 34770
rect 6358 34646 6368 34702
rect 6424 34646 6492 34702
rect 6548 34646 6616 34702
rect 6672 34646 6740 34702
rect 6796 34646 6864 34702
rect 6920 34646 6988 34702
rect 7044 34646 7112 34702
rect 7168 34646 7236 34702
rect 7292 34646 7360 34702
rect 7416 34646 7426 34702
rect 6358 34578 7426 34646
rect 6358 34522 6368 34578
rect 6424 34522 6492 34578
rect 6548 34522 6616 34578
rect 6672 34522 6740 34578
rect 6796 34522 6864 34578
rect 6920 34522 6988 34578
rect 7044 34522 7112 34578
rect 7168 34522 7236 34578
rect 7292 34522 7360 34578
rect 7416 34522 7426 34578
rect 6358 34454 7426 34522
rect 6358 34398 6368 34454
rect 6424 34398 6492 34454
rect 6548 34398 6616 34454
rect 6672 34398 6740 34454
rect 6796 34398 6864 34454
rect 6920 34398 6988 34454
rect 7044 34398 7112 34454
rect 7168 34398 7236 34454
rect 7292 34398 7360 34454
rect 7416 34398 7426 34454
rect 6358 34330 7426 34398
rect 6358 34274 6368 34330
rect 6424 34274 6492 34330
rect 6548 34274 6616 34330
rect 6672 34274 6740 34330
rect 6796 34274 6864 34330
rect 6920 34274 6988 34330
rect 7044 34274 7112 34330
rect 7168 34274 7236 34330
rect 7292 34274 7360 34330
rect 7416 34274 7426 34330
rect 6358 34206 7426 34274
rect 6358 34150 6368 34206
rect 6424 34150 6492 34206
rect 6548 34150 6616 34206
rect 6672 34150 6740 34206
rect 6796 34150 6864 34206
rect 6920 34150 6988 34206
rect 7044 34150 7112 34206
rect 7168 34150 7236 34206
rect 7292 34150 7360 34206
rect 7416 34150 7426 34206
rect 6358 34082 7426 34150
rect 6358 34026 6368 34082
rect 6424 34026 6492 34082
rect 6548 34026 6616 34082
rect 6672 34026 6740 34082
rect 6796 34026 6864 34082
rect 6920 34026 6988 34082
rect 7044 34026 7112 34082
rect 7168 34026 7236 34082
rect 7292 34026 7360 34082
rect 7416 34026 7426 34082
rect 6358 33958 7426 34026
rect 6358 33902 6368 33958
rect 6424 33902 6492 33958
rect 6548 33902 6616 33958
rect 6672 33902 6740 33958
rect 6796 33902 6864 33958
rect 6920 33902 6988 33958
rect 7044 33902 7112 33958
rect 7168 33902 7236 33958
rect 7292 33902 7360 33958
rect 7416 33902 7426 33958
rect 6358 33834 7426 33902
rect 6358 33778 6368 33834
rect 6424 33778 6492 33834
rect 6548 33778 6616 33834
rect 6672 33778 6740 33834
rect 6796 33778 6864 33834
rect 6920 33778 6988 33834
rect 7044 33778 7112 33834
rect 7168 33778 7236 33834
rect 7292 33778 7360 33834
rect 7416 33778 7426 33834
rect 6358 33710 7426 33778
rect 6358 33654 6368 33710
rect 6424 33654 6492 33710
rect 6548 33654 6616 33710
rect 6672 33654 6740 33710
rect 6796 33654 6864 33710
rect 6920 33654 6988 33710
rect 7044 33654 7112 33710
rect 7168 33654 7236 33710
rect 7292 33654 7360 33710
rect 7416 33654 7426 33710
rect 6358 33586 7426 33654
rect 6358 33530 6368 33586
rect 6424 33530 6492 33586
rect 6548 33530 6616 33586
rect 6672 33530 6740 33586
rect 6796 33530 6864 33586
rect 6920 33530 6988 33586
rect 7044 33530 7112 33586
rect 7168 33530 7236 33586
rect 7292 33530 7360 33586
rect 7416 33530 7426 33586
rect 6358 33462 7426 33530
rect 6358 33406 6368 33462
rect 6424 33406 6492 33462
rect 6548 33406 6616 33462
rect 6672 33406 6740 33462
rect 6796 33406 6864 33462
rect 6920 33406 6988 33462
rect 7044 33406 7112 33462
rect 7168 33406 7236 33462
rect 7292 33406 7360 33462
rect 7416 33406 7426 33462
rect 6358 33338 7426 33406
rect 6358 33282 6368 33338
rect 6424 33282 6492 33338
rect 6548 33282 6616 33338
rect 6672 33282 6740 33338
rect 6796 33282 6864 33338
rect 6920 33282 6988 33338
rect 7044 33282 7112 33338
rect 7168 33282 7236 33338
rect 7292 33282 7360 33338
rect 7416 33282 7426 33338
rect 6358 33214 7426 33282
rect 6358 33158 6368 33214
rect 6424 33158 6492 33214
rect 6548 33158 6616 33214
rect 6672 33158 6740 33214
rect 6796 33158 6864 33214
rect 6920 33158 6988 33214
rect 7044 33158 7112 33214
rect 7168 33158 7236 33214
rect 7292 33158 7360 33214
rect 7416 33158 7426 33214
rect 6358 33090 7426 33158
rect 6358 33034 6368 33090
rect 6424 33034 6492 33090
rect 6548 33034 6616 33090
rect 6672 33034 6740 33090
rect 6796 33034 6864 33090
rect 6920 33034 6988 33090
rect 7044 33034 7112 33090
rect 7168 33034 7236 33090
rect 7292 33034 7360 33090
rect 7416 33034 7426 33090
rect 6358 32966 7426 33034
rect 6358 32910 6368 32966
rect 6424 32910 6492 32966
rect 6548 32910 6616 32966
rect 6672 32910 6740 32966
rect 6796 32910 6864 32966
rect 6920 32910 6988 32966
rect 7044 32910 7112 32966
rect 7168 32910 7236 32966
rect 7292 32910 7360 32966
rect 7416 32910 7426 32966
rect 6358 32842 7426 32910
rect 6358 32786 6368 32842
rect 6424 32786 6492 32842
rect 6548 32786 6616 32842
rect 6672 32786 6740 32842
rect 6796 32786 6864 32842
rect 6920 32786 6988 32842
rect 7044 32786 7112 32842
rect 7168 32786 7236 32842
rect 7292 32786 7360 32842
rect 7416 32786 7426 32842
rect 6358 32718 7426 32786
rect 6358 32662 6368 32718
rect 6424 32662 6492 32718
rect 6548 32662 6616 32718
rect 6672 32662 6740 32718
rect 6796 32662 6864 32718
rect 6920 32662 6988 32718
rect 7044 32662 7112 32718
rect 7168 32662 7236 32718
rect 7292 32662 7360 32718
rect 7416 32662 7426 32718
rect 6358 32594 7426 32662
rect 6358 32538 6368 32594
rect 6424 32538 6492 32594
rect 6548 32538 6616 32594
rect 6672 32538 6740 32594
rect 6796 32538 6864 32594
rect 6920 32538 6988 32594
rect 7044 32538 7112 32594
rect 7168 32538 7236 32594
rect 7292 32538 7360 32594
rect 7416 32538 7426 32594
rect 6358 32470 7426 32538
rect 6358 32414 6368 32470
rect 6424 32414 6492 32470
rect 6548 32414 6616 32470
rect 6672 32414 6740 32470
rect 6796 32414 6864 32470
rect 6920 32414 6988 32470
rect 7044 32414 7112 32470
rect 7168 32414 7236 32470
rect 7292 32414 7360 32470
rect 7416 32414 7426 32470
rect 6358 32346 7426 32414
rect 6358 32290 6368 32346
rect 6424 32290 6492 32346
rect 6548 32290 6616 32346
rect 6672 32290 6740 32346
rect 6796 32290 6864 32346
rect 6920 32290 6988 32346
rect 7044 32290 7112 32346
rect 7168 32290 7236 32346
rect 7292 32290 7360 32346
rect 7416 32290 7426 32346
rect 6358 32222 7426 32290
rect 6358 32166 6368 32222
rect 6424 32166 6492 32222
rect 6548 32166 6616 32222
rect 6672 32166 6740 32222
rect 6796 32166 6864 32222
rect 6920 32166 6988 32222
rect 7044 32166 7112 32222
rect 7168 32166 7236 32222
rect 7292 32166 7360 32222
rect 7416 32166 7426 32222
rect 6358 32098 7426 32166
rect 6358 32042 6368 32098
rect 6424 32042 6492 32098
rect 6548 32042 6616 32098
rect 6672 32042 6740 32098
rect 6796 32042 6864 32098
rect 6920 32042 6988 32098
rect 7044 32042 7112 32098
rect 7168 32042 7236 32098
rect 7292 32042 7360 32098
rect 7416 32042 7426 32098
rect 6358 32032 7426 32042
rect 8741 34950 10553 34960
rect 8741 34894 8751 34950
rect 8807 34894 8875 34950
rect 8931 34894 8999 34950
rect 9055 34894 9123 34950
rect 9179 34894 9247 34950
rect 9303 34894 9371 34950
rect 9427 34894 9495 34950
rect 9551 34894 9619 34950
rect 9675 34894 9743 34950
rect 9799 34894 9867 34950
rect 9923 34894 9991 34950
rect 10047 34894 10115 34950
rect 10171 34894 10239 34950
rect 10295 34894 10363 34950
rect 10419 34894 10487 34950
rect 10543 34894 10553 34950
rect 8741 34826 10553 34894
rect 8741 34770 8751 34826
rect 8807 34770 8875 34826
rect 8931 34770 8999 34826
rect 9055 34770 9123 34826
rect 9179 34770 9247 34826
rect 9303 34770 9371 34826
rect 9427 34770 9495 34826
rect 9551 34770 9619 34826
rect 9675 34770 9743 34826
rect 9799 34770 9867 34826
rect 9923 34770 9991 34826
rect 10047 34770 10115 34826
rect 10171 34770 10239 34826
rect 10295 34770 10363 34826
rect 10419 34770 10487 34826
rect 10543 34770 10553 34826
rect 8741 34702 10553 34770
rect 8741 34646 8751 34702
rect 8807 34646 8875 34702
rect 8931 34646 8999 34702
rect 9055 34646 9123 34702
rect 9179 34646 9247 34702
rect 9303 34646 9371 34702
rect 9427 34646 9495 34702
rect 9551 34646 9619 34702
rect 9675 34646 9743 34702
rect 9799 34646 9867 34702
rect 9923 34646 9991 34702
rect 10047 34646 10115 34702
rect 10171 34646 10239 34702
rect 10295 34646 10363 34702
rect 10419 34646 10487 34702
rect 10543 34646 10553 34702
rect 8741 34578 10553 34646
rect 8741 34522 8751 34578
rect 8807 34522 8875 34578
rect 8931 34522 8999 34578
rect 9055 34522 9123 34578
rect 9179 34522 9247 34578
rect 9303 34522 9371 34578
rect 9427 34522 9495 34578
rect 9551 34522 9619 34578
rect 9675 34522 9743 34578
rect 9799 34522 9867 34578
rect 9923 34522 9991 34578
rect 10047 34522 10115 34578
rect 10171 34522 10239 34578
rect 10295 34522 10363 34578
rect 10419 34522 10487 34578
rect 10543 34522 10553 34578
rect 8741 34454 10553 34522
rect 8741 34398 8751 34454
rect 8807 34398 8875 34454
rect 8931 34398 8999 34454
rect 9055 34398 9123 34454
rect 9179 34398 9247 34454
rect 9303 34398 9371 34454
rect 9427 34398 9495 34454
rect 9551 34398 9619 34454
rect 9675 34398 9743 34454
rect 9799 34398 9867 34454
rect 9923 34398 9991 34454
rect 10047 34398 10115 34454
rect 10171 34398 10239 34454
rect 10295 34398 10363 34454
rect 10419 34398 10487 34454
rect 10543 34398 10553 34454
rect 8741 34330 10553 34398
rect 8741 34274 8751 34330
rect 8807 34274 8875 34330
rect 8931 34274 8999 34330
rect 9055 34274 9123 34330
rect 9179 34274 9247 34330
rect 9303 34274 9371 34330
rect 9427 34274 9495 34330
rect 9551 34274 9619 34330
rect 9675 34274 9743 34330
rect 9799 34274 9867 34330
rect 9923 34274 9991 34330
rect 10047 34274 10115 34330
rect 10171 34274 10239 34330
rect 10295 34274 10363 34330
rect 10419 34274 10487 34330
rect 10543 34274 10553 34330
rect 8741 34206 10553 34274
rect 8741 34150 8751 34206
rect 8807 34150 8875 34206
rect 8931 34150 8999 34206
rect 9055 34150 9123 34206
rect 9179 34150 9247 34206
rect 9303 34150 9371 34206
rect 9427 34150 9495 34206
rect 9551 34150 9619 34206
rect 9675 34150 9743 34206
rect 9799 34150 9867 34206
rect 9923 34150 9991 34206
rect 10047 34150 10115 34206
rect 10171 34150 10239 34206
rect 10295 34150 10363 34206
rect 10419 34150 10487 34206
rect 10543 34150 10553 34206
rect 8741 34082 10553 34150
rect 8741 34026 8751 34082
rect 8807 34026 8875 34082
rect 8931 34026 8999 34082
rect 9055 34026 9123 34082
rect 9179 34026 9247 34082
rect 9303 34026 9371 34082
rect 9427 34026 9495 34082
rect 9551 34026 9619 34082
rect 9675 34026 9743 34082
rect 9799 34026 9867 34082
rect 9923 34026 9991 34082
rect 10047 34026 10115 34082
rect 10171 34026 10239 34082
rect 10295 34026 10363 34082
rect 10419 34026 10487 34082
rect 10543 34026 10553 34082
rect 8741 33958 10553 34026
rect 8741 33902 8751 33958
rect 8807 33902 8875 33958
rect 8931 33902 8999 33958
rect 9055 33902 9123 33958
rect 9179 33902 9247 33958
rect 9303 33902 9371 33958
rect 9427 33902 9495 33958
rect 9551 33902 9619 33958
rect 9675 33902 9743 33958
rect 9799 33902 9867 33958
rect 9923 33902 9991 33958
rect 10047 33902 10115 33958
rect 10171 33902 10239 33958
rect 10295 33902 10363 33958
rect 10419 33902 10487 33958
rect 10543 33902 10553 33958
rect 8741 33834 10553 33902
rect 8741 33778 8751 33834
rect 8807 33778 8875 33834
rect 8931 33778 8999 33834
rect 9055 33778 9123 33834
rect 9179 33778 9247 33834
rect 9303 33778 9371 33834
rect 9427 33778 9495 33834
rect 9551 33778 9619 33834
rect 9675 33778 9743 33834
rect 9799 33778 9867 33834
rect 9923 33778 9991 33834
rect 10047 33778 10115 33834
rect 10171 33778 10239 33834
rect 10295 33778 10363 33834
rect 10419 33778 10487 33834
rect 10543 33778 10553 33834
rect 8741 33710 10553 33778
rect 8741 33654 8751 33710
rect 8807 33654 8875 33710
rect 8931 33654 8999 33710
rect 9055 33654 9123 33710
rect 9179 33654 9247 33710
rect 9303 33654 9371 33710
rect 9427 33654 9495 33710
rect 9551 33654 9619 33710
rect 9675 33654 9743 33710
rect 9799 33654 9867 33710
rect 9923 33654 9991 33710
rect 10047 33654 10115 33710
rect 10171 33654 10239 33710
rect 10295 33654 10363 33710
rect 10419 33654 10487 33710
rect 10543 33654 10553 33710
rect 8741 33586 10553 33654
rect 8741 33530 8751 33586
rect 8807 33530 8875 33586
rect 8931 33530 8999 33586
rect 9055 33530 9123 33586
rect 9179 33530 9247 33586
rect 9303 33530 9371 33586
rect 9427 33530 9495 33586
rect 9551 33530 9619 33586
rect 9675 33530 9743 33586
rect 9799 33530 9867 33586
rect 9923 33530 9991 33586
rect 10047 33530 10115 33586
rect 10171 33530 10239 33586
rect 10295 33530 10363 33586
rect 10419 33530 10487 33586
rect 10543 33530 10553 33586
rect 8741 33462 10553 33530
rect 8741 33406 8751 33462
rect 8807 33406 8875 33462
rect 8931 33406 8999 33462
rect 9055 33406 9123 33462
rect 9179 33406 9247 33462
rect 9303 33406 9371 33462
rect 9427 33406 9495 33462
rect 9551 33406 9619 33462
rect 9675 33406 9743 33462
rect 9799 33406 9867 33462
rect 9923 33406 9991 33462
rect 10047 33406 10115 33462
rect 10171 33406 10239 33462
rect 10295 33406 10363 33462
rect 10419 33406 10487 33462
rect 10543 33406 10553 33462
rect 8741 33338 10553 33406
rect 8741 33282 8751 33338
rect 8807 33282 8875 33338
rect 8931 33282 8999 33338
rect 9055 33282 9123 33338
rect 9179 33282 9247 33338
rect 9303 33282 9371 33338
rect 9427 33282 9495 33338
rect 9551 33282 9619 33338
rect 9675 33282 9743 33338
rect 9799 33282 9867 33338
rect 9923 33282 9991 33338
rect 10047 33282 10115 33338
rect 10171 33282 10239 33338
rect 10295 33282 10363 33338
rect 10419 33282 10487 33338
rect 10543 33282 10553 33338
rect 8741 33214 10553 33282
rect 8741 33158 8751 33214
rect 8807 33158 8875 33214
rect 8931 33158 8999 33214
rect 9055 33158 9123 33214
rect 9179 33158 9247 33214
rect 9303 33158 9371 33214
rect 9427 33158 9495 33214
rect 9551 33158 9619 33214
rect 9675 33158 9743 33214
rect 9799 33158 9867 33214
rect 9923 33158 9991 33214
rect 10047 33158 10115 33214
rect 10171 33158 10239 33214
rect 10295 33158 10363 33214
rect 10419 33158 10487 33214
rect 10543 33158 10553 33214
rect 8741 33090 10553 33158
rect 8741 33034 8751 33090
rect 8807 33034 8875 33090
rect 8931 33034 8999 33090
rect 9055 33034 9123 33090
rect 9179 33034 9247 33090
rect 9303 33034 9371 33090
rect 9427 33034 9495 33090
rect 9551 33034 9619 33090
rect 9675 33034 9743 33090
rect 9799 33034 9867 33090
rect 9923 33034 9991 33090
rect 10047 33034 10115 33090
rect 10171 33034 10239 33090
rect 10295 33034 10363 33090
rect 10419 33034 10487 33090
rect 10543 33034 10553 33090
rect 8741 32966 10553 33034
rect 8741 32910 8751 32966
rect 8807 32910 8875 32966
rect 8931 32910 8999 32966
rect 9055 32910 9123 32966
rect 9179 32910 9247 32966
rect 9303 32910 9371 32966
rect 9427 32910 9495 32966
rect 9551 32910 9619 32966
rect 9675 32910 9743 32966
rect 9799 32910 9867 32966
rect 9923 32910 9991 32966
rect 10047 32910 10115 32966
rect 10171 32910 10239 32966
rect 10295 32910 10363 32966
rect 10419 32910 10487 32966
rect 10543 32910 10553 32966
rect 8741 32842 10553 32910
rect 8741 32786 8751 32842
rect 8807 32786 8875 32842
rect 8931 32786 8999 32842
rect 9055 32786 9123 32842
rect 9179 32786 9247 32842
rect 9303 32786 9371 32842
rect 9427 32786 9495 32842
rect 9551 32786 9619 32842
rect 9675 32786 9743 32842
rect 9799 32786 9867 32842
rect 9923 32786 9991 32842
rect 10047 32786 10115 32842
rect 10171 32786 10239 32842
rect 10295 32786 10363 32842
rect 10419 32786 10487 32842
rect 10543 32786 10553 32842
rect 8741 32718 10553 32786
rect 8741 32662 8751 32718
rect 8807 32662 8875 32718
rect 8931 32662 8999 32718
rect 9055 32662 9123 32718
rect 9179 32662 9247 32718
rect 9303 32662 9371 32718
rect 9427 32662 9495 32718
rect 9551 32662 9619 32718
rect 9675 32662 9743 32718
rect 9799 32662 9867 32718
rect 9923 32662 9991 32718
rect 10047 32662 10115 32718
rect 10171 32662 10239 32718
rect 10295 32662 10363 32718
rect 10419 32662 10487 32718
rect 10543 32662 10553 32718
rect 8741 32594 10553 32662
rect 8741 32538 8751 32594
rect 8807 32538 8875 32594
rect 8931 32538 8999 32594
rect 9055 32538 9123 32594
rect 9179 32538 9247 32594
rect 9303 32538 9371 32594
rect 9427 32538 9495 32594
rect 9551 32538 9619 32594
rect 9675 32538 9743 32594
rect 9799 32538 9867 32594
rect 9923 32538 9991 32594
rect 10047 32538 10115 32594
rect 10171 32538 10239 32594
rect 10295 32538 10363 32594
rect 10419 32538 10487 32594
rect 10543 32538 10553 32594
rect 8741 32470 10553 32538
rect 8741 32414 8751 32470
rect 8807 32414 8875 32470
rect 8931 32414 8999 32470
rect 9055 32414 9123 32470
rect 9179 32414 9247 32470
rect 9303 32414 9371 32470
rect 9427 32414 9495 32470
rect 9551 32414 9619 32470
rect 9675 32414 9743 32470
rect 9799 32414 9867 32470
rect 9923 32414 9991 32470
rect 10047 32414 10115 32470
rect 10171 32414 10239 32470
rect 10295 32414 10363 32470
rect 10419 32414 10487 32470
rect 10543 32414 10553 32470
rect 8741 32346 10553 32414
rect 8741 32290 8751 32346
rect 8807 32290 8875 32346
rect 8931 32290 8999 32346
rect 9055 32290 9123 32346
rect 9179 32290 9247 32346
rect 9303 32290 9371 32346
rect 9427 32290 9495 32346
rect 9551 32290 9619 32346
rect 9675 32290 9743 32346
rect 9799 32290 9867 32346
rect 9923 32290 9991 32346
rect 10047 32290 10115 32346
rect 10171 32290 10239 32346
rect 10295 32290 10363 32346
rect 10419 32290 10487 32346
rect 10543 32290 10553 32346
rect 8741 32222 10553 32290
rect 8741 32166 8751 32222
rect 8807 32166 8875 32222
rect 8931 32166 8999 32222
rect 9055 32166 9123 32222
rect 9179 32166 9247 32222
rect 9303 32166 9371 32222
rect 9427 32166 9495 32222
rect 9551 32166 9619 32222
rect 9675 32166 9743 32222
rect 9799 32166 9867 32222
rect 9923 32166 9991 32222
rect 10047 32166 10115 32222
rect 10171 32166 10239 32222
rect 10295 32166 10363 32222
rect 10419 32166 10487 32222
rect 10543 32166 10553 32222
rect 8741 32098 10553 32166
rect 8741 32042 8751 32098
rect 8807 32042 8875 32098
rect 8931 32042 8999 32098
rect 9055 32042 9123 32098
rect 9179 32042 9247 32098
rect 9303 32042 9371 32098
rect 9427 32042 9495 32098
rect 9551 32042 9619 32098
rect 9675 32042 9743 32098
rect 9799 32042 9867 32098
rect 9923 32042 9991 32098
rect 10047 32042 10115 32098
rect 10171 32042 10239 32098
rect 10295 32042 10363 32098
rect 10419 32042 10487 32098
rect 10543 32042 10553 32098
rect 8741 32032 10553 32042
rect 12842 34950 13910 34960
rect 12842 34894 12852 34950
rect 12908 34894 12976 34950
rect 13032 34894 13100 34950
rect 13156 34894 13224 34950
rect 13280 34894 13348 34950
rect 13404 34894 13472 34950
rect 13528 34894 13596 34950
rect 13652 34894 13720 34950
rect 13776 34894 13844 34950
rect 13900 34894 13910 34950
rect 12842 34826 13910 34894
rect 12842 34770 12852 34826
rect 12908 34770 12976 34826
rect 13032 34770 13100 34826
rect 13156 34770 13224 34826
rect 13280 34770 13348 34826
rect 13404 34770 13472 34826
rect 13528 34770 13596 34826
rect 13652 34770 13720 34826
rect 13776 34770 13844 34826
rect 13900 34770 13910 34826
rect 12842 34702 13910 34770
rect 12842 34646 12852 34702
rect 12908 34646 12976 34702
rect 13032 34646 13100 34702
rect 13156 34646 13224 34702
rect 13280 34646 13348 34702
rect 13404 34646 13472 34702
rect 13528 34646 13596 34702
rect 13652 34646 13720 34702
rect 13776 34646 13844 34702
rect 13900 34646 13910 34702
rect 12842 34578 13910 34646
rect 12842 34522 12852 34578
rect 12908 34522 12976 34578
rect 13032 34522 13100 34578
rect 13156 34522 13224 34578
rect 13280 34522 13348 34578
rect 13404 34522 13472 34578
rect 13528 34522 13596 34578
rect 13652 34522 13720 34578
rect 13776 34522 13844 34578
rect 13900 34522 13910 34578
rect 12842 34454 13910 34522
rect 12842 34398 12852 34454
rect 12908 34398 12976 34454
rect 13032 34398 13100 34454
rect 13156 34398 13224 34454
rect 13280 34398 13348 34454
rect 13404 34398 13472 34454
rect 13528 34398 13596 34454
rect 13652 34398 13720 34454
rect 13776 34398 13844 34454
rect 13900 34398 13910 34454
rect 12842 34330 13910 34398
rect 12842 34274 12852 34330
rect 12908 34274 12976 34330
rect 13032 34274 13100 34330
rect 13156 34274 13224 34330
rect 13280 34274 13348 34330
rect 13404 34274 13472 34330
rect 13528 34274 13596 34330
rect 13652 34274 13720 34330
rect 13776 34274 13844 34330
rect 13900 34274 13910 34330
rect 12842 34206 13910 34274
rect 12842 34150 12852 34206
rect 12908 34150 12976 34206
rect 13032 34150 13100 34206
rect 13156 34150 13224 34206
rect 13280 34150 13348 34206
rect 13404 34150 13472 34206
rect 13528 34150 13596 34206
rect 13652 34150 13720 34206
rect 13776 34150 13844 34206
rect 13900 34150 13910 34206
rect 12842 34082 13910 34150
rect 12842 34026 12852 34082
rect 12908 34026 12976 34082
rect 13032 34026 13100 34082
rect 13156 34026 13224 34082
rect 13280 34026 13348 34082
rect 13404 34026 13472 34082
rect 13528 34026 13596 34082
rect 13652 34026 13720 34082
rect 13776 34026 13844 34082
rect 13900 34026 13910 34082
rect 12842 33958 13910 34026
rect 12842 33902 12852 33958
rect 12908 33902 12976 33958
rect 13032 33902 13100 33958
rect 13156 33902 13224 33958
rect 13280 33902 13348 33958
rect 13404 33902 13472 33958
rect 13528 33902 13596 33958
rect 13652 33902 13720 33958
rect 13776 33902 13844 33958
rect 13900 33902 13910 33958
rect 12842 33834 13910 33902
rect 12842 33778 12852 33834
rect 12908 33778 12976 33834
rect 13032 33778 13100 33834
rect 13156 33778 13224 33834
rect 13280 33778 13348 33834
rect 13404 33778 13472 33834
rect 13528 33778 13596 33834
rect 13652 33778 13720 33834
rect 13776 33778 13844 33834
rect 13900 33778 13910 33834
rect 12842 33710 13910 33778
rect 12842 33654 12852 33710
rect 12908 33654 12976 33710
rect 13032 33654 13100 33710
rect 13156 33654 13224 33710
rect 13280 33654 13348 33710
rect 13404 33654 13472 33710
rect 13528 33654 13596 33710
rect 13652 33654 13720 33710
rect 13776 33654 13844 33710
rect 13900 33654 13910 33710
rect 12842 33586 13910 33654
rect 12842 33530 12852 33586
rect 12908 33530 12976 33586
rect 13032 33530 13100 33586
rect 13156 33530 13224 33586
rect 13280 33530 13348 33586
rect 13404 33530 13472 33586
rect 13528 33530 13596 33586
rect 13652 33530 13720 33586
rect 13776 33530 13844 33586
rect 13900 33530 13910 33586
rect 12842 33462 13910 33530
rect 12842 33406 12852 33462
rect 12908 33406 12976 33462
rect 13032 33406 13100 33462
rect 13156 33406 13224 33462
rect 13280 33406 13348 33462
rect 13404 33406 13472 33462
rect 13528 33406 13596 33462
rect 13652 33406 13720 33462
rect 13776 33406 13844 33462
rect 13900 33406 13910 33462
rect 12842 33338 13910 33406
rect 12842 33282 12852 33338
rect 12908 33282 12976 33338
rect 13032 33282 13100 33338
rect 13156 33282 13224 33338
rect 13280 33282 13348 33338
rect 13404 33282 13472 33338
rect 13528 33282 13596 33338
rect 13652 33282 13720 33338
rect 13776 33282 13844 33338
rect 13900 33282 13910 33338
rect 12842 33214 13910 33282
rect 12842 33158 12852 33214
rect 12908 33158 12976 33214
rect 13032 33158 13100 33214
rect 13156 33158 13224 33214
rect 13280 33158 13348 33214
rect 13404 33158 13472 33214
rect 13528 33158 13596 33214
rect 13652 33158 13720 33214
rect 13776 33158 13844 33214
rect 13900 33158 13910 33214
rect 12842 33090 13910 33158
rect 12842 33034 12852 33090
rect 12908 33034 12976 33090
rect 13032 33034 13100 33090
rect 13156 33034 13224 33090
rect 13280 33034 13348 33090
rect 13404 33034 13472 33090
rect 13528 33034 13596 33090
rect 13652 33034 13720 33090
rect 13776 33034 13844 33090
rect 13900 33034 13910 33090
rect 12842 32966 13910 33034
rect 12842 32910 12852 32966
rect 12908 32910 12976 32966
rect 13032 32910 13100 32966
rect 13156 32910 13224 32966
rect 13280 32910 13348 32966
rect 13404 32910 13472 32966
rect 13528 32910 13596 32966
rect 13652 32910 13720 32966
rect 13776 32910 13844 32966
rect 13900 32910 13910 32966
rect 12842 32842 13910 32910
rect 12842 32786 12852 32842
rect 12908 32786 12976 32842
rect 13032 32786 13100 32842
rect 13156 32786 13224 32842
rect 13280 32786 13348 32842
rect 13404 32786 13472 32842
rect 13528 32786 13596 32842
rect 13652 32786 13720 32842
rect 13776 32786 13844 32842
rect 13900 32786 13910 32842
rect 12842 32718 13910 32786
rect 12842 32662 12852 32718
rect 12908 32662 12976 32718
rect 13032 32662 13100 32718
rect 13156 32662 13224 32718
rect 13280 32662 13348 32718
rect 13404 32662 13472 32718
rect 13528 32662 13596 32718
rect 13652 32662 13720 32718
rect 13776 32662 13844 32718
rect 13900 32662 13910 32718
rect 12842 32594 13910 32662
rect 12842 32538 12852 32594
rect 12908 32538 12976 32594
rect 13032 32538 13100 32594
rect 13156 32538 13224 32594
rect 13280 32538 13348 32594
rect 13404 32538 13472 32594
rect 13528 32538 13596 32594
rect 13652 32538 13720 32594
rect 13776 32538 13844 32594
rect 13900 32538 13910 32594
rect 12842 32470 13910 32538
rect 12842 32414 12852 32470
rect 12908 32414 12976 32470
rect 13032 32414 13100 32470
rect 13156 32414 13224 32470
rect 13280 32414 13348 32470
rect 13404 32414 13472 32470
rect 13528 32414 13596 32470
rect 13652 32414 13720 32470
rect 13776 32414 13844 32470
rect 13900 32414 13910 32470
rect 12842 32346 13910 32414
rect 12842 32290 12852 32346
rect 12908 32290 12976 32346
rect 13032 32290 13100 32346
rect 13156 32290 13224 32346
rect 13280 32290 13348 32346
rect 13404 32290 13472 32346
rect 13528 32290 13596 32346
rect 13652 32290 13720 32346
rect 13776 32290 13844 32346
rect 13900 32290 13910 32346
rect 12842 32222 13910 32290
rect 12842 32166 12852 32222
rect 12908 32166 12976 32222
rect 13032 32166 13100 32222
rect 13156 32166 13224 32222
rect 13280 32166 13348 32222
rect 13404 32166 13472 32222
rect 13528 32166 13596 32222
rect 13652 32166 13720 32222
rect 13776 32166 13844 32222
rect 13900 32166 13910 32222
rect 12842 32098 13910 32166
rect 12842 32042 12852 32098
rect 12908 32042 12976 32098
rect 13032 32042 13100 32098
rect 13156 32042 13224 32098
rect 13280 32042 13348 32098
rect 13404 32042 13472 32098
rect 13528 32042 13596 32098
rect 13652 32042 13720 32098
rect 13776 32042 13844 32098
rect 13900 32042 13910 32098
rect 12842 32032 13910 32042
rect 4129 32003 4205 32013
rect 2013 31906 2089 31974
rect 2013 31850 2023 31906
rect 2079 31850 2089 31906
rect 2013 31782 2089 31850
rect 2013 31726 2023 31782
rect 2079 31726 2089 31782
rect 2013 31658 2089 31726
rect 2013 31602 2023 31658
rect 2079 31602 2089 31658
rect 2013 31534 2089 31602
rect 2013 31478 2023 31534
rect 2079 31478 2089 31534
rect 2013 31410 2089 31478
rect 2013 31354 2023 31410
rect 2079 31354 2089 31410
rect 2013 31286 2089 31354
rect 2013 31230 2023 31286
rect 2079 31230 2089 31286
rect 2013 31162 2089 31230
rect 2013 31106 2023 31162
rect 2079 31106 2089 31162
rect 2013 31038 2089 31106
rect 2013 30982 2023 31038
rect 2079 30982 2089 31038
rect 2013 30914 2089 30982
rect 2013 30858 2023 30914
rect 2079 30858 2089 30914
rect 2013 30790 2089 30858
rect 2013 30734 2023 30790
rect 2079 30734 2089 30790
rect 2013 30666 2089 30734
rect 2013 30610 2023 30666
rect 2079 30610 2089 30666
rect 2013 30542 2089 30610
rect 2013 30486 2023 30542
rect 2079 30486 2089 30542
rect 2013 30418 2089 30486
rect 2013 30362 2023 30418
rect 2079 30362 2089 30418
rect 2013 30294 2089 30362
rect 2013 30238 2023 30294
rect 2079 30238 2089 30294
rect 2013 30170 2089 30238
rect 2013 30114 2023 30170
rect 2079 30114 2089 30170
rect 2013 30046 2089 30114
rect 2013 29990 2023 30046
rect 2079 29990 2089 30046
rect 2013 29922 2089 29990
rect 2013 29866 2023 29922
rect 2079 29866 2089 29922
rect 2013 29798 2089 29866
rect 2013 29742 2023 29798
rect 2079 29742 2089 29798
rect 2013 29674 2089 29742
rect 2013 29618 2023 29674
rect 2079 29618 2089 29674
rect 2013 29550 2089 29618
rect 2013 29494 2023 29550
rect 2079 29494 2089 29550
rect 2013 29426 2089 29494
rect 2013 29370 2023 29426
rect 2079 29370 2089 29426
rect 2013 29302 2089 29370
rect 2013 29246 2023 29302
rect 2079 29246 2089 29302
rect 2013 29178 2089 29246
rect 2013 29122 2023 29178
rect 2079 29122 2089 29178
rect 2013 29054 2089 29122
rect 2013 28998 2023 29054
rect 2079 28998 2089 29054
rect 1365 28879 1375 28935
rect 1431 28879 1441 28935
rect 1365 28811 1441 28879
rect 1365 28755 1375 28811
rect 1431 28755 1441 28811
rect 1365 28687 1441 28755
rect 1365 28631 1375 28687
rect 1431 28631 1441 28687
rect 1365 28563 1441 28631
rect 1365 28507 1375 28563
rect 1431 28507 1441 28563
rect 1365 28439 1441 28507
rect 1365 28383 1375 28439
rect 1431 28383 1441 28439
rect 1365 28315 1441 28383
rect 1365 28259 1375 28315
rect 1431 28259 1441 28315
rect 1365 28191 1441 28259
rect 1365 28135 1375 28191
rect 1431 28135 1441 28191
rect 1365 28067 1441 28135
rect 1365 28011 1375 28067
rect 1431 28011 1441 28067
rect 1365 27943 1441 28011
rect 1365 27887 1375 27943
rect 1431 27887 1441 27943
rect 1365 27819 1441 27887
rect 1365 27763 1375 27819
rect 1431 27763 1441 27819
rect 1365 27695 1441 27763
rect 1365 27639 1375 27695
rect 1431 27639 1441 27695
rect 1365 27571 1441 27639
rect 1365 27515 1375 27571
rect 1431 27515 1441 27571
rect 1365 27447 1441 27515
rect 1365 27391 1375 27447
rect 1431 27391 1441 27447
rect 1365 27323 1441 27391
rect 1365 27267 1375 27323
rect 1431 27267 1441 27323
rect 1365 27257 1441 27267
rect 1489 28922 1565 28932
rect 1489 28866 1499 28922
rect 1555 28866 1565 28922
rect 1489 28798 1565 28866
rect 2013 28930 2089 28998
rect 2013 28874 2023 28930
rect 2079 28874 2089 28930
rect 2013 28864 2089 28874
rect 4425 31750 6237 31760
rect 4425 31694 4435 31750
rect 4491 31694 4559 31750
rect 4615 31694 4683 31750
rect 4739 31694 4807 31750
rect 4863 31694 4931 31750
rect 4987 31694 5055 31750
rect 5111 31694 5179 31750
rect 5235 31694 5303 31750
rect 5359 31694 5427 31750
rect 5483 31694 5551 31750
rect 5607 31694 5675 31750
rect 5731 31694 5799 31750
rect 5855 31694 5923 31750
rect 5979 31694 6047 31750
rect 6103 31694 6171 31750
rect 6227 31694 6237 31750
rect 4425 31626 6237 31694
rect 4425 31570 4435 31626
rect 4491 31570 4559 31626
rect 4615 31570 4683 31626
rect 4739 31570 4807 31626
rect 4863 31570 4931 31626
rect 4987 31570 5055 31626
rect 5111 31570 5179 31626
rect 5235 31570 5303 31626
rect 5359 31570 5427 31626
rect 5483 31570 5551 31626
rect 5607 31570 5675 31626
rect 5731 31570 5799 31626
rect 5855 31570 5923 31626
rect 5979 31570 6047 31626
rect 6103 31570 6171 31626
rect 6227 31570 6237 31626
rect 4425 31502 6237 31570
rect 4425 31446 4435 31502
rect 4491 31446 4559 31502
rect 4615 31446 4683 31502
rect 4739 31446 4807 31502
rect 4863 31446 4931 31502
rect 4987 31446 5055 31502
rect 5111 31446 5179 31502
rect 5235 31446 5303 31502
rect 5359 31446 5427 31502
rect 5483 31446 5551 31502
rect 5607 31446 5675 31502
rect 5731 31446 5799 31502
rect 5855 31446 5923 31502
rect 5979 31446 6047 31502
rect 6103 31446 6171 31502
rect 6227 31446 6237 31502
rect 4425 31378 6237 31446
rect 4425 31322 4435 31378
rect 4491 31322 4559 31378
rect 4615 31322 4683 31378
rect 4739 31322 4807 31378
rect 4863 31322 4931 31378
rect 4987 31322 5055 31378
rect 5111 31322 5179 31378
rect 5235 31322 5303 31378
rect 5359 31322 5427 31378
rect 5483 31322 5551 31378
rect 5607 31322 5675 31378
rect 5731 31322 5799 31378
rect 5855 31322 5923 31378
rect 5979 31322 6047 31378
rect 6103 31322 6171 31378
rect 6227 31322 6237 31378
rect 4425 31254 6237 31322
rect 4425 31198 4435 31254
rect 4491 31198 4559 31254
rect 4615 31198 4683 31254
rect 4739 31198 4807 31254
rect 4863 31198 4931 31254
rect 4987 31198 5055 31254
rect 5111 31198 5179 31254
rect 5235 31198 5303 31254
rect 5359 31198 5427 31254
rect 5483 31198 5551 31254
rect 5607 31198 5675 31254
rect 5731 31198 5799 31254
rect 5855 31198 5923 31254
rect 5979 31198 6047 31254
rect 6103 31198 6171 31254
rect 6227 31198 6237 31254
rect 4425 31130 6237 31198
rect 4425 31074 4435 31130
rect 4491 31074 4559 31130
rect 4615 31074 4683 31130
rect 4739 31074 4807 31130
rect 4863 31074 4931 31130
rect 4987 31074 5055 31130
rect 5111 31074 5179 31130
rect 5235 31074 5303 31130
rect 5359 31074 5427 31130
rect 5483 31074 5551 31130
rect 5607 31074 5675 31130
rect 5731 31074 5799 31130
rect 5855 31074 5923 31130
rect 5979 31074 6047 31130
rect 6103 31074 6171 31130
rect 6227 31074 6237 31130
rect 4425 31006 6237 31074
rect 4425 30950 4435 31006
rect 4491 30950 4559 31006
rect 4615 30950 4683 31006
rect 4739 30950 4807 31006
rect 4863 30950 4931 31006
rect 4987 30950 5055 31006
rect 5111 30950 5179 31006
rect 5235 30950 5303 31006
rect 5359 30950 5427 31006
rect 5483 30950 5551 31006
rect 5607 30950 5675 31006
rect 5731 30950 5799 31006
rect 5855 30950 5923 31006
rect 5979 30950 6047 31006
rect 6103 30950 6171 31006
rect 6227 30950 6237 31006
rect 4425 30882 6237 30950
rect 4425 30826 4435 30882
rect 4491 30826 4559 30882
rect 4615 30826 4683 30882
rect 4739 30826 4807 30882
rect 4863 30826 4931 30882
rect 4987 30826 5055 30882
rect 5111 30826 5179 30882
rect 5235 30826 5303 30882
rect 5359 30826 5427 30882
rect 5483 30826 5551 30882
rect 5607 30826 5675 30882
rect 5731 30826 5799 30882
rect 5855 30826 5923 30882
rect 5979 30826 6047 30882
rect 6103 30826 6171 30882
rect 6227 30826 6237 30882
rect 4425 30758 6237 30826
rect 4425 30702 4435 30758
rect 4491 30702 4559 30758
rect 4615 30702 4683 30758
rect 4739 30702 4807 30758
rect 4863 30702 4931 30758
rect 4987 30702 5055 30758
rect 5111 30702 5179 30758
rect 5235 30702 5303 30758
rect 5359 30702 5427 30758
rect 5483 30702 5551 30758
rect 5607 30702 5675 30758
rect 5731 30702 5799 30758
rect 5855 30702 5923 30758
rect 5979 30702 6047 30758
rect 6103 30702 6171 30758
rect 6227 30702 6237 30758
rect 4425 30634 6237 30702
rect 4425 30578 4435 30634
rect 4491 30578 4559 30634
rect 4615 30578 4683 30634
rect 4739 30578 4807 30634
rect 4863 30578 4931 30634
rect 4987 30578 5055 30634
rect 5111 30578 5179 30634
rect 5235 30578 5303 30634
rect 5359 30578 5427 30634
rect 5483 30578 5551 30634
rect 5607 30578 5675 30634
rect 5731 30578 5799 30634
rect 5855 30578 5923 30634
rect 5979 30578 6047 30634
rect 6103 30578 6171 30634
rect 6227 30578 6237 30634
rect 4425 30510 6237 30578
rect 4425 30454 4435 30510
rect 4491 30454 4559 30510
rect 4615 30454 4683 30510
rect 4739 30454 4807 30510
rect 4863 30454 4931 30510
rect 4987 30454 5055 30510
rect 5111 30454 5179 30510
rect 5235 30454 5303 30510
rect 5359 30454 5427 30510
rect 5483 30454 5551 30510
rect 5607 30454 5675 30510
rect 5731 30454 5799 30510
rect 5855 30454 5923 30510
rect 5979 30454 6047 30510
rect 6103 30454 6171 30510
rect 6227 30454 6237 30510
rect 4425 30386 6237 30454
rect 4425 30330 4435 30386
rect 4491 30330 4559 30386
rect 4615 30330 4683 30386
rect 4739 30330 4807 30386
rect 4863 30330 4931 30386
rect 4987 30330 5055 30386
rect 5111 30330 5179 30386
rect 5235 30330 5303 30386
rect 5359 30330 5427 30386
rect 5483 30330 5551 30386
rect 5607 30330 5675 30386
rect 5731 30330 5799 30386
rect 5855 30330 5923 30386
rect 5979 30330 6047 30386
rect 6103 30330 6171 30386
rect 6227 30330 6237 30386
rect 4425 30262 6237 30330
rect 4425 30206 4435 30262
rect 4491 30206 4559 30262
rect 4615 30206 4683 30262
rect 4739 30206 4807 30262
rect 4863 30206 4931 30262
rect 4987 30206 5055 30262
rect 5111 30206 5179 30262
rect 5235 30206 5303 30262
rect 5359 30206 5427 30262
rect 5483 30206 5551 30262
rect 5607 30206 5675 30262
rect 5731 30206 5799 30262
rect 5855 30206 5923 30262
rect 5979 30206 6047 30262
rect 6103 30206 6171 30262
rect 6227 30206 6237 30262
rect 4425 30138 6237 30206
rect 4425 30082 4435 30138
rect 4491 30082 4559 30138
rect 4615 30082 4683 30138
rect 4739 30082 4807 30138
rect 4863 30082 4931 30138
rect 4987 30082 5055 30138
rect 5111 30082 5179 30138
rect 5235 30082 5303 30138
rect 5359 30082 5427 30138
rect 5483 30082 5551 30138
rect 5607 30082 5675 30138
rect 5731 30082 5799 30138
rect 5855 30082 5923 30138
rect 5979 30082 6047 30138
rect 6103 30082 6171 30138
rect 6227 30082 6237 30138
rect 4425 30014 6237 30082
rect 4425 29958 4435 30014
rect 4491 29958 4559 30014
rect 4615 29958 4683 30014
rect 4739 29958 4807 30014
rect 4863 29958 4931 30014
rect 4987 29958 5055 30014
rect 5111 29958 5179 30014
rect 5235 29958 5303 30014
rect 5359 29958 5427 30014
rect 5483 29958 5551 30014
rect 5607 29958 5675 30014
rect 5731 29958 5799 30014
rect 5855 29958 5923 30014
rect 5979 29958 6047 30014
rect 6103 29958 6171 30014
rect 6227 29958 6237 30014
rect 4425 29890 6237 29958
rect 4425 29834 4435 29890
rect 4491 29834 4559 29890
rect 4615 29834 4683 29890
rect 4739 29834 4807 29890
rect 4863 29834 4931 29890
rect 4987 29834 5055 29890
rect 5111 29834 5179 29890
rect 5235 29834 5303 29890
rect 5359 29834 5427 29890
rect 5483 29834 5551 29890
rect 5607 29834 5675 29890
rect 5731 29834 5799 29890
rect 5855 29834 5923 29890
rect 5979 29834 6047 29890
rect 6103 29834 6171 29890
rect 6227 29834 6237 29890
rect 4425 29766 6237 29834
rect 4425 29710 4435 29766
rect 4491 29710 4559 29766
rect 4615 29710 4683 29766
rect 4739 29710 4807 29766
rect 4863 29710 4931 29766
rect 4987 29710 5055 29766
rect 5111 29710 5179 29766
rect 5235 29710 5303 29766
rect 5359 29710 5427 29766
rect 5483 29710 5551 29766
rect 5607 29710 5675 29766
rect 5731 29710 5799 29766
rect 5855 29710 5923 29766
rect 5979 29710 6047 29766
rect 6103 29710 6171 29766
rect 6227 29710 6237 29766
rect 4425 29642 6237 29710
rect 4425 29586 4435 29642
rect 4491 29586 4559 29642
rect 4615 29586 4683 29642
rect 4739 29586 4807 29642
rect 4863 29586 4931 29642
rect 4987 29586 5055 29642
rect 5111 29586 5179 29642
rect 5235 29586 5303 29642
rect 5359 29586 5427 29642
rect 5483 29586 5551 29642
rect 5607 29586 5675 29642
rect 5731 29586 5799 29642
rect 5855 29586 5923 29642
rect 5979 29586 6047 29642
rect 6103 29586 6171 29642
rect 6227 29586 6237 29642
rect 4425 29518 6237 29586
rect 4425 29462 4435 29518
rect 4491 29462 4559 29518
rect 4615 29462 4683 29518
rect 4739 29462 4807 29518
rect 4863 29462 4931 29518
rect 4987 29462 5055 29518
rect 5111 29462 5179 29518
rect 5235 29462 5303 29518
rect 5359 29462 5427 29518
rect 5483 29462 5551 29518
rect 5607 29462 5675 29518
rect 5731 29462 5799 29518
rect 5855 29462 5923 29518
rect 5979 29462 6047 29518
rect 6103 29462 6171 29518
rect 6227 29462 6237 29518
rect 4425 29394 6237 29462
rect 4425 29338 4435 29394
rect 4491 29338 4559 29394
rect 4615 29338 4683 29394
rect 4739 29338 4807 29394
rect 4863 29338 4931 29394
rect 4987 29338 5055 29394
rect 5111 29338 5179 29394
rect 5235 29338 5303 29394
rect 5359 29338 5427 29394
rect 5483 29338 5551 29394
rect 5607 29338 5675 29394
rect 5731 29338 5799 29394
rect 5855 29338 5923 29394
rect 5979 29338 6047 29394
rect 6103 29338 6171 29394
rect 6227 29338 6237 29394
rect 4425 29270 6237 29338
rect 4425 29214 4435 29270
rect 4491 29214 4559 29270
rect 4615 29214 4683 29270
rect 4739 29214 4807 29270
rect 4863 29214 4931 29270
rect 4987 29214 5055 29270
rect 5111 29214 5179 29270
rect 5235 29214 5303 29270
rect 5359 29214 5427 29270
rect 5483 29214 5551 29270
rect 5607 29214 5675 29270
rect 5731 29214 5799 29270
rect 5855 29214 5923 29270
rect 5979 29214 6047 29270
rect 6103 29214 6171 29270
rect 6227 29214 6237 29270
rect 4425 29146 6237 29214
rect 4425 29090 4435 29146
rect 4491 29090 4559 29146
rect 4615 29090 4683 29146
rect 4739 29090 4807 29146
rect 4863 29090 4931 29146
rect 4987 29090 5055 29146
rect 5111 29090 5179 29146
rect 5235 29090 5303 29146
rect 5359 29090 5427 29146
rect 5483 29090 5551 29146
rect 5607 29090 5675 29146
rect 5731 29090 5799 29146
rect 5855 29090 5923 29146
rect 5979 29090 6047 29146
rect 6103 29090 6171 29146
rect 6227 29090 6237 29146
rect 4425 29022 6237 29090
rect 4425 28966 4435 29022
rect 4491 28966 4559 29022
rect 4615 28966 4683 29022
rect 4739 28966 4807 29022
rect 4863 28966 4931 29022
rect 4987 28966 5055 29022
rect 5111 28966 5179 29022
rect 5235 28966 5303 29022
rect 5359 28966 5427 29022
rect 5483 28966 5551 29022
rect 5607 28966 5675 29022
rect 5731 28966 5799 29022
rect 5855 28966 5923 29022
rect 5979 28966 6047 29022
rect 6103 28966 6171 29022
rect 6227 28966 6237 29022
rect 4425 28898 6237 28966
rect 4425 28842 4435 28898
rect 4491 28842 4559 28898
rect 4615 28842 4683 28898
rect 4739 28842 4807 28898
rect 4863 28842 4931 28898
rect 4987 28842 5055 28898
rect 5111 28842 5179 28898
rect 5235 28842 5303 28898
rect 5359 28842 5427 28898
rect 5483 28842 5551 28898
rect 5607 28842 5675 28898
rect 5731 28842 5799 28898
rect 5855 28842 5923 28898
rect 5979 28842 6047 28898
rect 6103 28842 6171 28898
rect 6227 28842 6237 28898
rect 4425 28832 6237 28842
rect 7552 31750 8620 31760
rect 7552 31694 7562 31750
rect 7618 31694 7686 31750
rect 7742 31694 7810 31750
rect 7866 31694 7934 31750
rect 7990 31694 8058 31750
rect 8114 31694 8182 31750
rect 8238 31694 8306 31750
rect 8362 31694 8430 31750
rect 8486 31694 8554 31750
rect 8610 31694 8620 31750
rect 7552 31626 8620 31694
rect 7552 31570 7562 31626
rect 7618 31570 7686 31626
rect 7742 31570 7810 31626
rect 7866 31570 7934 31626
rect 7990 31570 8058 31626
rect 8114 31570 8182 31626
rect 8238 31570 8306 31626
rect 8362 31570 8430 31626
rect 8486 31570 8554 31626
rect 8610 31570 8620 31626
rect 7552 31502 8620 31570
rect 7552 31446 7562 31502
rect 7618 31446 7686 31502
rect 7742 31446 7810 31502
rect 7866 31446 7934 31502
rect 7990 31446 8058 31502
rect 8114 31446 8182 31502
rect 8238 31446 8306 31502
rect 8362 31446 8430 31502
rect 8486 31446 8554 31502
rect 8610 31446 8620 31502
rect 7552 31378 8620 31446
rect 7552 31322 7562 31378
rect 7618 31322 7686 31378
rect 7742 31322 7810 31378
rect 7866 31322 7934 31378
rect 7990 31322 8058 31378
rect 8114 31322 8182 31378
rect 8238 31322 8306 31378
rect 8362 31322 8430 31378
rect 8486 31322 8554 31378
rect 8610 31322 8620 31378
rect 7552 31254 8620 31322
rect 7552 31198 7562 31254
rect 7618 31198 7686 31254
rect 7742 31198 7810 31254
rect 7866 31198 7934 31254
rect 7990 31198 8058 31254
rect 8114 31198 8182 31254
rect 8238 31198 8306 31254
rect 8362 31198 8430 31254
rect 8486 31198 8554 31254
rect 8610 31198 8620 31254
rect 7552 31130 8620 31198
rect 7552 31074 7562 31130
rect 7618 31074 7686 31130
rect 7742 31074 7810 31130
rect 7866 31074 7934 31130
rect 7990 31074 8058 31130
rect 8114 31074 8182 31130
rect 8238 31074 8306 31130
rect 8362 31074 8430 31130
rect 8486 31074 8554 31130
rect 8610 31074 8620 31130
rect 7552 31006 8620 31074
rect 7552 30950 7562 31006
rect 7618 30950 7686 31006
rect 7742 30950 7810 31006
rect 7866 30950 7934 31006
rect 7990 30950 8058 31006
rect 8114 30950 8182 31006
rect 8238 30950 8306 31006
rect 8362 30950 8430 31006
rect 8486 30950 8554 31006
rect 8610 30950 8620 31006
rect 7552 30882 8620 30950
rect 7552 30826 7562 30882
rect 7618 30826 7686 30882
rect 7742 30826 7810 30882
rect 7866 30826 7934 30882
rect 7990 30826 8058 30882
rect 8114 30826 8182 30882
rect 8238 30826 8306 30882
rect 8362 30826 8430 30882
rect 8486 30826 8554 30882
rect 8610 30826 8620 30882
rect 7552 30758 8620 30826
rect 7552 30702 7562 30758
rect 7618 30702 7686 30758
rect 7742 30702 7810 30758
rect 7866 30702 7934 30758
rect 7990 30702 8058 30758
rect 8114 30702 8182 30758
rect 8238 30702 8306 30758
rect 8362 30702 8430 30758
rect 8486 30702 8554 30758
rect 8610 30702 8620 30758
rect 7552 30634 8620 30702
rect 7552 30578 7562 30634
rect 7618 30578 7686 30634
rect 7742 30578 7810 30634
rect 7866 30578 7934 30634
rect 7990 30578 8058 30634
rect 8114 30578 8182 30634
rect 8238 30578 8306 30634
rect 8362 30578 8430 30634
rect 8486 30578 8554 30634
rect 8610 30578 8620 30634
rect 7552 30510 8620 30578
rect 7552 30454 7562 30510
rect 7618 30454 7686 30510
rect 7742 30454 7810 30510
rect 7866 30454 7934 30510
rect 7990 30454 8058 30510
rect 8114 30454 8182 30510
rect 8238 30454 8306 30510
rect 8362 30454 8430 30510
rect 8486 30454 8554 30510
rect 8610 30454 8620 30510
rect 7552 30386 8620 30454
rect 7552 30330 7562 30386
rect 7618 30330 7686 30386
rect 7742 30330 7810 30386
rect 7866 30330 7934 30386
rect 7990 30330 8058 30386
rect 8114 30330 8182 30386
rect 8238 30330 8306 30386
rect 8362 30330 8430 30386
rect 8486 30330 8554 30386
rect 8610 30330 8620 30386
rect 7552 30262 8620 30330
rect 7552 30206 7562 30262
rect 7618 30206 7686 30262
rect 7742 30206 7810 30262
rect 7866 30206 7934 30262
rect 7990 30206 8058 30262
rect 8114 30206 8182 30262
rect 8238 30206 8306 30262
rect 8362 30206 8430 30262
rect 8486 30206 8554 30262
rect 8610 30206 8620 30262
rect 7552 30138 8620 30206
rect 7552 30082 7562 30138
rect 7618 30082 7686 30138
rect 7742 30082 7810 30138
rect 7866 30082 7934 30138
rect 7990 30082 8058 30138
rect 8114 30082 8182 30138
rect 8238 30082 8306 30138
rect 8362 30082 8430 30138
rect 8486 30082 8554 30138
rect 8610 30082 8620 30138
rect 7552 30014 8620 30082
rect 7552 29958 7562 30014
rect 7618 29958 7686 30014
rect 7742 29958 7810 30014
rect 7866 29958 7934 30014
rect 7990 29958 8058 30014
rect 8114 29958 8182 30014
rect 8238 29958 8306 30014
rect 8362 29958 8430 30014
rect 8486 29958 8554 30014
rect 8610 29958 8620 30014
rect 7552 29890 8620 29958
rect 7552 29834 7562 29890
rect 7618 29834 7686 29890
rect 7742 29834 7810 29890
rect 7866 29834 7934 29890
rect 7990 29834 8058 29890
rect 8114 29834 8182 29890
rect 8238 29834 8306 29890
rect 8362 29834 8430 29890
rect 8486 29834 8554 29890
rect 8610 29834 8620 29890
rect 7552 29766 8620 29834
rect 7552 29710 7562 29766
rect 7618 29710 7686 29766
rect 7742 29710 7810 29766
rect 7866 29710 7934 29766
rect 7990 29710 8058 29766
rect 8114 29710 8182 29766
rect 8238 29710 8306 29766
rect 8362 29710 8430 29766
rect 8486 29710 8554 29766
rect 8610 29710 8620 29766
rect 7552 29642 8620 29710
rect 7552 29586 7562 29642
rect 7618 29586 7686 29642
rect 7742 29586 7810 29642
rect 7866 29586 7934 29642
rect 7990 29586 8058 29642
rect 8114 29586 8182 29642
rect 8238 29586 8306 29642
rect 8362 29586 8430 29642
rect 8486 29586 8554 29642
rect 8610 29586 8620 29642
rect 7552 29518 8620 29586
rect 7552 29462 7562 29518
rect 7618 29462 7686 29518
rect 7742 29462 7810 29518
rect 7866 29462 7934 29518
rect 7990 29462 8058 29518
rect 8114 29462 8182 29518
rect 8238 29462 8306 29518
rect 8362 29462 8430 29518
rect 8486 29462 8554 29518
rect 8610 29462 8620 29518
rect 7552 29394 8620 29462
rect 7552 29338 7562 29394
rect 7618 29338 7686 29394
rect 7742 29338 7810 29394
rect 7866 29338 7934 29394
rect 7990 29338 8058 29394
rect 8114 29338 8182 29394
rect 8238 29338 8306 29394
rect 8362 29338 8430 29394
rect 8486 29338 8554 29394
rect 8610 29338 8620 29394
rect 7552 29270 8620 29338
rect 7552 29214 7562 29270
rect 7618 29214 7686 29270
rect 7742 29214 7810 29270
rect 7866 29214 7934 29270
rect 7990 29214 8058 29270
rect 8114 29214 8182 29270
rect 8238 29214 8306 29270
rect 8362 29214 8430 29270
rect 8486 29214 8554 29270
rect 8610 29214 8620 29270
rect 7552 29146 8620 29214
rect 7552 29090 7562 29146
rect 7618 29090 7686 29146
rect 7742 29090 7810 29146
rect 7866 29090 7934 29146
rect 7990 29090 8058 29146
rect 8114 29090 8182 29146
rect 8238 29090 8306 29146
rect 8362 29090 8430 29146
rect 8486 29090 8554 29146
rect 8610 29090 8620 29146
rect 7552 29022 8620 29090
rect 7552 28966 7562 29022
rect 7618 28966 7686 29022
rect 7742 28966 7810 29022
rect 7866 28966 7934 29022
rect 7990 28966 8058 29022
rect 8114 28966 8182 29022
rect 8238 28966 8306 29022
rect 8362 28966 8430 29022
rect 8486 28966 8554 29022
rect 8610 28966 8620 29022
rect 7552 28898 8620 28966
rect 7552 28842 7562 28898
rect 7618 28842 7686 28898
rect 7742 28842 7810 28898
rect 7866 28842 7934 28898
rect 7990 28842 8058 28898
rect 8114 28842 8182 28898
rect 8238 28842 8306 28898
rect 8362 28842 8430 28898
rect 8486 28842 8554 28898
rect 8610 28842 8620 28898
rect 7552 28832 8620 28842
rect 10669 31750 12481 31760
rect 10669 31694 10679 31750
rect 10735 31694 10803 31750
rect 10859 31694 10927 31750
rect 10983 31694 11051 31750
rect 11107 31694 11175 31750
rect 11231 31694 11299 31750
rect 11355 31694 11423 31750
rect 11479 31694 11547 31750
rect 11603 31694 11671 31750
rect 11727 31694 11795 31750
rect 11851 31694 11919 31750
rect 11975 31694 12043 31750
rect 12099 31694 12167 31750
rect 12223 31694 12291 31750
rect 12347 31694 12415 31750
rect 12471 31694 12481 31750
rect 10669 31626 12481 31694
rect 10669 31570 10679 31626
rect 10735 31570 10803 31626
rect 10859 31570 10927 31626
rect 10983 31570 11051 31626
rect 11107 31570 11175 31626
rect 11231 31570 11299 31626
rect 11355 31570 11423 31626
rect 11479 31570 11547 31626
rect 11603 31570 11671 31626
rect 11727 31570 11795 31626
rect 11851 31570 11919 31626
rect 11975 31570 12043 31626
rect 12099 31570 12167 31626
rect 12223 31570 12291 31626
rect 12347 31570 12415 31626
rect 12471 31570 12481 31626
rect 10669 31502 12481 31570
rect 10669 31446 10679 31502
rect 10735 31446 10803 31502
rect 10859 31446 10927 31502
rect 10983 31446 11051 31502
rect 11107 31446 11175 31502
rect 11231 31446 11299 31502
rect 11355 31446 11423 31502
rect 11479 31446 11547 31502
rect 11603 31446 11671 31502
rect 11727 31446 11795 31502
rect 11851 31446 11919 31502
rect 11975 31446 12043 31502
rect 12099 31446 12167 31502
rect 12223 31446 12291 31502
rect 12347 31446 12415 31502
rect 12471 31446 12481 31502
rect 10669 31378 12481 31446
rect 10669 31322 10679 31378
rect 10735 31322 10803 31378
rect 10859 31322 10927 31378
rect 10983 31322 11051 31378
rect 11107 31322 11175 31378
rect 11231 31322 11299 31378
rect 11355 31322 11423 31378
rect 11479 31322 11547 31378
rect 11603 31322 11671 31378
rect 11727 31322 11795 31378
rect 11851 31322 11919 31378
rect 11975 31322 12043 31378
rect 12099 31322 12167 31378
rect 12223 31322 12291 31378
rect 12347 31322 12415 31378
rect 12471 31322 12481 31378
rect 10669 31254 12481 31322
rect 10669 31198 10679 31254
rect 10735 31198 10803 31254
rect 10859 31198 10927 31254
rect 10983 31198 11051 31254
rect 11107 31198 11175 31254
rect 11231 31198 11299 31254
rect 11355 31198 11423 31254
rect 11479 31198 11547 31254
rect 11603 31198 11671 31254
rect 11727 31198 11795 31254
rect 11851 31198 11919 31254
rect 11975 31198 12043 31254
rect 12099 31198 12167 31254
rect 12223 31198 12291 31254
rect 12347 31198 12415 31254
rect 12471 31198 12481 31254
rect 10669 31130 12481 31198
rect 10669 31074 10679 31130
rect 10735 31074 10803 31130
rect 10859 31074 10927 31130
rect 10983 31074 11051 31130
rect 11107 31074 11175 31130
rect 11231 31074 11299 31130
rect 11355 31074 11423 31130
rect 11479 31074 11547 31130
rect 11603 31074 11671 31130
rect 11727 31074 11795 31130
rect 11851 31074 11919 31130
rect 11975 31074 12043 31130
rect 12099 31074 12167 31130
rect 12223 31074 12291 31130
rect 12347 31074 12415 31130
rect 12471 31074 12481 31130
rect 10669 31006 12481 31074
rect 10669 30950 10679 31006
rect 10735 30950 10803 31006
rect 10859 30950 10927 31006
rect 10983 30950 11051 31006
rect 11107 30950 11175 31006
rect 11231 30950 11299 31006
rect 11355 30950 11423 31006
rect 11479 30950 11547 31006
rect 11603 30950 11671 31006
rect 11727 30950 11795 31006
rect 11851 30950 11919 31006
rect 11975 30950 12043 31006
rect 12099 30950 12167 31006
rect 12223 30950 12291 31006
rect 12347 30950 12415 31006
rect 12471 30950 12481 31006
rect 10669 30882 12481 30950
rect 10669 30826 10679 30882
rect 10735 30826 10803 30882
rect 10859 30826 10927 30882
rect 10983 30826 11051 30882
rect 11107 30826 11175 30882
rect 11231 30826 11299 30882
rect 11355 30826 11423 30882
rect 11479 30826 11547 30882
rect 11603 30826 11671 30882
rect 11727 30826 11795 30882
rect 11851 30826 11919 30882
rect 11975 30826 12043 30882
rect 12099 30826 12167 30882
rect 12223 30826 12291 30882
rect 12347 30826 12415 30882
rect 12471 30826 12481 30882
rect 10669 30758 12481 30826
rect 10669 30702 10679 30758
rect 10735 30702 10803 30758
rect 10859 30702 10927 30758
rect 10983 30702 11051 30758
rect 11107 30702 11175 30758
rect 11231 30702 11299 30758
rect 11355 30702 11423 30758
rect 11479 30702 11547 30758
rect 11603 30702 11671 30758
rect 11727 30702 11795 30758
rect 11851 30702 11919 30758
rect 11975 30702 12043 30758
rect 12099 30702 12167 30758
rect 12223 30702 12291 30758
rect 12347 30702 12415 30758
rect 12471 30702 12481 30758
rect 10669 30634 12481 30702
rect 10669 30578 10679 30634
rect 10735 30578 10803 30634
rect 10859 30578 10927 30634
rect 10983 30578 11051 30634
rect 11107 30578 11175 30634
rect 11231 30578 11299 30634
rect 11355 30578 11423 30634
rect 11479 30578 11547 30634
rect 11603 30578 11671 30634
rect 11727 30578 11795 30634
rect 11851 30578 11919 30634
rect 11975 30578 12043 30634
rect 12099 30578 12167 30634
rect 12223 30578 12291 30634
rect 12347 30578 12415 30634
rect 12471 30578 12481 30634
rect 10669 30510 12481 30578
rect 10669 30454 10679 30510
rect 10735 30454 10803 30510
rect 10859 30454 10927 30510
rect 10983 30454 11051 30510
rect 11107 30454 11175 30510
rect 11231 30454 11299 30510
rect 11355 30454 11423 30510
rect 11479 30454 11547 30510
rect 11603 30454 11671 30510
rect 11727 30454 11795 30510
rect 11851 30454 11919 30510
rect 11975 30454 12043 30510
rect 12099 30454 12167 30510
rect 12223 30454 12291 30510
rect 12347 30454 12415 30510
rect 12471 30454 12481 30510
rect 10669 30386 12481 30454
rect 10669 30330 10679 30386
rect 10735 30330 10803 30386
rect 10859 30330 10927 30386
rect 10983 30330 11051 30386
rect 11107 30330 11175 30386
rect 11231 30330 11299 30386
rect 11355 30330 11423 30386
rect 11479 30330 11547 30386
rect 11603 30330 11671 30386
rect 11727 30330 11795 30386
rect 11851 30330 11919 30386
rect 11975 30330 12043 30386
rect 12099 30330 12167 30386
rect 12223 30330 12291 30386
rect 12347 30330 12415 30386
rect 12471 30330 12481 30386
rect 10669 30262 12481 30330
rect 10669 30206 10679 30262
rect 10735 30206 10803 30262
rect 10859 30206 10927 30262
rect 10983 30206 11051 30262
rect 11107 30206 11175 30262
rect 11231 30206 11299 30262
rect 11355 30206 11423 30262
rect 11479 30206 11547 30262
rect 11603 30206 11671 30262
rect 11727 30206 11795 30262
rect 11851 30206 11919 30262
rect 11975 30206 12043 30262
rect 12099 30206 12167 30262
rect 12223 30206 12291 30262
rect 12347 30206 12415 30262
rect 12471 30206 12481 30262
rect 10669 30138 12481 30206
rect 10669 30082 10679 30138
rect 10735 30082 10803 30138
rect 10859 30082 10927 30138
rect 10983 30082 11051 30138
rect 11107 30082 11175 30138
rect 11231 30082 11299 30138
rect 11355 30082 11423 30138
rect 11479 30082 11547 30138
rect 11603 30082 11671 30138
rect 11727 30082 11795 30138
rect 11851 30082 11919 30138
rect 11975 30082 12043 30138
rect 12099 30082 12167 30138
rect 12223 30082 12291 30138
rect 12347 30082 12415 30138
rect 12471 30082 12481 30138
rect 10669 30014 12481 30082
rect 10669 29958 10679 30014
rect 10735 29958 10803 30014
rect 10859 29958 10927 30014
rect 10983 29958 11051 30014
rect 11107 29958 11175 30014
rect 11231 29958 11299 30014
rect 11355 29958 11423 30014
rect 11479 29958 11547 30014
rect 11603 29958 11671 30014
rect 11727 29958 11795 30014
rect 11851 29958 11919 30014
rect 11975 29958 12043 30014
rect 12099 29958 12167 30014
rect 12223 29958 12291 30014
rect 12347 29958 12415 30014
rect 12471 29958 12481 30014
rect 10669 29890 12481 29958
rect 10669 29834 10679 29890
rect 10735 29834 10803 29890
rect 10859 29834 10927 29890
rect 10983 29834 11051 29890
rect 11107 29834 11175 29890
rect 11231 29834 11299 29890
rect 11355 29834 11423 29890
rect 11479 29834 11547 29890
rect 11603 29834 11671 29890
rect 11727 29834 11795 29890
rect 11851 29834 11919 29890
rect 11975 29834 12043 29890
rect 12099 29834 12167 29890
rect 12223 29834 12291 29890
rect 12347 29834 12415 29890
rect 12471 29834 12481 29890
rect 10669 29766 12481 29834
rect 10669 29710 10679 29766
rect 10735 29710 10803 29766
rect 10859 29710 10927 29766
rect 10983 29710 11051 29766
rect 11107 29710 11175 29766
rect 11231 29710 11299 29766
rect 11355 29710 11423 29766
rect 11479 29710 11547 29766
rect 11603 29710 11671 29766
rect 11727 29710 11795 29766
rect 11851 29710 11919 29766
rect 11975 29710 12043 29766
rect 12099 29710 12167 29766
rect 12223 29710 12291 29766
rect 12347 29710 12415 29766
rect 12471 29710 12481 29766
rect 10669 29642 12481 29710
rect 10669 29586 10679 29642
rect 10735 29586 10803 29642
rect 10859 29586 10927 29642
rect 10983 29586 11051 29642
rect 11107 29586 11175 29642
rect 11231 29586 11299 29642
rect 11355 29586 11423 29642
rect 11479 29586 11547 29642
rect 11603 29586 11671 29642
rect 11727 29586 11795 29642
rect 11851 29586 11919 29642
rect 11975 29586 12043 29642
rect 12099 29586 12167 29642
rect 12223 29586 12291 29642
rect 12347 29586 12415 29642
rect 12471 29586 12481 29642
rect 10669 29518 12481 29586
rect 10669 29462 10679 29518
rect 10735 29462 10803 29518
rect 10859 29462 10927 29518
rect 10983 29462 11051 29518
rect 11107 29462 11175 29518
rect 11231 29462 11299 29518
rect 11355 29462 11423 29518
rect 11479 29462 11547 29518
rect 11603 29462 11671 29518
rect 11727 29462 11795 29518
rect 11851 29462 11919 29518
rect 11975 29462 12043 29518
rect 12099 29462 12167 29518
rect 12223 29462 12291 29518
rect 12347 29462 12415 29518
rect 12471 29462 12481 29518
rect 10669 29394 12481 29462
rect 10669 29338 10679 29394
rect 10735 29338 10803 29394
rect 10859 29338 10927 29394
rect 10983 29338 11051 29394
rect 11107 29338 11175 29394
rect 11231 29338 11299 29394
rect 11355 29338 11423 29394
rect 11479 29338 11547 29394
rect 11603 29338 11671 29394
rect 11727 29338 11795 29394
rect 11851 29338 11919 29394
rect 11975 29338 12043 29394
rect 12099 29338 12167 29394
rect 12223 29338 12291 29394
rect 12347 29338 12415 29394
rect 12471 29338 12481 29394
rect 10669 29270 12481 29338
rect 10669 29214 10679 29270
rect 10735 29214 10803 29270
rect 10859 29214 10927 29270
rect 10983 29214 11051 29270
rect 11107 29214 11175 29270
rect 11231 29214 11299 29270
rect 11355 29214 11423 29270
rect 11479 29214 11547 29270
rect 11603 29214 11671 29270
rect 11727 29214 11795 29270
rect 11851 29214 11919 29270
rect 11975 29214 12043 29270
rect 12099 29214 12167 29270
rect 12223 29214 12291 29270
rect 12347 29214 12415 29270
rect 12471 29214 12481 29270
rect 10669 29146 12481 29214
rect 10669 29090 10679 29146
rect 10735 29090 10803 29146
rect 10859 29090 10927 29146
rect 10983 29090 11051 29146
rect 11107 29090 11175 29146
rect 11231 29090 11299 29146
rect 11355 29090 11423 29146
rect 11479 29090 11547 29146
rect 11603 29090 11671 29146
rect 11727 29090 11795 29146
rect 11851 29090 11919 29146
rect 11975 29090 12043 29146
rect 12099 29090 12167 29146
rect 12223 29090 12291 29146
rect 12347 29090 12415 29146
rect 12471 29090 12481 29146
rect 10669 29022 12481 29090
rect 10669 28966 10679 29022
rect 10735 28966 10803 29022
rect 10859 28966 10927 29022
rect 10983 28966 11051 29022
rect 11107 28966 11175 29022
rect 11231 28966 11299 29022
rect 11355 28966 11423 29022
rect 11479 28966 11547 29022
rect 11603 28966 11671 29022
rect 11727 28966 11795 29022
rect 11851 28966 11919 29022
rect 11975 28966 12043 29022
rect 12099 28966 12167 29022
rect 12223 28966 12291 29022
rect 12347 28966 12415 29022
rect 12471 28966 12481 29022
rect 10669 28898 12481 28966
rect 10669 28842 10679 28898
rect 10735 28842 10803 28898
rect 10859 28842 10927 28898
rect 10983 28842 11051 28898
rect 11107 28842 11175 28898
rect 11231 28842 11299 28898
rect 11355 28842 11423 28898
rect 11479 28842 11547 28898
rect 11603 28842 11671 28898
rect 11727 28842 11795 28898
rect 11851 28842 11919 28898
rect 11975 28842 12043 28898
rect 12099 28842 12167 28898
rect 12223 28842 12291 28898
rect 12347 28842 12415 28898
rect 12471 28842 12481 28898
rect 10669 28832 12481 28842
rect 1489 28742 1499 28798
rect 1555 28742 1565 28798
rect 1489 28674 1565 28742
rect 1489 28618 1499 28674
rect 1555 28618 1565 28674
rect 1489 28550 1565 28618
rect 1489 28494 1499 28550
rect 1555 28494 1565 28550
rect 1489 28426 1565 28494
rect 1489 28370 1499 28426
rect 1555 28370 1565 28426
rect 1489 28302 1565 28370
rect 1489 28246 1499 28302
rect 1555 28246 1565 28302
rect 1489 28178 1565 28246
rect 1489 28122 1499 28178
rect 1555 28122 1565 28178
rect 1489 28054 1565 28122
rect 1489 27998 1499 28054
rect 1555 27998 1565 28054
rect 1489 27930 1565 27998
rect 1489 27874 1499 27930
rect 1555 27874 1565 27930
rect 1489 27806 1565 27874
rect 1489 27750 1499 27806
rect 1555 27750 1565 27806
rect 1489 27682 1565 27750
rect 1489 27626 1499 27682
rect 1555 27626 1565 27682
rect 1489 27558 1565 27626
rect 1489 27502 1499 27558
rect 1555 27502 1565 27558
rect 1489 27434 1565 27502
rect 1489 27378 1499 27434
rect 1555 27378 1565 27434
rect 1489 27310 1565 27378
rect 1489 27254 1499 27310
rect 1555 27254 1565 27310
rect 1613 28808 1689 28818
rect 1613 28752 1623 28808
rect 1679 28752 1689 28808
rect 1613 28684 1689 28752
rect 1613 28628 1623 28684
rect 1679 28628 1689 28684
rect 1613 28560 1689 28628
rect 1613 28504 1623 28560
rect 1679 28504 1689 28560
rect 1613 28436 1689 28504
rect 1613 28380 1623 28436
rect 1679 28380 1689 28436
rect 1613 28312 1689 28380
rect 1613 28256 1623 28312
rect 1679 28256 1689 28312
rect 1613 28188 1689 28256
rect 1613 28132 1623 28188
rect 1679 28132 1689 28188
rect 1613 28064 1689 28132
rect 1613 28008 1623 28064
rect 1679 28008 1689 28064
rect 1613 27940 1689 28008
rect 1613 27884 1623 27940
rect 1679 27884 1689 27940
rect 1613 27816 1689 27884
rect 1613 27760 1623 27816
rect 1679 27760 1689 27816
rect 1613 27692 1689 27760
rect 1613 27636 1623 27692
rect 1679 27636 1689 27692
rect 1613 27568 1689 27636
rect 1613 27512 1623 27568
rect 1679 27512 1689 27568
rect 1613 27444 1689 27512
rect 1613 27388 1623 27444
rect 1679 27388 1689 27444
rect 1613 27320 1689 27388
rect 1613 27264 1623 27320
rect 1679 27264 1689 27320
rect 1613 27254 1689 27264
rect 1737 28653 1813 28663
rect 1737 28597 1747 28653
rect 1803 28597 1813 28653
rect 1737 28529 1813 28597
rect 1737 28473 1747 28529
rect 1803 28473 1813 28529
rect 1737 28405 1813 28473
rect 1737 28349 1747 28405
rect 1803 28349 1813 28405
rect 1737 28281 1813 28349
rect 1737 28225 1747 28281
rect 1803 28225 1813 28281
rect 1737 28157 1813 28225
rect 1737 28101 1747 28157
rect 1803 28101 1813 28157
rect 1737 28033 1813 28101
rect 1737 27977 1747 28033
rect 1803 27977 1813 28033
rect 1737 27909 1813 27977
rect 1737 27853 1747 27909
rect 1803 27853 1813 27909
rect 1737 27785 1813 27853
rect 1737 27729 1747 27785
rect 1803 27729 1813 27785
rect 1737 27661 1813 27729
rect 1737 27605 1747 27661
rect 1803 27605 1813 27661
rect 1737 27537 1813 27605
rect 1737 27481 1747 27537
rect 1803 27481 1813 27537
rect 1737 27413 1813 27481
rect 1737 27357 1747 27413
rect 1803 27357 1813 27413
rect 1737 27289 1813 27357
rect 1489 27244 1565 27254
rect 1737 27233 1747 27289
rect 1803 27233 1813 27289
rect 1861 28539 1937 28549
rect 1861 28483 1871 28539
rect 1927 28483 1937 28539
rect 1861 28415 1937 28483
rect 1861 28359 1871 28415
rect 1927 28359 1937 28415
rect 1861 28291 1937 28359
rect 1861 28235 1871 28291
rect 1927 28235 1937 28291
rect 1861 28167 1937 28235
rect 1861 28111 1871 28167
rect 1927 28111 1937 28167
rect 1861 28043 1937 28111
rect 1861 27987 1871 28043
rect 1927 27987 1937 28043
rect 1861 27919 1937 27987
rect 1861 27863 1871 27919
rect 1927 27863 1937 27919
rect 1861 27795 1937 27863
rect 1861 27739 1871 27795
rect 1927 27739 1937 27795
rect 1861 27671 1937 27739
rect 1861 27615 1871 27671
rect 1927 27615 1937 27671
rect 1861 27547 1937 27615
rect 1861 27491 1871 27547
rect 1927 27491 1937 27547
rect 1861 27423 1937 27491
rect 1861 27367 1871 27423
rect 1927 27367 1937 27423
rect 1861 27299 1937 27367
rect 1861 27243 1871 27299
rect 1927 27243 1937 27299
rect 1861 27233 1937 27243
rect 1985 28537 2061 28547
rect 1985 28481 1995 28537
rect 2051 28481 2061 28537
rect 1985 28413 2061 28481
rect 1985 28357 1995 28413
rect 2051 28357 2061 28413
rect 1985 28289 2061 28357
rect 1985 28233 1995 28289
rect 2051 28233 2061 28289
rect 1985 28165 2061 28233
rect 1985 28109 1995 28165
rect 2051 28109 2061 28165
rect 1985 28041 2061 28109
rect 1985 27985 1995 28041
rect 2051 27985 2061 28041
rect 1985 27917 2061 27985
rect 1985 27861 1995 27917
rect 2051 27861 2061 27917
rect 1985 27793 2061 27861
rect 1985 27737 1995 27793
rect 2051 27737 2061 27793
rect 1985 27669 2061 27737
rect 1985 27613 1995 27669
rect 2051 27613 2061 27669
rect 1985 27545 2061 27613
rect 1985 27489 1995 27545
rect 2051 27489 2061 27545
rect 1985 27421 2061 27489
rect 1985 27365 1995 27421
rect 2051 27365 2061 27421
rect 1985 27297 2061 27365
rect 1985 27241 1995 27297
rect 2051 27241 2061 27297
rect 1737 27223 1813 27233
rect 1985 27231 2061 27241
rect 4425 28544 6237 28554
rect 4425 28488 4435 28544
rect 4491 28488 4559 28544
rect 4615 28488 4683 28544
rect 4739 28488 4807 28544
rect 4863 28488 4931 28544
rect 4987 28488 5055 28544
rect 5111 28488 5179 28544
rect 5235 28488 5303 28544
rect 5359 28488 5427 28544
rect 5483 28488 5551 28544
rect 5607 28488 5675 28544
rect 5731 28488 5799 28544
rect 5855 28488 5923 28544
rect 5979 28488 6047 28544
rect 6103 28488 6171 28544
rect 6227 28488 6237 28544
rect 4425 28420 6237 28488
rect 4425 28364 4435 28420
rect 4491 28364 4559 28420
rect 4615 28364 4683 28420
rect 4739 28364 4807 28420
rect 4863 28364 4931 28420
rect 4987 28364 5055 28420
rect 5111 28364 5179 28420
rect 5235 28364 5303 28420
rect 5359 28364 5427 28420
rect 5483 28364 5551 28420
rect 5607 28364 5675 28420
rect 5731 28364 5799 28420
rect 5855 28364 5923 28420
rect 5979 28364 6047 28420
rect 6103 28364 6171 28420
rect 6227 28364 6237 28420
rect 4425 28296 6237 28364
rect 4425 28240 4435 28296
rect 4491 28240 4559 28296
rect 4615 28240 4683 28296
rect 4739 28240 4807 28296
rect 4863 28240 4931 28296
rect 4987 28240 5055 28296
rect 5111 28240 5179 28296
rect 5235 28240 5303 28296
rect 5359 28240 5427 28296
rect 5483 28240 5551 28296
rect 5607 28240 5675 28296
rect 5731 28240 5799 28296
rect 5855 28240 5923 28296
rect 5979 28240 6047 28296
rect 6103 28240 6171 28296
rect 6227 28240 6237 28296
rect 4425 28172 6237 28240
rect 4425 28116 4435 28172
rect 4491 28116 4559 28172
rect 4615 28116 4683 28172
rect 4739 28116 4807 28172
rect 4863 28116 4931 28172
rect 4987 28116 5055 28172
rect 5111 28116 5179 28172
rect 5235 28116 5303 28172
rect 5359 28116 5427 28172
rect 5483 28116 5551 28172
rect 5607 28116 5675 28172
rect 5731 28116 5799 28172
rect 5855 28116 5923 28172
rect 5979 28116 6047 28172
rect 6103 28116 6171 28172
rect 6227 28116 6237 28172
rect 4425 28048 6237 28116
rect 4425 27992 4435 28048
rect 4491 27992 4559 28048
rect 4615 27992 4683 28048
rect 4739 27992 4807 28048
rect 4863 27992 4931 28048
rect 4987 27992 5055 28048
rect 5111 27992 5179 28048
rect 5235 27992 5303 28048
rect 5359 27992 5427 28048
rect 5483 27992 5551 28048
rect 5607 27992 5675 28048
rect 5731 27992 5799 28048
rect 5855 27992 5923 28048
rect 5979 27992 6047 28048
rect 6103 27992 6171 28048
rect 6227 27992 6237 28048
rect 4425 27924 6237 27992
rect 4425 27868 4435 27924
rect 4491 27868 4559 27924
rect 4615 27868 4683 27924
rect 4739 27868 4807 27924
rect 4863 27868 4931 27924
rect 4987 27868 5055 27924
rect 5111 27868 5179 27924
rect 5235 27868 5303 27924
rect 5359 27868 5427 27924
rect 5483 27868 5551 27924
rect 5607 27868 5675 27924
rect 5731 27868 5799 27924
rect 5855 27868 5923 27924
rect 5979 27868 6047 27924
rect 6103 27868 6171 27924
rect 6227 27868 6237 27924
rect 4425 27800 6237 27868
rect 4425 27744 4435 27800
rect 4491 27744 4559 27800
rect 4615 27744 4683 27800
rect 4739 27744 4807 27800
rect 4863 27744 4931 27800
rect 4987 27744 5055 27800
rect 5111 27744 5179 27800
rect 5235 27744 5303 27800
rect 5359 27744 5427 27800
rect 5483 27744 5551 27800
rect 5607 27744 5675 27800
rect 5731 27744 5799 27800
rect 5855 27744 5923 27800
rect 5979 27744 6047 27800
rect 6103 27744 6171 27800
rect 6227 27744 6237 27800
rect 4425 27676 6237 27744
rect 4425 27620 4435 27676
rect 4491 27620 4559 27676
rect 4615 27620 4683 27676
rect 4739 27620 4807 27676
rect 4863 27620 4931 27676
rect 4987 27620 5055 27676
rect 5111 27620 5179 27676
rect 5235 27620 5303 27676
rect 5359 27620 5427 27676
rect 5483 27620 5551 27676
rect 5607 27620 5675 27676
rect 5731 27620 5799 27676
rect 5855 27620 5923 27676
rect 5979 27620 6047 27676
rect 6103 27620 6171 27676
rect 6227 27620 6237 27676
rect 4425 27552 6237 27620
rect 4425 27496 4435 27552
rect 4491 27496 4559 27552
rect 4615 27496 4683 27552
rect 4739 27496 4807 27552
rect 4863 27496 4931 27552
rect 4987 27496 5055 27552
rect 5111 27496 5179 27552
rect 5235 27496 5303 27552
rect 5359 27496 5427 27552
rect 5483 27496 5551 27552
rect 5607 27496 5675 27552
rect 5731 27496 5799 27552
rect 5855 27496 5923 27552
rect 5979 27496 6047 27552
rect 6103 27496 6171 27552
rect 6227 27496 6237 27552
rect 4425 27428 6237 27496
rect 4425 27372 4435 27428
rect 4491 27372 4559 27428
rect 4615 27372 4683 27428
rect 4739 27372 4807 27428
rect 4863 27372 4931 27428
rect 4987 27372 5055 27428
rect 5111 27372 5179 27428
rect 5235 27372 5303 27428
rect 5359 27372 5427 27428
rect 5483 27372 5551 27428
rect 5607 27372 5675 27428
rect 5731 27372 5799 27428
rect 5855 27372 5923 27428
rect 5979 27372 6047 27428
rect 6103 27372 6171 27428
rect 6227 27372 6237 27428
rect 4425 27304 6237 27372
rect 4425 27248 4435 27304
rect 4491 27248 4559 27304
rect 4615 27248 4683 27304
rect 4739 27248 4807 27304
rect 4863 27248 4931 27304
rect 4987 27248 5055 27304
rect 5111 27248 5179 27304
rect 5235 27248 5303 27304
rect 5359 27248 5427 27304
rect 5483 27248 5551 27304
rect 5607 27248 5675 27304
rect 5731 27248 5799 27304
rect 5855 27248 5923 27304
rect 5979 27248 6047 27304
rect 6103 27248 6171 27304
rect 6227 27248 6237 27304
rect 4425 27238 6237 27248
rect 7552 28544 8620 28554
rect 7552 28488 7562 28544
rect 7618 28488 7686 28544
rect 7742 28488 7810 28544
rect 7866 28488 7934 28544
rect 7990 28488 8058 28544
rect 8114 28488 8182 28544
rect 8238 28488 8306 28544
rect 8362 28488 8430 28544
rect 8486 28488 8554 28544
rect 8610 28488 8620 28544
rect 7552 28420 8620 28488
rect 7552 28364 7562 28420
rect 7618 28364 7686 28420
rect 7742 28364 7810 28420
rect 7866 28364 7934 28420
rect 7990 28364 8058 28420
rect 8114 28364 8182 28420
rect 8238 28364 8306 28420
rect 8362 28364 8430 28420
rect 8486 28364 8554 28420
rect 8610 28364 8620 28420
rect 7552 28296 8620 28364
rect 7552 28240 7562 28296
rect 7618 28240 7686 28296
rect 7742 28240 7810 28296
rect 7866 28240 7934 28296
rect 7990 28240 8058 28296
rect 8114 28240 8182 28296
rect 8238 28240 8306 28296
rect 8362 28240 8430 28296
rect 8486 28240 8554 28296
rect 8610 28240 8620 28296
rect 7552 28172 8620 28240
rect 7552 28116 7562 28172
rect 7618 28116 7686 28172
rect 7742 28116 7810 28172
rect 7866 28116 7934 28172
rect 7990 28116 8058 28172
rect 8114 28116 8182 28172
rect 8238 28116 8306 28172
rect 8362 28116 8430 28172
rect 8486 28116 8554 28172
rect 8610 28116 8620 28172
rect 7552 28048 8620 28116
rect 7552 27992 7562 28048
rect 7618 27992 7686 28048
rect 7742 27992 7810 28048
rect 7866 27992 7934 28048
rect 7990 27992 8058 28048
rect 8114 27992 8182 28048
rect 8238 27992 8306 28048
rect 8362 27992 8430 28048
rect 8486 27992 8554 28048
rect 8610 27992 8620 28048
rect 7552 27924 8620 27992
rect 7552 27868 7562 27924
rect 7618 27868 7686 27924
rect 7742 27868 7810 27924
rect 7866 27868 7934 27924
rect 7990 27868 8058 27924
rect 8114 27868 8182 27924
rect 8238 27868 8306 27924
rect 8362 27868 8430 27924
rect 8486 27868 8554 27924
rect 8610 27868 8620 27924
rect 7552 27800 8620 27868
rect 7552 27744 7562 27800
rect 7618 27744 7686 27800
rect 7742 27744 7810 27800
rect 7866 27744 7934 27800
rect 7990 27744 8058 27800
rect 8114 27744 8182 27800
rect 8238 27744 8306 27800
rect 8362 27744 8430 27800
rect 8486 27744 8554 27800
rect 8610 27744 8620 27800
rect 7552 27676 8620 27744
rect 7552 27620 7562 27676
rect 7618 27620 7686 27676
rect 7742 27620 7810 27676
rect 7866 27620 7934 27676
rect 7990 27620 8058 27676
rect 8114 27620 8182 27676
rect 8238 27620 8306 27676
rect 8362 27620 8430 27676
rect 8486 27620 8554 27676
rect 8610 27620 8620 27676
rect 7552 27552 8620 27620
rect 7552 27496 7562 27552
rect 7618 27496 7686 27552
rect 7742 27496 7810 27552
rect 7866 27496 7934 27552
rect 7990 27496 8058 27552
rect 8114 27496 8182 27552
rect 8238 27496 8306 27552
rect 8362 27496 8430 27552
rect 8486 27496 8554 27552
rect 8610 27496 8620 27552
rect 7552 27428 8620 27496
rect 7552 27372 7562 27428
rect 7618 27372 7686 27428
rect 7742 27372 7810 27428
rect 7866 27372 7934 27428
rect 7990 27372 8058 27428
rect 8114 27372 8182 27428
rect 8238 27372 8306 27428
rect 8362 27372 8430 27428
rect 8486 27372 8554 27428
rect 8610 27372 8620 27428
rect 7552 27304 8620 27372
rect 7552 27248 7562 27304
rect 7618 27248 7686 27304
rect 7742 27248 7810 27304
rect 7866 27248 7934 27304
rect 7990 27248 8058 27304
rect 8114 27248 8182 27304
rect 8238 27248 8306 27304
rect 8362 27248 8430 27304
rect 8486 27248 8554 27304
rect 8610 27248 8620 27304
rect 7552 27238 8620 27248
rect 10669 28544 12481 28554
rect 10669 28488 10679 28544
rect 10735 28488 10803 28544
rect 10859 28488 10927 28544
rect 10983 28488 11051 28544
rect 11107 28488 11175 28544
rect 11231 28488 11299 28544
rect 11355 28488 11423 28544
rect 11479 28488 11547 28544
rect 11603 28488 11671 28544
rect 11727 28488 11795 28544
rect 11851 28488 11919 28544
rect 11975 28488 12043 28544
rect 12099 28488 12167 28544
rect 12223 28488 12291 28544
rect 12347 28488 12415 28544
rect 12471 28488 12481 28544
rect 10669 28420 12481 28488
rect 10669 28364 10679 28420
rect 10735 28364 10803 28420
rect 10859 28364 10927 28420
rect 10983 28364 11051 28420
rect 11107 28364 11175 28420
rect 11231 28364 11299 28420
rect 11355 28364 11423 28420
rect 11479 28364 11547 28420
rect 11603 28364 11671 28420
rect 11727 28364 11795 28420
rect 11851 28364 11919 28420
rect 11975 28364 12043 28420
rect 12099 28364 12167 28420
rect 12223 28364 12291 28420
rect 12347 28364 12415 28420
rect 12471 28364 12481 28420
rect 10669 28296 12481 28364
rect 10669 28240 10679 28296
rect 10735 28240 10803 28296
rect 10859 28240 10927 28296
rect 10983 28240 11051 28296
rect 11107 28240 11175 28296
rect 11231 28240 11299 28296
rect 11355 28240 11423 28296
rect 11479 28240 11547 28296
rect 11603 28240 11671 28296
rect 11727 28240 11795 28296
rect 11851 28240 11919 28296
rect 11975 28240 12043 28296
rect 12099 28240 12167 28296
rect 12223 28240 12291 28296
rect 12347 28240 12415 28296
rect 12471 28240 12481 28296
rect 10669 28172 12481 28240
rect 10669 28116 10679 28172
rect 10735 28116 10803 28172
rect 10859 28116 10927 28172
rect 10983 28116 11051 28172
rect 11107 28116 11175 28172
rect 11231 28116 11299 28172
rect 11355 28116 11423 28172
rect 11479 28116 11547 28172
rect 11603 28116 11671 28172
rect 11727 28116 11795 28172
rect 11851 28116 11919 28172
rect 11975 28116 12043 28172
rect 12099 28116 12167 28172
rect 12223 28116 12291 28172
rect 12347 28116 12415 28172
rect 12471 28116 12481 28172
rect 10669 28048 12481 28116
rect 10669 27992 10679 28048
rect 10735 27992 10803 28048
rect 10859 27992 10927 28048
rect 10983 27992 11051 28048
rect 11107 27992 11175 28048
rect 11231 27992 11299 28048
rect 11355 27992 11423 28048
rect 11479 27992 11547 28048
rect 11603 27992 11671 28048
rect 11727 27992 11795 28048
rect 11851 27992 11919 28048
rect 11975 27992 12043 28048
rect 12099 27992 12167 28048
rect 12223 27992 12291 28048
rect 12347 27992 12415 28048
rect 12471 27992 12481 28048
rect 10669 27924 12481 27992
rect 10669 27868 10679 27924
rect 10735 27868 10803 27924
rect 10859 27868 10927 27924
rect 10983 27868 11051 27924
rect 11107 27868 11175 27924
rect 11231 27868 11299 27924
rect 11355 27868 11423 27924
rect 11479 27868 11547 27924
rect 11603 27868 11671 27924
rect 11727 27868 11795 27924
rect 11851 27868 11919 27924
rect 11975 27868 12043 27924
rect 12099 27868 12167 27924
rect 12223 27868 12291 27924
rect 12347 27868 12415 27924
rect 12471 27868 12481 27924
rect 10669 27800 12481 27868
rect 10669 27744 10679 27800
rect 10735 27744 10803 27800
rect 10859 27744 10927 27800
rect 10983 27744 11051 27800
rect 11107 27744 11175 27800
rect 11231 27744 11299 27800
rect 11355 27744 11423 27800
rect 11479 27744 11547 27800
rect 11603 27744 11671 27800
rect 11727 27744 11795 27800
rect 11851 27744 11919 27800
rect 11975 27744 12043 27800
rect 12099 27744 12167 27800
rect 12223 27744 12291 27800
rect 12347 27744 12415 27800
rect 12471 27744 12481 27800
rect 10669 27676 12481 27744
rect 10669 27620 10679 27676
rect 10735 27620 10803 27676
rect 10859 27620 10927 27676
rect 10983 27620 11051 27676
rect 11107 27620 11175 27676
rect 11231 27620 11299 27676
rect 11355 27620 11423 27676
rect 11479 27620 11547 27676
rect 11603 27620 11671 27676
rect 11727 27620 11795 27676
rect 11851 27620 11919 27676
rect 11975 27620 12043 27676
rect 12099 27620 12167 27676
rect 12223 27620 12291 27676
rect 12347 27620 12415 27676
rect 12471 27620 12481 27676
rect 10669 27552 12481 27620
rect 10669 27496 10679 27552
rect 10735 27496 10803 27552
rect 10859 27496 10927 27552
rect 10983 27496 11051 27552
rect 11107 27496 11175 27552
rect 11231 27496 11299 27552
rect 11355 27496 11423 27552
rect 11479 27496 11547 27552
rect 11603 27496 11671 27552
rect 11727 27496 11795 27552
rect 11851 27496 11919 27552
rect 11975 27496 12043 27552
rect 12099 27496 12167 27552
rect 12223 27496 12291 27552
rect 12347 27496 12415 27552
rect 12471 27496 12481 27552
rect 10669 27428 12481 27496
rect 10669 27372 10679 27428
rect 10735 27372 10803 27428
rect 10859 27372 10927 27428
rect 10983 27372 11051 27428
rect 11107 27372 11175 27428
rect 11231 27372 11299 27428
rect 11355 27372 11423 27428
rect 11479 27372 11547 27428
rect 11603 27372 11671 27428
rect 11727 27372 11795 27428
rect 11851 27372 11919 27428
rect 11975 27372 12043 27428
rect 12099 27372 12167 27428
rect 12223 27372 12291 27428
rect 12347 27372 12415 27428
rect 12471 27372 12481 27428
rect 10669 27304 12481 27372
rect 10669 27248 10679 27304
rect 10735 27248 10803 27304
rect 10859 27248 10927 27304
rect 10983 27248 11051 27304
rect 11107 27248 11175 27304
rect 11231 27248 11299 27304
rect 11355 27248 11423 27304
rect 11479 27248 11547 27304
rect 11603 27248 11671 27304
rect 11727 27248 11795 27304
rect 11851 27248 11919 27304
rect 11975 27248 12043 27304
rect 12099 27248 12167 27304
rect 12223 27248 12291 27304
rect 12347 27248 12415 27304
rect 12471 27248 12481 27304
rect 10669 27238 12481 27248
rect 2497 26944 4309 26954
rect 2497 26888 2507 26944
rect 2563 26888 2631 26944
rect 2687 26888 2755 26944
rect 2811 26888 2879 26944
rect 2935 26888 3003 26944
rect 3059 26888 3127 26944
rect 3183 26888 3251 26944
rect 3307 26888 3375 26944
rect 3431 26888 3499 26944
rect 3555 26888 3623 26944
rect 3679 26888 3747 26944
rect 3803 26888 3871 26944
rect 3927 26888 3995 26944
rect 4051 26888 4119 26944
rect 4175 26888 4243 26944
rect 4299 26888 4309 26944
rect 2497 26820 4309 26888
rect 2497 26764 2507 26820
rect 2563 26764 2631 26820
rect 2687 26764 2755 26820
rect 2811 26764 2879 26820
rect 2935 26764 3003 26820
rect 3059 26764 3127 26820
rect 3183 26764 3251 26820
rect 3307 26764 3375 26820
rect 3431 26764 3499 26820
rect 3555 26764 3623 26820
rect 3679 26764 3747 26820
rect 3803 26764 3871 26820
rect 3927 26764 3995 26820
rect 4051 26764 4119 26820
rect 4175 26764 4243 26820
rect 4299 26764 4309 26820
rect 2497 26696 4309 26764
rect 2497 26640 2507 26696
rect 2563 26640 2631 26696
rect 2687 26640 2755 26696
rect 2811 26640 2879 26696
rect 2935 26640 3003 26696
rect 3059 26640 3127 26696
rect 3183 26640 3251 26696
rect 3307 26640 3375 26696
rect 3431 26640 3499 26696
rect 3555 26640 3623 26696
rect 3679 26640 3747 26696
rect 3803 26640 3871 26696
rect 3927 26640 3995 26696
rect 4051 26640 4119 26696
rect 4175 26640 4243 26696
rect 4299 26640 4309 26696
rect 2497 26572 4309 26640
rect 2497 26516 2507 26572
rect 2563 26516 2631 26572
rect 2687 26516 2755 26572
rect 2811 26516 2879 26572
rect 2935 26516 3003 26572
rect 3059 26516 3127 26572
rect 3183 26516 3251 26572
rect 3307 26516 3375 26572
rect 3431 26516 3499 26572
rect 3555 26516 3623 26572
rect 3679 26516 3747 26572
rect 3803 26516 3871 26572
rect 3927 26516 3995 26572
rect 4051 26516 4119 26572
rect 4175 26516 4243 26572
rect 4299 26516 4309 26572
rect 2497 26448 4309 26516
rect 2497 26392 2507 26448
rect 2563 26392 2631 26448
rect 2687 26392 2755 26448
rect 2811 26392 2879 26448
rect 2935 26392 3003 26448
rect 3059 26392 3127 26448
rect 3183 26392 3251 26448
rect 3307 26392 3375 26448
rect 3431 26392 3499 26448
rect 3555 26392 3623 26448
rect 3679 26392 3747 26448
rect 3803 26392 3871 26448
rect 3927 26392 3995 26448
rect 4051 26392 4119 26448
rect 4175 26392 4243 26448
rect 4299 26392 4309 26448
rect 2497 26324 4309 26392
rect 2497 26268 2507 26324
rect 2563 26268 2631 26324
rect 2687 26268 2755 26324
rect 2811 26268 2879 26324
rect 2935 26268 3003 26324
rect 3059 26268 3127 26324
rect 3183 26268 3251 26324
rect 3307 26268 3375 26324
rect 3431 26268 3499 26324
rect 3555 26268 3623 26324
rect 3679 26268 3747 26324
rect 3803 26268 3871 26324
rect 3927 26268 3995 26324
rect 4051 26268 4119 26324
rect 4175 26268 4243 26324
rect 4299 26268 4309 26324
rect 2497 26200 4309 26268
rect 2497 26144 2507 26200
rect 2563 26144 2631 26200
rect 2687 26144 2755 26200
rect 2811 26144 2879 26200
rect 2935 26144 3003 26200
rect 3059 26144 3127 26200
rect 3183 26144 3251 26200
rect 3307 26144 3375 26200
rect 3431 26144 3499 26200
rect 3555 26144 3623 26200
rect 3679 26144 3747 26200
rect 3803 26144 3871 26200
rect 3927 26144 3995 26200
rect 4051 26144 4119 26200
rect 4175 26144 4243 26200
rect 4299 26144 4309 26200
rect 2497 26076 4309 26144
rect 2497 26020 2507 26076
rect 2563 26020 2631 26076
rect 2687 26020 2755 26076
rect 2811 26020 2879 26076
rect 2935 26020 3003 26076
rect 3059 26020 3127 26076
rect 3183 26020 3251 26076
rect 3307 26020 3375 26076
rect 3431 26020 3499 26076
rect 3555 26020 3623 26076
rect 3679 26020 3747 26076
rect 3803 26020 3871 26076
rect 3927 26020 3995 26076
rect 4051 26020 4119 26076
rect 4175 26020 4243 26076
rect 4299 26020 4309 26076
rect 2497 25952 4309 26020
rect 2497 25896 2507 25952
rect 2563 25896 2631 25952
rect 2687 25896 2755 25952
rect 2811 25896 2879 25952
rect 2935 25896 3003 25952
rect 3059 25896 3127 25952
rect 3183 25896 3251 25952
rect 3307 25896 3375 25952
rect 3431 25896 3499 25952
rect 3555 25896 3623 25952
rect 3679 25896 3747 25952
rect 3803 25896 3871 25952
rect 3927 25896 3995 25952
rect 4051 25896 4119 25952
rect 4175 25896 4243 25952
rect 4299 25896 4309 25952
rect 2497 25828 4309 25896
rect 2497 25772 2507 25828
rect 2563 25772 2631 25828
rect 2687 25772 2755 25828
rect 2811 25772 2879 25828
rect 2935 25772 3003 25828
rect 3059 25772 3127 25828
rect 3183 25772 3251 25828
rect 3307 25772 3375 25828
rect 3431 25772 3499 25828
rect 3555 25772 3623 25828
rect 3679 25772 3747 25828
rect 3803 25772 3871 25828
rect 3927 25772 3995 25828
rect 4051 25772 4119 25828
rect 4175 25772 4243 25828
rect 4299 25772 4309 25828
rect 2497 25704 4309 25772
rect 2497 25648 2507 25704
rect 2563 25648 2631 25704
rect 2687 25648 2755 25704
rect 2811 25648 2879 25704
rect 2935 25648 3003 25704
rect 3059 25648 3127 25704
rect 3183 25648 3251 25704
rect 3307 25648 3375 25704
rect 3431 25648 3499 25704
rect 3555 25648 3623 25704
rect 3679 25648 3747 25704
rect 3803 25648 3871 25704
rect 3927 25648 3995 25704
rect 4051 25648 4119 25704
rect 4175 25648 4243 25704
rect 4299 25648 4309 25704
rect 2497 25638 4309 25648
rect 6358 26944 7426 26954
rect 6358 26888 6368 26944
rect 6424 26888 6492 26944
rect 6548 26888 6616 26944
rect 6672 26888 6740 26944
rect 6796 26888 6864 26944
rect 6920 26888 6988 26944
rect 7044 26888 7112 26944
rect 7168 26888 7236 26944
rect 7292 26888 7360 26944
rect 7416 26888 7426 26944
rect 6358 26820 7426 26888
rect 6358 26764 6368 26820
rect 6424 26764 6492 26820
rect 6548 26764 6616 26820
rect 6672 26764 6740 26820
rect 6796 26764 6864 26820
rect 6920 26764 6988 26820
rect 7044 26764 7112 26820
rect 7168 26764 7236 26820
rect 7292 26764 7360 26820
rect 7416 26764 7426 26820
rect 6358 26696 7426 26764
rect 6358 26640 6368 26696
rect 6424 26640 6492 26696
rect 6548 26640 6616 26696
rect 6672 26640 6740 26696
rect 6796 26640 6864 26696
rect 6920 26640 6988 26696
rect 7044 26640 7112 26696
rect 7168 26640 7236 26696
rect 7292 26640 7360 26696
rect 7416 26640 7426 26696
rect 6358 26572 7426 26640
rect 6358 26516 6368 26572
rect 6424 26516 6492 26572
rect 6548 26516 6616 26572
rect 6672 26516 6740 26572
rect 6796 26516 6864 26572
rect 6920 26516 6988 26572
rect 7044 26516 7112 26572
rect 7168 26516 7236 26572
rect 7292 26516 7360 26572
rect 7416 26516 7426 26572
rect 6358 26448 7426 26516
rect 6358 26392 6368 26448
rect 6424 26392 6492 26448
rect 6548 26392 6616 26448
rect 6672 26392 6740 26448
rect 6796 26392 6864 26448
rect 6920 26392 6988 26448
rect 7044 26392 7112 26448
rect 7168 26392 7236 26448
rect 7292 26392 7360 26448
rect 7416 26392 7426 26448
rect 6358 26324 7426 26392
rect 6358 26268 6368 26324
rect 6424 26268 6492 26324
rect 6548 26268 6616 26324
rect 6672 26268 6740 26324
rect 6796 26268 6864 26324
rect 6920 26268 6988 26324
rect 7044 26268 7112 26324
rect 7168 26268 7236 26324
rect 7292 26268 7360 26324
rect 7416 26268 7426 26324
rect 6358 26200 7426 26268
rect 6358 26144 6368 26200
rect 6424 26144 6492 26200
rect 6548 26144 6616 26200
rect 6672 26144 6740 26200
rect 6796 26144 6864 26200
rect 6920 26144 6988 26200
rect 7044 26144 7112 26200
rect 7168 26144 7236 26200
rect 7292 26144 7360 26200
rect 7416 26144 7426 26200
rect 6358 26076 7426 26144
rect 6358 26020 6368 26076
rect 6424 26020 6492 26076
rect 6548 26020 6616 26076
rect 6672 26020 6740 26076
rect 6796 26020 6864 26076
rect 6920 26020 6988 26076
rect 7044 26020 7112 26076
rect 7168 26020 7236 26076
rect 7292 26020 7360 26076
rect 7416 26020 7426 26076
rect 6358 25952 7426 26020
rect 6358 25896 6368 25952
rect 6424 25896 6492 25952
rect 6548 25896 6616 25952
rect 6672 25896 6740 25952
rect 6796 25896 6864 25952
rect 6920 25896 6988 25952
rect 7044 25896 7112 25952
rect 7168 25896 7236 25952
rect 7292 25896 7360 25952
rect 7416 25896 7426 25952
rect 6358 25828 7426 25896
rect 6358 25772 6368 25828
rect 6424 25772 6492 25828
rect 6548 25772 6616 25828
rect 6672 25772 6740 25828
rect 6796 25772 6864 25828
rect 6920 25772 6988 25828
rect 7044 25772 7112 25828
rect 7168 25772 7236 25828
rect 7292 25772 7360 25828
rect 7416 25772 7426 25828
rect 6358 25704 7426 25772
rect 6358 25648 6368 25704
rect 6424 25648 6492 25704
rect 6548 25648 6616 25704
rect 6672 25648 6740 25704
rect 6796 25648 6864 25704
rect 6920 25648 6988 25704
rect 7044 25648 7112 25704
rect 7168 25648 7236 25704
rect 7292 25648 7360 25704
rect 7416 25648 7426 25704
rect 6358 25638 7426 25648
rect 8741 26944 10553 26954
rect 8741 26888 8751 26944
rect 8807 26888 8875 26944
rect 8931 26888 8999 26944
rect 9055 26888 9123 26944
rect 9179 26888 9247 26944
rect 9303 26888 9371 26944
rect 9427 26888 9495 26944
rect 9551 26888 9619 26944
rect 9675 26888 9743 26944
rect 9799 26888 9867 26944
rect 9923 26888 9991 26944
rect 10047 26888 10115 26944
rect 10171 26888 10239 26944
rect 10295 26888 10363 26944
rect 10419 26888 10487 26944
rect 10543 26888 10553 26944
rect 8741 26820 10553 26888
rect 8741 26764 8751 26820
rect 8807 26764 8875 26820
rect 8931 26764 8999 26820
rect 9055 26764 9123 26820
rect 9179 26764 9247 26820
rect 9303 26764 9371 26820
rect 9427 26764 9495 26820
rect 9551 26764 9619 26820
rect 9675 26764 9743 26820
rect 9799 26764 9867 26820
rect 9923 26764 9991 26820
rect 10047 26764 10115 26820
rect 10171 26764 10239 26820
rect 10295 26764 10363 26820
rect 10419 26764 10487 26820
rect 10543 26764 10553 26820
rect 8741 26696 10553 26764
rect 8741 26640 8751 26696
rect 8807 26640 8875 26696
rect 8931 26640 8999 26696
rect 9055 26640 9123 26696
rect 9179 26640 9247 26696
rect 9303 26640 9371 26696
rect 9427 26640 9495 26696
rect 9551 26640 9619 26696
rect 9675 26640 9743 26696
rect 9799 26640 9867 26696
rect 9923 26640 9991 26696
rect 10047 26640 10115 26696
rect 10171 26640 10239 26696
rect 10295 26640 10363 26696
rect 10419 26640 10487 26696
rect 10543 26640 10553 26696
rect 8741 26572 10553 26640
rect 8741 26516 8751 26572
rect 8807 26516 8875 26572
rect 8931 26516 8999 26572
rect 9055 26516 9123 26572
rect 9179 26516 9247 26572
rect 9303 26516 9371 26572
rect 9427 26516 9495 26572
rect 9551 26516 9619 26572
rect 9675 26516 9743 26572
rect 9799 26516 9867 26572
rect 9923 26516 9991 26572
rect 10047 26516 10115 26572
rect 10171 26516 10239 26572
rect 10295 26516 10363 26572
rect 10419 26516 10487 26572
rect 10543 26516 10553 26572
rect 8741 26448 10553 26516
rect 8741 26392 8751 26448
rect 8807 26392 8875 26448
rect 8931 26392 8999 26448
rect 9055 26392 9123 26448
rect 9179 26392 9247 26448
rect 9303 26392 9371 26448
rect 9427 26392 9495 26448
rect 9551 26392 9619 26448
rect 9675 26392 9743 26448
rect 9799 26392 9867 26448
rect 9923 26392 9991 26448
rect 10047 26392 10115 26448
rect 10171 26392 10239 26448
rect 10295 26392 10363 26448
rect 10419 26392 10487 26448
rect 10543 26392 10553 26448
rect 8741 26324 10553 26392
rect 8741 26268 8751 26324
rect 8807 26268 8875 26324
rect 8931 26268 8999 26324
rect 9055 26268 9123 26324
rect 9179 26268 9247 26324
rect 9303 26268 9371 26324
rect 9427 26268 9495 26324
rect 9551 26268 9619 26324
rect 9675 26268 9743 26324
rect 9799 26268 9867 26324
rect 9923 26268 9991 26324
rect 10047 26268 10115 26324
rect 10171 26268 10239 26324
rect 10295 26268 10363 26324
rect 10419 26268 10487 26324
rect 10543 26268 10553 26324
rect 8741 26200 10553 26268
rect 8741 26144 8751 26200
rect 8807 26144 8875 26200
rect 8931 26144 8999 26200
rect 9055 26144 9123 26200
rect 9179 26144 9247 26200
rect 9303 26144 9371 26200
rect 9427 26144 9495 26200
rect 9551 26144 9619 26200
rect 9675 26144 9743 26200
rect 9799 26144 9867 26200
rect 9923 26144 9991 26200
rect 10047 26144 10115 26200
rect 10171 26144 10239 26200
rect 10295 26144 10363 26200
rect 10419 26144 10487 26200
rect 10543 26144 10553 26200
rect 8741 26076 10553 26144
rect 8741 26020 8751 26076
rect 8807 26020 8875 26076
rect 8931 26020 8999 26076
rect 9055 26020 9123 26076
rect 9179 26020 9247 26076
rect 9303 26020 9371 26076
rect 9427 26020 9495 26076
rect 9551 26020 9619 26076
rect 9675 26020 9743 26076
rect 9799 26020 9867 26076
rect 9923 26020 9991 26076
rect 10047 26020 10115 26076
rect 10171 26020 10239 26076
rect 10295 26020 10363 26076
rect 10419 26020 10487 26076
rect 10543 26020 10553 26076
rect 8741 25952 10553 26020
rect 8741 25896 8751 25952
rect 8807 25896 8875 25952
rect 8931 25896 8999 25952
rect 9055 25896 9123 25952
rect 9179 25896 9247 25952
rect 9303 25896 9371 25952
rect 9427 25896 9495 25952
rect 9551 25896 9619 25952
rect 9675 25896 9743 25952
rect 9799 25896 9867 25952
rect 9923 25896 9991 25952
rect 10047 25896 10115 25952
rect 10171 25896 10239 25952
rect 10295 25896 10363 25952
rect 10419 25896 10487 25952
rect 10543 25896 10553 25952
rect 8741 25828 10553 25896
rect 8741 25772 8751 25828
rect 8807 25772 8875 25828
rect 8931 25772 8999 25828
rect 9055 25772 9123 25828
rect 9179 25772 9247 25828
rect 9303 25772 9371 25828
rect 9427 25772 9495 25828
rect 9551 25772 9619 25828
rect 9675 25772 9743 25828
rect 9799 25772 9867 25828
rect 9923 25772 9991 25828
rect 10047 25772 10115 25828
rect 10171 25772 10239 25828
rect 10295 25772 10363 25828
rect 10419 25772 10487 25828
rect 10543 25772 10553 25828
rect 8741 25704 10553 25772
rect 8741 25648 8751 25704
rect 8807 25648 8875 25704
rect 8931 25648 8999 25704
rect 9055 25648 9123 25704
rect 9179 25648 9247 25704
rect 9303 25648 9371 25704
rect 9427 25648 9495 25704
rect 9551 25648 9619 25704
rect 9675 25648 9743 25704
rect 9799 25648 9867 25704
rect 9923 25648 9991 25704
rect 10047 25648 10115 25704
rect 10171 25648 10239 25704
rect 10295 25648 10363 25704
rect 10419 25648 10487 25704
rect 10543 25648 10553 25704
rect 8741 25638 10553 25648
rect 12842 26944 13910 26954
rect 12842 26888 12852 26944
rect 12908 26888 12976 26944
rect 13032 26888 13100 26944
rect 13156 26888 13224 26944
rect 13280 26888 13348 26944
rect 13404 26888 13472 26944
rect 13528 26888 13596 26944
rect 13652 26888 13720 26944
rect 13776 26888 13844 26944
rect 13900 26888 13910 26944
rect 12842 26820 13910 26888
rect 12842 26764 12852 26820
rect 12908 26764 12976 26820
rect 13032 26764 13100 26820
rect 13156 26764 13224 26820
rect 13280 26764 13348 26820
rect 13404 26764 13472 26820
rect 13528 26764 13596 26820
rect 13652 26764 13720 26820
rect 13776 26764 13844 26820
rect 13900 26764 13910 26820
rect 12842 26696 13910 26764
rect 12842 26640 12852 26696
rect 12908 26640 12976 26696
rect 13032 26640 13100 26696
rect 13156 26640 13224 26696
rect 13280 26640 13348 26696
rect 13404 26640 13472 26696
rect 13528 26640 13596 26696
rect 13652 26640 13720 26696
rect 13776 26640 13844 26696
rect 13900 26640 13910 26696
rect 12842 26572 13910 26640
rect 12842 26516 12852 26572
rect 12908 26516 12976 26572
rect 13032 26516 13100 26572
rect 13156 26516 13224 26572
rect 13280 26516 13348 26572
rect 13404 26516 13472 26572
rect 13528 26516 13596 26572
rect 13652 26516 13720 26572
rect 13776 26516 13844 26572
rect 13900 26516 13910 26572
rect 12842 26448 13910 26516
rect 12842 26392 12852 26448
rect 12908 26392 12976 26448
rect 13032 26392 13100 26448
rect 13156 26392 13224 26448
rect 13280 26392 13348 26448
rect 13404 26392 13472 26448
rect 13528 26392 13596 26448
rect 13652 26392 13720 26448
rect 13776 26392 13844 26448
rect 13900 26392 13910 26448
rect 12842 26324 13910 26392
rect 12842 26268 12852 26324
rect 12908 26268 12976 26324
rect 13032 26268 13100 26324
rect 13156 26268 13224 26324
rect 13280 26268 13348 26324
rect 13404 26268 13472 26324
rect 13528 26268 13596 26324
rect 13652 26268 13720 26324
rect 13776 26268 13844 26324
rect 13900 26268 13910 26324
rect 12842 26200 13910 26268
rect 12842 26144 12852 26200
rect 12908 26144 12976 26200
rect 13032 26144 13100 26200
rect 13156 26144 13224 26200
rect 13280 26144 13348 26200
rect 13404 26144 13472 26200
rect 13528 26144 13596 26200
rect 13652 26144 13720 26200
rect 13776 26144 13844 26200
rect 13900 26144 13910 26200
rect 12842 26076 13910 26144
rect 12842 26020 12852 26076
rect 12908 26020 12976 26076
rect 13032 26020 13100 26076
rect 13156 26020 13224 26076
rect 13280 26020 13348 26076
rect 13404 26020 13472 26076
rect 13528 26020 13596 26076
rect 13652 26020 13720 26076
rect 13776 26020 13844 26076
rect 13900 26020 13910 26076
rect 12842 25952 13910 26020
rect 12842 25896 12852 25952
rect 12908 25896 12976 25952
rect 13032 25896 13100 25952
rect 13156 25896 13224 25952
rect 13280 25896 13348 25952
rect 13404 25896 13472 25952
rect 13528 25896 13596 25952
rect 13652 25896 13720 25952
rect 13776 25896 13844 25952
rect 13900 25896 13910 25952
rect 12842 25828 13910 25896
rect 12842 25772 12852 25828
rect 12908 25772 12976 25828
rect 13032 25772 13100 25828
rect 13156 25772 13224 25828
rect 13280 25772 13348 25828
rect 13404 25772 13472 25828
rect 13528 25772 13596 25828
rect 13652 25772 13720 25828
rect 13776 25772 13844 25828
rect 13900 25772 13910 25828
rect 12842 25704 13910 25772
rect 12842 25648 12852 25704
rect 12908 25648 12976 25704
rect 13032 25648 13100 25704
rect 13156 25648 13224 25704
rect 13280 25648 13348 25704
rect 13404 25648 13472 25704
rect 13528 25648 13596 25704
rect 13652 25648 13720 25704
rect 13776 25648 13844 25704
rect 13900 25648 13910 25704
rect 12842 25638 13910 25648
rect 1068 25350 2136 25360
rect 1068 25294 1078 25350
rect 1134 25294 1202 25350
rect 1258 25294 1326 25350
rect 1382 25294 1450 25350
rect 1506 25294 1574 25350
rect 1630 25294 1698 25350
rect 1754 25294 1822 25350
rect 1878 25294 1946 25350
rect 2002 25294 2070 25350
rect 2126 25294 2136 25350
rect 1068 25226 2136 25294
rect 1068 25170 1078 25226
rect 1134 25170 1202 25226
rect 1258 25170 1326 25226
rect 1382 25170 1450 25226
rect 1506 25170 1574 25226
rect 1630 25170 1698 25226
rect 1754 25170 1822 25226
rect 1878 25170 1946 25226
rect 2002 25170 2070 25226
rect 2126 25170 2136 25226
rect 1068 25102 2136 25170
rect 1068 25046 1078 25102
rect 1134 25046 1202 25102
rect 1258 25046 1326 25102
rect 1382 25046 1450 25102
rect 1506 25046 1574 25102
rect 1630 25046 1698 25102
rect 1754 25046 1822 25102
rect 1878 25046 1946 25102
rect 2002 25046 2070 25102
rect 2126 25046 2136 25102
rect 1068 24978 2136 25046
rect 1068 24922 1078 24978
rect 1134 24922 1202 24978
rect 1258 24922 1326 24978
rect 1382 24922 1450 24978
rect 1506 24922 1574 24978
rect 1630 24922 1698 24978
rect 1754 24922 1822 24978
rect 1878 24922 1946 24978
rect 2002 24922 2070 24978
rect 2126 24922 2136 24978
rect 1068 24854 2136 24922
rect 1068 24798 1078 24854
rect 1134 24798 1202 24854
rect 1258 24798 1326 24854
rect 1382 24798 1450 24854
rect 1506 24798 1574 24854
rect 1630 24798 1698 24854
rect 1754 24798 1822 24854
rect 1878 24798 1946 24854
rect 2002 24798 2070 24854
rect 2126 24798 2136 24854
rect 1068 24730 2136 24798
rect 1068 24674 1078 24730
rect 1134 24674 1202 24730
rect 1258 24674 1326 24730
rect 1382 24674 1450 24730
rect 1506 24674 1574 24730
rect 1630 24674 1698 24730
rect 1754 24674 1822 24730
rect 1878 24674 1946 24730
rect 2002 24674 2070 24730
rect 2126 24674 2136 24730
rect 1068 24606 2136 24674
rect 1068 24550 1078 24606
rect 1134 24550 1202 24606
rect 1258 24550 1326 24606
rect 1382 24550 1450 24606
rect 1506 24550 1574 24606
rect 1630 24550 1698 24606
rect 1754 24550 1822 24606
rect 1878 24550 1946 24606
rect 2002 24550 2070 24606
rect 2126 24550 2136 24606
rect 1068 24482 2136 24550
rect 1068 24426 1078 24482
rect 1134 24426 1202 24482
rect 1258 24426 1326 24482
rect 1382 24426 1450 24482
rect 1506 24426 1574 24482
rect 1630 24426 1698 24482
rect 1754 24426 1822 24482
rect 1878 24426 1946 24482
rect 2002 24426 2070 24482
rect 2126 24426 2136 24482
rect 1068 24358 2136 24426
rect 1068 24302 1078 24358
rect 1134 24302 1202 24358
rect 1258 24302 1326 24358
rect 1382 24302 1450 24358
rect 1506 24302 1574 24358
rect 1630 24302 1698 24358
rect 1754 24302 1822 24358
rect 1878 24302 1946 24358
rect 2002 24302 2070 24358
rect 2126 24302 2136 24358
rect 1068 24234 2136 24302
rect 1068 24178 1078 24234
rect 1134 24178 1202 24234
rect 1258 24178 1326 24234
rect 1382 24178 1450 24234
rect 1506 24178 1574 24234
rect 1630 24178 1698 24234
rect 1754 24178 1822 24234
rect 1878 24178 1946 24234
rect 2002 24178 2070 24234
rect 2126 24178 2136 24234
rect 1068 24110 2136 24178
rect 1068 24054 1078 24110
rect 1134 24054 1202 24110
rect 1258 24054 1326 24110
rect 1382 24054 1450 24110
rect 1506 24054 1574 24110
rect 1630 24054 1698 24110
rect 1754 24054 1822 24110
rect 1878 24054 1946 24110
rect 2002 24054 2070 24110
rect 2126 24054 2136 24110
rect 1068 23986 2136 24054
rect 1068 23930 1078 23986
rect 1134 23930 1202 23986
rect 1258 23930 1326 23986
rect 1382 23930 1450 23986
rect 1506 23930 1574 23986
rect 1630 23930 1698 23986
rect 1754 23930 1822 23986
rect 1878 23930 1946 23986
rect 2002 23930 2070 23986
rect 2126 23930 2136 23986
rect 1068 23862 2136 23930
rect 1068 23806 1078 23862
rect 1134 23806 1202 23862
rect 1258 23806 1326 23862
rect 1382 23806 1450 23862
rect 1506 23806 1574 23862
rect 1630 23806 1698 23862
rect 1754 23806 1822 23862
rect 1878 23806 1946 23862
rect 2002 23806 2070 23862
rect 2126 23806 2136 23862
rect 1068 23738 2136 23806
rect 1068 23682 1078 23738
rect 1134 23682 1202 23738
rect 1258 23682 1326 23738
rect 1382 23682 1450 23738
rect 1506 23682 1574 23738
rect 1630 23682 1698 23738
rect 1754 23682 1822 23738
rect 1878 23682 1946 23738
rect 2002 23682 2070 23738
rect 2126 23682 2136 23738
rect 1068 23614 2136 23682
rect 1068 23558 1078 23614
rect 1134 23558 1202 23614
rect 1258 23558 1326 23614
rect 1382 23558 1450 23614
rect 1506 23558 1574 23614
rect 1630 23558 1698 23614
rect 1754 23558 1822 23614
rect 1878 23558 1946 23614
rect 2002 23558 2070 23614
rect 2126 23558 2136 23614
rect 1068 23490 2136 23558
rect 1068 23434 1078 23490
rect 1134 23434 1202 23490
rect 1258 23434 1326 23490
rect 1382 23434 1450 23490
rect 1506 23434 1574 23490
rect 1630 23434 1698 23490
rect 1754 23434 1822 23490
rect 1878 23434 1946 23490
rect 2002 23434 2070 23490
rect 2126 23434 2136 23490
rect 1068 23366 2136 23434
rect 1068 23310 1078 23366
rect 1134 23310 1202 23366
rect 1258 23310 1326 23366
rect 1382 23310 1450 23366
rect 1506 23310 1574 23366
rect 1630 23310 1698 23366
rect 1754 23310 1822 23366
rect 1878 23310 1946 23366
rect 2002 23310 2070 23366
rect 2126 23310 2136 23366
rect 1068 23242 2136 23310
rect 1068 23186 1078 23242
rect 1134 23186 1202 23242
rect 1258 23186 1326 23242
rect 1382 23186 1450 23242
rect 1506 23186 1574 23242
rect 1630 23186 1698 23242
rect 1754 23186 1822 23242
rect 1878 23186 1946 23242
rect 2002 23186 2070 23242
rect 2126 23186 2136 23242
rect 1068 23118 2136 23186
rect 1068 23062 1078 23118
rect 1134 23062 1202 23118
rect 1258 23062 1326 23118
rect 1382 23062 1450 23118
rect 1506 23062 1574 23118
rect 1630 23062 1698 23118
rect 1754 23062 1822 23118
rect 1878 23062 1946 23118
rect 2002 23062 2070 23118
rect 2126 23062 2136 23118
rect 1068 22994 2136 23062
rect 1068 22938 1078 22994
rect 1134 22938 1202 22994
rect 1258 22938 1326 22994
rect 1382 22938 1450 22994
rect 1506 22938 1574 22994
rect 1630 22938 1698 22994
rect 1754 22938 1822 22994
rect 1878 22938 1946 22994
rect 2002 22938 2070 22994
rect 2126 22938 2136 22994
rect 1068 22870 2136 22938
rect 1068 22814 1078 22870
rect 1134 22814 1202 22870
rect 1258 22814 1326 22870
rect 1382 22814 1450 22870
rect 1506 22814 1574 22870
rect 1630 22814 1698 22870
rect 1754 22814 1822 22870
rect 1878 22814 1946 22870
rect 2002 22814 2070 22870
rect 2126 22814 2136 22870
rect 1068 22746 2136 22814
rect 1068 22690 1078 22746
rect 1134 22690 1202 22746
rect 1258 22690 1326 22746
rect 1382 22690 1450 22746
rect 1506 22690 1574 22746
rect 1630 22690 1698 22746
rect 1754 22690 1822 22746
rect 1878 22690 1946 22746
rect 2002 22690 2070 22746
rect 2126 22690 2136 22746
rect 1068 22622 2136 22690
rect 1068 22566 1078 22622
rect 1134 22566 1202 22622
rect 1258 22566 1326 22622
rect 1382 22566 1450 22622
rect 1506 22566 1574 22622
rect 1630 22566 1698 22622
rect 1754 22566 1822 22622
rect 1878 22566 1946 22622
rect 2002 22566 2070 22622
rect 2126 22566 2136 22622
rect 1068 22498 2136 22566
rect 1068 22442 1078 22498
rect 1134 22442 1202 22498
rect 1258 22442 1326 22498
rect 1382 22442 1450 22498
rect 1506 22442 1574 22498
rect 1630 22442 1698 22498
rect 1754 22442 1822 22498
rect 1878 22442 1946 22498
rect 2002 22442 2070 22498
rect 2126 22442 2136 22498
rect 1068 22432 2136 22442
rect 4425 25350 6237 25360
rect 4425 25294 4435 25350
rect 4491 25294 4559 25350
rect 4615 25294 4683 25350
rect 4739 25294 4807 25350
rect 4863 25294 4931 25350
rect 4987 25294 5055 25350
rect 5111 25294 5179 25350
rect 5235 25294 5303 25350
rect 5359 25294 5427 25350
rect 5483 25294 5551 25350
rect 5607 25294 5675 25350
rect 5731 25294 5799 25350
rect 5855 25294 5923 25350
rect 5979 25294 6047 25350
rect 6103 25294 6171 25350
rect 6227 25294 6237 25350
rect 4425 25226 6237 25294
rect 4425 25170 4435 25226
rect 4491 25170 4559 25226
rect 4615 25170 4683 25226
rect 4739 25170 4807 25226
rect 4863 25170 4931 25226
rect 4987 25170 5055 25226
rect 5111 25170 5179 25226
rect 5235 25170 5303 25226
rect 5359 25170 5427 25226
rect 5483 25170 5551 25226
rect 5607 25170 5675 25226
rect 5731 25170 5799 25226
rect 5855 25170 5923 25226
rect 5979 25170 6047 25226
rect 6103 25170 6171 25226
rect 6227 25170 6237 25226
rect 4425 25102 6237 25170
rect 4425 25046 4435 25102
rect 4491 25046 4559 25102
rect 4615 25046 4683 25102
rect 4739 25046 4807 25102
rect 4863 25046 4931 25102
rect 4987 25046 5055 25102
rect 5111 25046 5179 25102
rect 5235 25046 5303 25102
rect 5359 25046 5427 25102
rect 5483 25046 5551 25102
rect 5607 25046 5675 25102
rect 5731 25046 5799 25102
rect 5855 25046 5923 25102
rect 5979 25046 6047 25102
rect 6103 25046 6171 25102
rect 6227 25046 6237 25102
rect 4425 24978 6237 25046
rect 4425 24922 4435 24978
rect 4491 24922 4559 24978
rect 4615 24922 4683 24978
rect 4739 24922 4807 24978
rect 4863 24922 4931 24978
rect 4987 24922 5055 24978
rect 5111 24922 5179 24978
rect 5235 24922 5303 24978
rect 5359 24922 5427 24978
rect 5483 24922 5551 24978
rect 5607 24922 5675 24978
rect 5731 24922 5799 24978
rect 5855 24922 5923 24978
rect 5979 24922 6047 24978
rect 6103 24922 6171 24978
rect 6227 24922 6237 24978
rect 4425 24854 6237 24922
rect 4425 24798 4435 24854
rect 4491 24798 4559 24854
rect 4615 24798 4683 24854
rect 4739 24798 4807 24854
rect 4863 24798 4931 24854
rect 4987 24798 5055 24854
rect 5111 24798 5179 24854
rect 5235 24798 5303 24854
rect 5359 24798 5427 24854
rect 5483 24798 5551 24854
rect 5607 24798 5675 24854
rect 5731 24798 5799 24854
rect 5855 24798 5923 24854
rect 5979 24798 6047 24854
rect 6103 24798 6171 24854
rect 6227 24798 6237 24854
rect 4425 24730 6237 24798
rect 4425 24674 4435 24730
rect 4491 24674 4559 24730
rect 4615 24674 4683 24730
rect 4739 24674 4807 24730
rect 4863 24674 4931 24730
rect 4987 24674 5055 24730
rect 5111 24674 5179 24730
rect 5235 24674 5303 24730
rect 5359 24674 5427 24730
rect 5483 24674 5551 24730
rect 5607 24674 5675 24730
rect 5731 24674 5799 24730
rect 5855 24674 5923 24730
rect 5979 24674 6047 24730
rect 6103 24674 6171 24730
rect 6227 24674 6237 24730
rect 4425 24606 6237 24674
rect 4425 24550 4435 24606
rect 4491 24550 4559 24606
rect 4615 24550 4683 24606
rect 4739 24550 4807 24606
rect 4863 24550 4931 24606
rect 4987 24550 5055 24606
rect 5111 24550 5179 24606
rect 5235 24550 5303 24606
rect 5359 24550 5427 24606
rect 5483 24550 5551 24606
rect 5607 24550 5675 24606
rect 5731 24550 5799 24606
rect 5855 24550 5923 24606
rect 5979 24550 6047 24606
rect 6103 24550 6171 24606
rect 6227 24550 6237 24606
rect 4425 24482 6237 24550
rect 4425 24426 4435 24482
rect 4491 24426 4559 24482
rect 4615 24426 4683 24482
rect 4739 24426 4807 24482
rect 4863 24426 4931 24482
rect 4987 24426 5055 24482
rect 5111 24426 5179 24482
rect 5235 24426 5303 24482
rect 5359 24426 5427 24482
rect 5483 24426 5551 24482
rect 5607 24426 5675 24482
rect 5731 24426 5799 24482
rect 5855 24426 5923 24482
rect 5979 24426 6047 24482
rect 6103 24426 6171 24482
rect 6227 24426 6237 24482
rect 4425 24358 6237 24426
rect 4425 24302 4435 24358
rect 4491 24302 4559 24358
rect 4615 24302 4683 24358
rect 4739 24302 4807 24358
rect 4863 24302 4931 24358
rect 4987 24302 5055 24358
rect 5111 24302 5179 24358
rect 5235 24302 5303 24358
rect 5359 24302 5427 24358
rect 5483 24302 5551 24358
rect 5607 24302 5675 24358
rect 5731 24302 5799 24358
rect 5855 24302 5923 24358
rect 5979 24302 6047 24358
rect 6103 24302 6171 24358
rect 6227 24302 6237 24358
rect 4425 24234 6237 24302
rect 4425 24178 4435 24234
rect 4491 24178 4559 24234
rect 4615 24178 4683 24234
rect 4739 24178 4807 24234
rect 4863 24178 4931 24234
rect 4987 24178 5055 24234
rect 5111 24178 5179 24234
rect 5235 24178 5303 24234
rect 5359 24178 5427 24234
rect 5483 24178 5551 24234
rect 5607 24178 5675 24234
rect 5731 24178 5799 24234
rect 5855 24178 5923 24234
rect 5979 24178 6047 24234
rect 6103 24178 6171 24234
rect 6227 24178 6237 24234
rect 4425 24110 6237 24178
rect 4425 24054 4435 24110
rect 4491 24054 4559 24110
rect 4615 24054 4683 24110
rect 4739 24054 4807 24110
rect 4863 24054 4931 24110
rect 4987 24054 5055 24110
rect 5111 24054 5179 24110
rect 5235 24054 5303 24110
rect 5359 24054 5427 24110
rect 5483 24054 5551 24110
rect 5607 24054 5675 24110
rect 5731 24054 5799 24110
rect 5855 24054 5923 24110
rect 5979 24054 6047 24110
rect 6103 24054 6171 24110
rect 6227 24054 6237 24110
rect 4425 23986 6237 24054
rect 4425 23930 4435 23986
rect 4491 23930 4559 23986
rect 4615 23930 4683 23986
rect 4739 23930 4807 23986
rect 4863 23930 4931 23986
rect 4987 23930 5055 23986
rect 5111 23930 5179 23986
rect 5235 23930 5303 23986
rect 5359 23930 5427 23986
rect 5483 23930 5551 23986
rect 5607 23930 5675 23986
rect 5731 23930 5799 23986
rect 5855 23930 5923 23986
rect 5979 23930 6047 23986
rect 6103 23930 6171 23986
rect 6227 23930 6237 23986
rect 4425 23862 6237 23930
rect 4425 23806 4435 23862
rect 4491 23806 4559 23862
rect 4615 23806 4683 23862
rect 4739 23806 4807 23862
rect 4863 23806 4931 23862
rect 4987 23806 5055 23862
rect 5111 23806 5179 23862
rect 5235 23806 5303 23862
rect 5359 23806 5427 23862
rect 5483 23806 5551 23862
rect 5607 23806 5675 23862
rect 5731 23806 5799 23862
rect 5855 23806 5923 23862
rect 5979 23806 6047 23862
rect 6103 23806 6171 23862
rect 6227 23806 6237 23862
rect 4425 23738 6237 23806
rect 4425 23682 4435 23738
rect 4491 23682 4559 23738
rect 4615 23682 4683 23738
rect 4739 23682 4807 23738
rect 4863 23682 4931 23738
rect 4987 23682 5055 23738
rect 5111 23682 5179 23738
rect 5235 23682 5303 23738
rect 5359 23682 5427 23738
rect 5483 23682 5551 23738
rect 5607 23682 5675 23738
rect 5731 23682 5799 23738
rect 5855 23682 5923 23738
rect 5979 23682 6047 23738
rect 6103 23682 6171 23738
rect 6227 23682 6237 23738
rect 4425 23614 6237 23682
rect 4425 23558 4435 23614
rect 4491 23558 4559 23614
rect 4615 23558 4683 23614
rect 4739 23558 4807 23614
rect 4863 23558 4931 23614
rect 4987 23558 5055 23614
rect 5111 23558 5179 23614
rect 5235 23558 5303 23614
rect 5359 23558 5427 23614
rect 5483 23558 5551 23614
rect 5607 23558 5675 23614
rect 5731 23558 5799 23614
rect 5855 23558 5923 23614
rect 5979 23558 6047 23614
rect 6103 23558 6171 23614
rect 6227 23558 6237 23614
rect 4425 23490 6237 23558
rect 4425 23434 4435 23490
rect 4491 23434 4559 23490
rect 4615 23434 4683 23490
rect 4739 23434 4807 23490
rect 4863 23434 4931 23490
rect 4987 23434 5055 23490
rect 5111 23434 5179 23490
rect 5235 23434 5303 23490
rect 5359 23434 5427 23490
rect 5483 23434 5551 23490
rect 5607 23434 5675 23490
rect 5731 23434 5799 23490
rect 5855 23434 5923 23490
rect 5979 23434 6047 23490
rect 6103 23434 6171 23490
rect 6227 23434 6237 23490
rect 4425 23366 6237 23434
rect 4425 23310 4435 23366
rect 4491 23310 4559 23366
rect 4615 23310 4683 23366
rect 4739 23310 4807 23366
rect 4863 23310 4931 23366
rect 4987 23310 5055 23366
rect 5111 23310 5179 23366
rect 5235 23310 5303 23366
rect 5359 23310 5427 23366
rect 5483 23310 5551 23366
rect 5607 23310 5675 23366
rect 5731 23310 5799 23366
rect 5855 23310 5923 23366
rect 5979 23310 6047 23366
rect 6103 23310 6171 23366
rect 6227 23310 6237 23366
rect 4425 23242 6237 23310
rect 4425 23186 4435 23242
rect 4491 23186 4559 23242
rect 4615 23186 4683 23242
rect 4739 23186 4807 23242
rect 4863 23186 4931 23242
rect 4987 23186 5055 23242
rect 5111 23186 5179 23242
rect 5235 23186 5303 23242
rect 5359 23186 5427 23242
rect 5483 23186 5551 23242
rect 5607 23186 5675 23242
rect 5731 23186 5799 23242
rect 5855 23186 5923 23242
rect 5979 23186 6047 23242
rect 6103 23186 6171 23242
rect 6227 23186 6237 23242
rect 4425 23118 6237 23186
rect 4425 23062 4435 23118
rect 4491 23062 4559 23118
rect 4615 23062 4683 23118
rect 4739 23062 4807 23118
rect 4863 23062 4931 23118
rect 4987 23062 5055 23118
rect 5111 23062 5179 23118
rect 5235 23062 5303 23118
rect 5359 23062 5427 23118
rect 5483 23062 5551 23118
rect 5607 23062 5675 23118
rect 5731 23062 5799 23118
rect 5855 23062 5923 23118
rect 5979 23062 6047 23118
rect 6103 23062 6171 23118
rect 6227 23062 6237 23118
rect 4425 22994 6237 23062
rect 4425 22938 4435 22994
rect 4491 22938 4559 22994
rect 4615 22938 4683 22994
rect 4739 22938 4807 22994
rect 4863 22938 4931 22994
rect 4987 22938 5055 22994
rect 5111 22938 5179 22994
rect 5235 22938 5303 22994
rect 5359 22938 5427 22994
rect 5483 22938 5551 22994
rect 5607 22938 5675 22994
rect 5731 22938 5799 22994
rect 5855 22938 5923 22994
rect 5979 22938 6047 22994
rect 6103 22938 6171 22994
rect 6227 22938 6237 22994
rect 4425 22870 6237 22938
rect 4425 22814 4435 22870
rect 4491 22814 4559 22870
rect 4615 22814 4683 22870
rect 4739 22814 4807 22870
rect 4863 22814 4931 22870
rect 4987 22814 5055 22870
rect 5111 22814 5179 22870
rect 5235 22814 5303 22870
rect 5359 22814 5427 22870
rect 5483 22814 5551 22870
rect 5607 22814 5675 22870
rect 5731 22814 5799 22870
rect 5855 22814 5923 22870
rect 5979 22814 6047 22870
rect 6103 22814 6171 22870
rect 6227 22814 6237 22870
rect 4425 22746 6237 22814
rect 4425 22690 4435 22746
rect 4491 22690 4559 22746
rect 4615 22690 4683 22746
rect 4739 22690 4807 22746
rect 4863 22690 4931 22746
rect 4987 22690 5055 22746
rect 5111 22690 5179 22746
rect 5235 22690 5303 22746
rect 5359 22690 5427 22746
rect 5483 22690 5551 22746
rect 5607 22690 5675 22746
rect 5731 22690 5799 22746
rect 5855 22690 5923 22746
rect 5979 22690 6047 22746
rect 6103 22690 6171 22746
rect 6227 22690 6237 22746
rect 4425 22622 6237 22690
rect 4425 22566 4435 22622
rect 4491 22566 4559 22622
rect 4615 22566 4683 22622
rect 4739 22566 4807 22622
rect 4863 22566 4931 22622
rect 4987 22566 5055 22622
rect 5111 22566 5179 22622
rect 5235 22566 5303 22622
rect 5359 22566 5427 22622
rect 5483 22566 5551 22622
rect 5607 22566 5675 22622
rect 5731 22566 5799 22622
rect 5855 22566 5923 22622
rect 5979 22566 6047 22622
rect 6103 22566 6171 22622
rect 6227 22566 6237 22622
rect 4425 22498 6237 22566
rect 4425 22442 4435 22498
rect 4491 22442 4559 22498
rect 4615 22442 4683 22498
rect 4739 22442 4807 22498
rect 4863 22442 4931 22498
rect 4987 22442 5055 22498
rect 5111 22442 5179 22498
rect 5235 22442 5303 22498
rect 5359 22442 5427 22498
rect 5483 22442 5551 22498
rect 5607 22442 5675 22498
rect 5731 22442 5799 22498
rect 5855 22442 5923 22498
rect 5979 22442 6047 22498
rect 6103 22442 6171 22498
rect 6227 22442 6237 22498
rect 4425 22432 6237 22442
rect 7552 25350 8620 25360
rect 7552 25294 7562 25350
rect 7618 25294 7686 25350
rect 7742 25294 7810 25350
rect 7866 25294 7934 25350
rect 7990 25294 8058 25350
rect 8114 25294 8182 25350
rect 8238 25294 8306 25350
rect 8362 25294 8430 25350
rect 8486 25294 8554 25350
rect 8610 25294 8620 25350
rect 7552 25226 8620 25294
rect 7552 25170 7562 25226
rect 7618 25170 7686 25226
rect 7742 25170 7810 25226
rect 7866 25170 7934 25226
rect 7990 25170 8058 25226
rect 8114 25170 8182 25226
rect 8238 25170 8306 25226
rect 8362 25170 8430 25226
rect 8486 25170 8554 25226
rect 8610 25170 8620 25226
rect 7552 25102 8620 25170
rect 7552 25046 7562 25102
rect 7618 25046 7686 25102
rect 7742 25046 7810 25102
rect 7866 25046 7934 25102
rect 7990 25046 8058 25102
rect 8114 25046 8182 25102
rect 8238 25046 8306 25102
rect 8362 25046 8430 25102
rect 8486 25046 8554 25102
rect 8610 25046 8620 25102
rect 7552 24978 8620 25046
rect 7552 24922 7562 24978
rect 7618 24922 7686 24978
rect 7742 24922 7810 24978
rect 7866 24922 7934 24978
rect 7990 24922 8058 24978
rect 8114 24922 8182 24978
rect 8238 24922 8306 24978
rect 8362 24922 8430 24978
rect 8486 24922 8554 24978
rect 8610 24922 8620 24978
rect 7552 24854 8620 24922
rect 7552 24798 7562 24854
rect 7618 24798 7686 24854
rect 7742 24798 7810 24854
rect 7866 24798 7934 24854
rect 7990 24798 8058 24854
rect 8114 24798 8182 24854
rect 8238 24798 8306 24854
rect 8362 24798 8430 24854
rect 8486 24798 8554 24854
rect 8610 24798 8620 24854
rect 7552 24730 8620 24798
rect 7552 24674 7562 24730
rect 7618 24674 7686 24730
rect 7742 24674 7810 24730
rect 7866 24674 7934 24730
rect 7990 24674 8058 24730
rect 8114 24674 8182 24730
rect 8238 24674 8306 24730
rect 8362 24674 8430 24730
rect 8486 24674 8554 24730
rect 8610 24674 8620 24730
rect 7552 24606 8620 24674
rect 7552 24550 7562 24606
rect 7618 24550 7686 24606
rect 7742 24550 7810 24606
rect 7866 24550 7934 24606
rect 7990 24550 8058 24606
rect 8114 24550 8182 24606
rect 8238 24550 8306 24606
rect 8362 24550 8430 24606
rect 8486 24550 8554 24606
rect 8610 24550 8620 24606
rect 7552 24482 8620 24550
rect 7552 24426 7562 24482
rect 7618 24426 7686 24482
rect 7742 24426 7810 24482
rect 7866 24426 7934 24482
rect 7990 24426 8058 24482
rect 8114 24426 8182 24482
rect 8238 24426 8306 24482
rect 8362 24426 8430 24482
rect 8486 24426 8554 24482
rect 8610 24426 8620 24482
rect 7552 24358 8620 24426
rect 7552 24302 7562 24358
rect 7618 24302 7686 24358
rect 7742 24302 7810 24358
rect 7866 24302 7934 24358
rect 7990 24302 8058 24358
rect 8114 24302 8182 24358
rect 8238 24302 8306 24358
rect 8362 24302 8430 24358
rect 8486 24302 8554 24358
rect 8610 24302 8620 24358
rect 7552 24234 8620 24302
rect 7552 24178 7562 24234
rect 7618 24178 7686 24234
rect 7742 24178 7810 24234
rect 7866 24178 7934 24234
rect 7990 24178 8058 24234
rect 8114 24178 8182 24234
rect 8238 24178 8306 24234
rect 8362 24178 8430 24234
rect 8486 24178 8554 24234
rect 8610 24178 8620 24234
rect 7552 24110 8620 24178
rect 7552 24054 7562 24110
rect 7618 24054 7686 24110
rect 7742 24054 7810 24110
rect 7866 24054 7934 24110
rect 7990 24054 8058 24110
rect 8114 24054 8182 24110
rect 8238 24054 8306 24110
rect 8362 24054 8430 24110
rect 8486 24054 8554 24110
rect 8610 24054 8620 24110
rect 7552 23986 8620 24054
rect 7552 23930 7562 23986
rect 7618 23930 7686 23986
rect 7742 23930 7810 23986
rect 7866 23930 7934 23986
rect 7990 23930 8058 23986
rect 8114 23930 8182 23986
rect 8238 23930 8306 23986
rect 8362 23930 8430 23986
rect 8486 23930 8554 23986
rect 8610 23930 8620 23986
rect 7552 23862 8620 23930
rect 7552 23806 7562 23862
rect 7618 23806 7686 23862
rect 7742 23806 7810 23862
rect 7866 23806 7934 23862
rect 7990 23806 8058 23862
rect 8114 23806 8182 23862
rect 8238 23806 8306 23862
rect 8362 23806 8430 23862
rect 8486 23806 8554 23862
rect 8610 23806 8620 23862
rect 7552 23738 8620 23806
rect 7552 23682 7562 23738
rect 7618 23682 7686 23738
rect 7742 23682 7810 23738
rect 7866 23682 7934 23738
rect 7990 23682 8058 23738
rect 8114 23682 8182 23738
rect 8238 23682 8306 23738
rect 8362 23682 8430 23738
rect 8486 23682 8554 23738
rect 8610 23682 8620 23738
rect 7552 23614 8620 23682
rect 7552 23558 7562 23614
rect 7618 23558 7686 23614
rect 7742 23558 7810 23614
rect 7866 23558 7934 23614
rect 7990 23558 8058 23614
rect 8114 23558 8182 23614
rect 8238 23558 8306 23614
rect 8362 23558 8430 23614
rect 8486 23558 8554 23614
rect 8610 23558 8620 23614
rect 7552 23490 8620 23558
rect 7552 23434 7562 23490
rect 7618 23434 7686 23490
rect 7742 23434 7810 23490
rect 7866 23434 7934 23490
rect 7990 23434 8058 23490
rect 8114 23434 8182 23490
rect 8238 23434 8306 23490
rect 8362 23434 8430 23490
rect 8486 23434 8554 23490
rect 8610 23434 8620 23490
rect 7552 23366 8620 23434
rect 7552 23310 7562 23366
rect 7618 23310 7686 23366
rect 7742 23310 7810 23366
rect 7866 23310 7934 23366
rect 7990 23310 8058 23366
rect 8114 23310 8182 23366
rect 8238 23310 8306 23366
rect 8362 23310 8430 23366
rect 8486 23310 8554 23366
rect 8610 23310 8620 23366
rect 7552 23242 8620 23310
rect 7552 23186 7562 23242
rect 7618 23186 7686 23242
rect 7742 23186 7810 23242
rect 7866 23186 7934 23242
rect 7990 23186 8058 23242
rect 8114 23186 8182 23242
rect 8238 23186 8306 23242
rect 8362 23186 8430 23242
rect 8486 23186 8554 23242
rect 8610 23186 8620 23242
rect 7552 23118 8620 23186
rect 7552 23062 7562 23118
rect 7618 23062 7686 23118
rect 7742 23062 7810 23118
rect 7866 23062 7934 23118
rect 7990 23062 8058 23118
rect 8114 23062 8182 23118
rect 8238 23062 8306 23118
rect 8362 23062 8430 23118
rect 8486 23062 8554 23118
rect 8610 23062 8620 23118
rect 7552 22994 8620 23062
rect 7552 22938 7562 22994
rect 7618 22938 7686 22994
rect 7742 22938 7810 22994
rect 7866 22938 7934 22994
rect 7990 22938 8058 22994
rect 8114 22938 8182 22994
rect 8238 22938 8306 22994
rect 8362 22938 8430 22994
rect 8486 22938 8554 22994
rect 8610 22938 8620 22994
rect 7552 22870 8620 22938
rect 7552 22814 7562 22870
rect 7618 22814 7686 22870
rect 7742 22814 7810 22870
rect 7866 22814 7934 22870
rect 7990 22814 8058 22870
rect 8114 22814 8182 22870
rect 8238 22814 8306 22870
rect 8362 22814 8430 22870
rect 8486 22814 8554 22870
rect 8610 22814 8620 22870
rect 7552 22746 8620 22814
rect 7552 22690 7562 22746
rect 7618 22690 7686 22746
rect 7742 22690 7810 22746
rect 7866 22690 7934 22746
rect 7990 22690 8058 22746
rect 8114 22690 8182 22746
rect 8238 22690 8306 22746
rect 8362 22690 8430 22746
rect 8486 22690 8554 22746
rect 8610 22690 8620 22746
rect 7552 22622 8620 22690
rect 7552 22566 7562 22622
rect 7618 22566 7686 22622
rect 7742 22566 7810 22622
rect 7866 22566 7934 22622
rect 7990 22566 8058 22622
rect 8114 22566 8182 22622
rect 8238 22566 8306 22622
rect 8362 22566 8430 22622
rect 8486 22566 8554 22622
rect 8610 22566 8620 22622
rect 7552 22498 8620 22566
rect 7552 22442 7562 22498
rect 7618 22442 7686 22498
rect 7742 22442 7810 22498
rect 7866 22442 7934 22498
rect 7990 22442 8058 22498
rect 8114 22442 8182 22498
rect 8238 22442 8306 22498
rect 8362 22442 8430 22498
rect 8486 22442 8554 22498
rect 8610 22442 8620 22498
rect 7552 22432 8620 22442
rect 10669 25350 12481 25360
rect 10669 25294 10679 25350
rect 10735 25294 10803 25350
rect 10859 25294 10927 25350
rect 10983 25294 11051 25350
rect 11107 25294 11175 25350
rect 11231 25294 11299 25350
rect 11355 25294 11423 25350
rect 11479 25294 11547 25350
rect 11603 25294 11671 25350
rect 11727 25294 11795 25350
rect 11851 25294 11919 25350
rect 11975 25294 12043 25350
rect 12099 25294 12167 25350
rect 12223 25294 12291 25350
rect 12347 25294 12415 25350
rect 12471 25294 12481 25350
rect 10669 25226 12481 25294
rect 10669 25170 10679 25226
rect 10735 25170 10803 25226
rect 10859 25170 10927 25226
rect 10983 25170 11051 25226
rect 11107 25170 11175 25226
rect 11231 25170 11299 25226
rect 11355 25170 11423 25226
rect 11479 25170 11547 25226
rect 11603 25170 11671 25226
rect 11727 25170 11795 25226
rect 11851 25170 11919 25226
rect 11975 25170 12043 25226
rect 12099 25170 12167 25226
rect 12223 25170 12291 25226
rect 12347 25170 12415 25226
rect 12471 25170 12481 25226
rect 10669 25102 12481 25170
rect 10669 25046 10679 25102
rect 10735 25046 10803 25102
rect 10859 25046 10927 25102
rect 10983 25046 11051 25102
rect 11107 25046 11175 25102
rect 11231 25046 11299 25102
rect 11355 25046 11423 25102
rect 11479 25046 11547 25102
rect 11603 25046 11671 25102
rect 11727 25046 11795 25102
rect 11851 25046 11919 25102
rect 11975 25046 12043 25102
rect 12099 25046 12167 25102
rect 12223 25046 12291 25102
rect 12347 25046 12415 25102
rect 12471 25046 12481 25102
rect 10669 24978 12481 25046
rect 10669 24922 10679 24978
rect 10735 24922 10803 24978
rect 10859 24922 10927 24978
rect 10983 24922 11051 24978
rect 11107 24922 11175 24978
rect 11231 24922 11299 24978
rect 11355 24922 11423 24978
rect 11479 24922 11547 24978
rect 11603 24922 11671 24978
rect 11727 24922 11795 24978
rect 11851 24922 11919 24978
rect 11975 24922 12043 24978
rect 12099 24922 12167 24978
rect 12223 24922 12291 24978
rect 12347 24922 12415 24978
rect 12471 24922 12481 24978
rect 10669 24854 12481 24922
rect 10669 24798 10679 24854
rect 10735 24798 10803 24854
rect 10859 24798 10927 24854
rect 10983 24798 11051 24854
rect 11107 24798 11175 24854
rect 11231 24798 11299 24854
rect 11355 24798 11423 24854
rect 11479 24798 11547 24854
rect 11603 24798 11671 24854
rect 11727 24798 11795 24854
rect 11851 24798 11919 24854
rect 11975 24798 12043 24854
rect 12099 24798 12167 24854
rect 12223 24798 12291 24854
rect 12347 24798 12415 24854
rect 12471 24798 12481 24854
rect 10669 24730 12481 24798
rect 10669 24674 10679 24730
rect 10735 24674 10803 24730
rect 10859 24674 10927 24730
rect 10983 24674 11051 24730
rect 11107 24674 11175 24730
rect 11231 24674 11299 24730
rect 11355 24674 11423 24730
rect 11479 24674 11547 24730
rect 11603 24674 11671 24730
rect 11727 24674 11795 24730
rect 11851 24674 11919 24730
rect 11975 24674 12043 24730
rect 12099 24674 12167 24730
rect 12223 24674 12291 24730
rect 12347 24674 12415 24730
rect 12471 24674 12481 24730
rect 10669 24606 12481 24674
rect 10669 24550 10679 24606
rect 10735 24550 10803 24606
rect 10859 24550 10927 24606
rect 10983 24550 11051 24606
rect 11107 24550 11175 24606
rect 11231 24550 11299 24606
rect 11355 24550 11423 24606
rect 11479 24550 11547 24606
rect 11603 24550 11671 24606
rect 11727 24550 11795 24606
rect 11851 24550 11919 24606
rect 11975 24550 12043 24606
rect 12099 24550 12167 24606
rect 12223 24550 12291 24606
rect 12347 24550 12415 24606
rect 12471 24550 12481 24606
rect 10669 24482 12481 24550
rect 10669 24426 10679 24482
rect 10735 24426 10803 24482
rect 10859 24426 10927 24482
rect 10983 24426 11051 24482
rect 11107 24426 11175 24482
rect 11231 24426 11299 24482
rect 11355 24426 11423 24482
rect 11479 24426 11547 24482
rect 11603 24426 11671 24482
rect 11727 24426 11795 24482
rect 11851 24426 11919 24482
rect 11975 24426 12043 24482
rect 12099 24426 12167 24482
rect 12223 24426 12291 24482
rect 12347 24426 12415 24482
rect 12471 24426 12481 24482
rect 10669 24358 12481 24426
rect 10669 24302 10679 24358
rect 10735 24302 10803 24358
rect 10859 24302 10927 24358
rect 10983 24302 11051 24358
rect 11107 24302 11175 24358
rect 11231 24302 11299 24358
rect 11355 24302 11423 24358
rect 11479 24302 11547 24358
rect 11603 24302 11671 24358
rect 11727 24302 11795 24358
rect 11851 24302 11919 24358
rect 11975 24302 12043 24358
rect 12099 24302 12167 24358
rect 12223 24302 12291 24358
rect 12347 24302 12415 24358
rect 12471 24302 12481 24358
rect 10669 24234 12481 24302
rect 10669 24178 10679 24234
rect 10735 24178 10803 24234
rect 10859 24178 10927 24234
rect 10983 24178 11051 24234
rect 11107 24178 11175 24234
rect 11231 24178 11299 24234
rect 11355 24178 11423 24234
rect 11479 24178 11547 24234
rect 11603 24178 11671 24234
rect 11727 24178 11795 24234
rect 11851 24178 11919 24234
rect 11975 24178 12043 24234
rect 12099 24178 12167 24234
rect 12223 24178 12291 24234
rect 12347 24178 12415 24234
rect 12471 24178 12481 24234
rect 10669 24110 12481 24178
rect 10669 24054 10679 24110
rect 10735 24054 10803 24110
rect 10859 24054 10927 24110
rect 10983 24054 11051 24110
rect 11107 24054 11175 24110
rect 11231 24054 11299 24110
rect 11355 24054 11423 24110
rect 11479 24054 11547 24110
rect 11603 24054 11671 24110
rect 11727 24054 11795 24110
rect 11851 24054 11919 24110
rect 11975 24054 12043 24110
rect 12099 24054 12167 24110
rect 12223 24054 12291 24110
rect 12347 24054 12415 24110
rect 12471 24054 12481 24110
rect 10669 23986 12481 24054
rect 10669 23930 10679 23986
rect 10735 23930 10803 23986
rect 10859 23930 10927 23986
rect 10983 23930 11051 23986
rect 11107 23930 11175 23986
rect 11231 23930 11299 23986
rect 11355 23930 11423 23986
rect 11479 23930 11547 23986
rect 11603 23930 11671 23986
rect 11727 23930 11795 23986
rect 11851 23930 11919 23986
rect 11975 23930 12043 23986
rect 12099 23930 12167 23986
rect 12223 23930 12291 23986
rect 12347 23930 12415 23986
rect 12471 23930 12481 23986
rect 10669 23862 12481 23930
rect 10669 23806 10679 23862
rect 10735 23806 10803 23862
rect 10859 23806 10927 23862
rect 10983 23806 11051 23862
rect 11107 23806 11175 23862
rect 11231 23806 11299 23862
rect 11355 23806 11423 23862
rect 11479 23806 11547 23862
rect 11603 23806 11671 23862
rect 11727 23806 11795 23862
rect 11851 23806 11919 23862
rect 11975 23806 12043 23862
rect 12099 23806 12167 23862
rect 12223 23806 12291 23862
rect 12347 23806 12415 23862
rect 12471 23806 12481 23862
rect 10669 23738 12481 23806
rect 10669 23682 10679 23738
rect 10735 23682 10803 23738
rect 10859 23682 10927 23738
rect 10983 23682 11051 23738
rect 11107 23682 11175 23738
rect 11231 23682 11299 23738
rect 11355 23682 11423 23738
rect 11479 23682 11547 23738
rect 11603 23682 11671 23738
rect 11727 23682 11795 23738
rect 11851 23682 11919 23738
rect 11975 23682 12043 23738
rect 12099 23682 12167 23738
rect 12223 23682 12291 23738
rect 12347 23682 12415 23738
rect 12471 23682 12481 23738
rect 10669 23614 12481 23682
rect 10669 23558 10679 23614
rect 10735 23558 10803 23614
rect 10859 23558 10927 23614
rect 10983 23558 11051 23614
rect 11107 23558 11175 23614
rect 11231 23558 11299 23614
rect 11355 23558 11423 23614
rect 11479 23558 11547 23614
rect 11603 23558 11671 23614
rect 11727 23558 11795 23614
rect 11851 23558 11919 23614
rect 11975 23558 12043 23614
rect 12099 23558 12167 23614
rect 12223 23558 12291 23614
rect 12347 23558 12415 23614
rect 12471 23558 12481 23614
rect 10669 23490 12481 23558
rect 10669 23434 10679 23490
rect 10735 23434 10803 23490
rect 10859 23434 10927 23490
rect 10983 23434 11051 23490
rect 11107 23434 11175 23490
rect 11231 23434 11299 23490
rect 11355 23434 11423 23490
rect 11479 23434 11547 23490
rect 11603 23434 11671 23490
rect 11727 23434 11795 23490
rect 11851 23434 11919 23490
rect 11975 23434 12043 23490
rect 12099 23434 12167 23490
rect 12223 23434 12291 23490
rect 12347 23434 12415 23490
rect 12471 23434 12481 23490
rect 10669 23366 12481 23434
rect 10669 23310 10679 23366
rect 10735 23310 10803 23366
rect 10859 23310 10927 23366
rect 10983 23310 11051 23366
rect 11107 23310 11175 23366
rect 11231 23310 11299 23366
rect 11355 23310 11423 23366
rect 11479 23310 11547 23366
rect 11603 23310 11671 23366
rect 11727 23310 11795 23366
rect 11851 23310 11919 23366
rect 11975 23310 12043 23366
rect 12099 23310 12167 23366
rect 12223 23310 12291 23366
rect 12347 23310 12415 23366
rect 12471 23310 12481 23366
rect 10669 23242 12481 23310
rect 10669 23186 10679 23242
rect 10735 23186 10803 23242
rect 10859 23186 10927 23242
rect 10983 23186 11051 23242
rect 11107 23186 11175 23242
rect 11231 23186 11299 23242
rect 11355 23186 11423 23242
rect 11479 23186 11547 23242
rect 11603 23186 11671 23242
rect 11727 23186 11795 23242
rect 11851 23186 11919 23242
rect 11975 23186 12043 23242
rect 12099 23186 12167 23242
rect 12223 23186 12291 23242
rect 12347 23186 12415 23242
rect 12471 23186 12481 23242
rect 10669 23118 12481 23186
rect 10669 23062 10679 23118
rect 10735 23062 10803 23118
rect 10859 23062 10927 23118
rect 10983 23062 11051 23118
rect 11107 23062 11175 23118
rect 11231 23062 11299 23118
rect 11355 23062 11423 23118
rect 11479 23062 11547 23118
rect 11603 23062 11671 23118
rect 11727 23062 11795 23118
rect 11851 23062 11919 23118
rect 11975 23062 12043 23118
rect 12099 23062 12167 23118
rect 12223 23062 12291 23118
rect 12347 23062 12415 23118
rect 12471 23062 12481 23118
rect 10669 22994 12481 23062
rect 10669 22938 10679 22994
rect 10735 22938 10803 22994
rect 10859 22938 10927 22994
rect 10983 22938 11051 22994
rect 11107 22938 11175 22994
rect 11231 22938 11299 22994
rect 11355 22938 11423 22994
rect 11479 22938 11547 22994
rect 11603 22938 11671 22994
rect 11727 22938 11795 22994
rect 11851 22938 11919 22994
rect 11975 22938 12043 22994
rect 12099 22938 12167 22994
rect 12223 22938 12291 22994
rect 12347 22938 12415 22994
rect 12471 22938 12481 22994
rect 10669 22870 12481 22938
rect 10669 22814 10679 22870
rect 10735 22814 10803 22870
rect 10859 22814 10927 22870
rect 10983 22814 11051 22870
rect 11107 22814 11175 22870
rect 11231 22814 11299 22870
rect 11355 22814 11423 22870
rect 11479 22814 11547 22870
rect 11603 22814 11671 22870
rect 11727 22814 11795 22870
rect 11851 22814 11919 22870
rect 11975 22814 12043 22870
rect 12099 22814 12167 22870
rect 12223 22814 12291 22870
rect 12347 22814 12415 22870
rect 12471 22814 12481 22870
rect 10669 22746 12481 22814
rect 10669 22690 10679 22746
rect 10735 22690 10803 22746
rect 10859 22690 10927 22746
rect 10983 22690 11051 22746
rect 11107 22690 11175 22746
rect 11231 22690 11299 22746
rect 11355 22690 11423 22746
rect 11479 22690 11547 22746
rect 11603 22690 11671 22746
rect 11727 22690 11795 22746
rect 11851 22690 11919 22746
rect 11975 22690 12043 22746
rect 12099 22690 12167 22746
rect 12223 22690 12291 22746
rect 12347 22690 12415 22746
rect 12471 22690 12481 22746
rect 10669 22622 12481 22690
rect 10669 22566 10679 22622
rect 10735 22566 10803 22622
rect 10859 22566 10927 22622
rect 10983 22566 11051 22622
rect 11107 22566 11175 22622
rect 11231 22566 11299 22622
rect 11355 22566 11423 22622
rect 11479 22566 11547 22622
rect 11603 22566 11671 22622
rect 11727 22566 11795 22622
rect 11851 22566 11919 22622
rect 11975 22566 12043 22622
rect 12099 22566 12167 22622
rect 12223 22566 12291 22622
rect 12347 22566 12415 22622
rect 12471 22566 12481 22622
rect 10669 22498 12481 22566
rect 10669 22442 10679 22498
rect 10735 22442 10803 22498
rect 10859 22442 10927 22498
rect 10983 22442 11051 22498
rect 11107 22442 11175 22498
rect 11231 22442 11299 22498
rect 11355 22442 11423 22498
rect 11479 22442 11547 22498
rect 11603 22442 11671 22498
rect 11727 22442 11795 22498
rect 11851 22442 11919 22498
rect 11975 22442 12043 22498
rect 12099 22442 12167 22498
rect 12223 22442 12291 22498
rect 12347 22442 12415 22498
rect 12471 22442 12481 22498
rect 10669 22432 12481 22442
rect 1068 22150 2136 22160
rect 1068 22094 1078 22150
rect 1134 22094 1202 22150
rect 1258 22094 1326 22150
rect 1382 22094 1450 22150
rect 1506 22094 1574 22150
rect 1630 22094 1698 22150
rect 1754 22094 1822 22150
rect 1878 22094 1946 22150
rect 2002 22094 2070 22150
rect 2126 22094 2136 22150
rect 1068 22026 2136 22094
rect 1068 21970 1078 22026
rect 1134 21970 1202 22026
rect 1258 21970 1326 22026
rect 1382 21970 1450 22026
rect 1506 21970 1574 22026
rect 1630 21970 1698 22026
rect 1754 21970 1822 22026
rect 1878 21970 1946 22026
rect 2002 21970 2070 22026
rect 2126 21970 2136 22026
rect 1068 21902 2136 21970
rect 1068 21846 1078 21902
rect 1134 21846 1202 21902
rect 1258 21846 1326 21902
rect 1382 21846 1450 21902
rect 1506 21846 1574 21902
rect 1630 21846 1698 21902
rect 1754 21846 1822 21902
rect 1878 21846 1946 21902
rect 2002 21846 2070 21902
rect 2126 21846 2136 21902
rect 1068 21778 2136 21846
rect 1068 21722 1078 21778
rect 1134 21722 1202 21778
rect 1258 21722 1326 21778
rect 1382 21722 1450 21778
rect 1506 21722 1574 21778
rect 1630 21722 1698 21778
rect 1754 21722 1822 21778
rect 1878 21722 1946 21778
rect 2002 21722 2070 21778
rect 2126 21722 2136 21778
rect 1068 21654 2136 21722
rect 1068 21598 1078 21654
rect 1134 21598 1202 21654
rect 1258 21598 1326 21654
rect 1382 21598 1450 21654
rect 1506 21598 1574 21654
rect 1630 21598 1698 21654
rect 1754 21598 1822 21654
rect 1878 21598 1946 21654
rect 2002 21598 2070 21654
rect 2126 21598 2136 21654
rect 1068 21530 2136 21598
rect 1068 21474 1078 21530
rect 1134 21474 1202 21530
rect 1258 21474 1326 21530
rect 1382 21474 1450 21530
rect 1506 21474 1574 21530
rect 1630 21474 1698 21530
rect 1754 21474 1822 21530
rect 1878 21474 1946 21530
rect 2002 21474 2070 21530
rect 2126 21474 2136 21530
rect 1068 21406 2136 21474
rect 1068 21350 1078 21406
rect 1134 21350 1202 21406
rect 1258 21350 1326 21406
rect 1382 21350 1450 21406
rect 1506 21350 1574 21406
rect 1630 21350 1698 21406
rect 1754 21350 1822 21406
rect 1878 21350 1946 21406
rect 2002 21350 2070 21406
rect 2126 21350 2136 21406
rect 1068 21282 2136 21350
rect 1068 21226 1078 21282
rect 1134 21226 1202 21282
rect 1258 21226 1326 21282
rect 1382 21226 1450 21282
rect 1506 21226 1574 21282
rect 1630 21226 1698 21282
rect 1754 21226 1822 21282
rect 1878 21226 1946 21282
rect 2002 21226 2070 21282
rect 2126 21226 2136 21282
rect 1068 21158 2136 21226
rect 1068 21102 1078 21158
rect 1134 21102 1202 21158
rect 1258 21102 1326 21158
rect 1382 21102 1450 21158
rect 1506 21102 1574 21158
rect 1630 21102 1698 21158
rect 1754 21102 1822 21158
rect 1878 21102 1946 21158
rect 2002 21102 2070 21158
rect 2126 21102 2136 21158
rect 1068 21034 2136 21102
rect 1068 20978 1078 21034
rect 1134 20978 1202 21034
rect 1258 20978 1326 21034
rect 1382 20978 1450 21034
rect 1506 20978 1574 21034
rect 1630 20978 1698 21034
rect 1754 20978 1822 21034
rect 1878 20978 1946 21034
rect 2002 20978 2070 21034
rect 2126 20978 2136 21034
rect 1068 20910 2136 20978
rect 1068 20854 1078 20910
rect 1134 20854 1202 20910
rect 1258 20854 1326 20910
rect 1382 20854 1450 20910
rect 1506 20854 1574 20910
rect 1630 20854 1698 20910
rect 1754 20854 1822 20910
rect 1878 20854 1946 20910
rect 2002 20854 2070 20910
rect 2126 20854 2136 20910
rect 1068 20786 2136 20854
rect 1068 20730 1078 20786
rect 1134 20730 1202 20786
rect 1258 20730 1326 20786
rect 1382 20730 1450 20786
rect 1506 20730 1574 20786
rect 1630 20730 1698 20786
rect 1754 20730 1822 20786
rect 1878 20730 1946 20786
rect 2002 20730 2070 20786
rect 2126 20730 2136 20786
rect 1068 20662 2136 20730
rect 1068 20606 1078 20662
rect 1134 20606 1202 20662
rect 1258 20606 1326 20662
rect 1382 20606 1450 20662
rect 1506 20606 1574 20662
rect 1630 20606 1698 20662
rect 1754 20606 1822 20662
rect 1878 20606 1946 20662
rect 2002 20606 2070 20662
rect 2126 20606 2136 20662
rect 1068 20538 2136 20606
rect 1068 20482 1078 20538
rect 1134 20482 1202 20538
rect 1258 20482 1326 20538
rect 1382 20482 1450 20538
rect 1506 20482 1574 20538
rect 1630 20482 1698 20538
rect 1754 20482 1822 20538
rect 1878 20482 1946 20538
rect 2002 20482 2070 20538
rect 2126 20482 2136 20538
rect 1068 20414 2136 20482
rect 1068 20358 1078 20414
rect 1134 20358 1202 20414
rect 1258 20358 1326 20414
rect 1382 20358 1450 20414
rect 1506 20358 1574 20414
rect 1630 20358 1698 20414
rect 1754 20358 1822 20414
rect 1878 20358 1946 20414
rect 2002 20358 2070 20414
rect 2126 20358 2136 20414
rect 1068 20290 2136 20358
rect 1068 20234 1078 20290
rect 1134 20234 1202 20290
rect 1258 20234 1326 20290
rect 1382 20234 1450 20290
rect 1506 20234 1574 20290
rect 1630 20234 1698 20290
rect 1754 20234 1822 20290
rect 1878 20234 1946 20290
rect 2002 20234 2070 20290
rect 2126 20234 2136 20290
rect 1068 20166 2136 20234
rect 1068 20110 1078 20166
rect 1134 20110 1202 20166
rect 1258 20110 1326 20166
rect 1382 20110 1450 20166
rect 1506 20110 1574 20166
rect 1630 20110 1698 20166
rect 1754 20110 1822 20166
rect 1878 20110 1946 20166
rect 2002 20110 2070 20166
rect 2126 20110 2136 20166
rect 1068 20042 2136 20110
rect 1068 19986 1078 20042
rect 1134 19986 1202 20042
rect 1258 19986 1326 20042
rect 1382 19986 1450 20042
rect 1506 19986 1574 20042
rect 1630 19986 1698 20042
rect 1754 19986 1822 20042
rect 1878 19986 1946 20042
rect 2002 19986 2070 20042
rect 2126 19986 2136 20042
rect 1068 19918 2136 19986
rect 1068 19862 1078 19918
rect 1134 19862 1202 19918
rect 1258 19862 1326 19918
rect 1382 19862 1450 19918
rect 1506 19862 1574 19918
rect 1630 19862 1698 19918
rect 1754 19862 1822 19918
rect 1878 19862 1946 19918
rect 2002 19862 2070 19918
rect 2126 19862 2136 19918
rect 1068 19794 2136 19862
rect 1068 19738 1078 19794
rect 1134 19738 1202 19794
rect 1258 19738 1326 19794
rect 1382 19738 1450 19794
rect 1506 19738 1574 19794
rect 1630 19738 1698 19794
rect 1754 19738 1822 19794
rect 1878 19738 1946 19794
rect 2002 19738 2070 19794
rect 2126 19738 2136 19794
rect 1068 19670 2136 19738
rect 1068 19614 1078 19670
rect 1134 19614 1202 19670
rect 1258 19614 1326 19670
rect 1382 19614 1450 19670
rect 1506 19614 1574 19670
rect 1630 19614 1698 19670
rect 1754 19614 1822 19670
rect 1878 19614 1946 19670
rect 2002 19614 2070 19670
rect 2126 19614 2136 19670
rect 1068 19546 2136 19614
rect 1068 19490 1078 19546
rect 1134 19490 1202 19546
rect 1258 19490 1326 19546
rect 1382 19490 1450 19546
rect 1506 19490 1574 19546
rect 1630 19490 1698 19546
rect 1754 19490 1822 19546
rect 1878 19490 1946 19546
rect 2002 19490 2070 19546
rect 2126 19490 2136 19546
rect 1068 19422 2136 19490
rect 1068 19366 1078 19422
rect 1134 19366 1202 19422
rect 1258 19366 1326 19422
rect 1382 19366 1450 19422
rect 1506 19366 1574 19422
rect 1630 19366 1698 19422
rect 1754 19366 1822 19422
rect 1878 19366 1946 19422
rect 2002 19366 2070 19422
rect 2126 19366 2136 19422
rect 1068 19298 2136 19366
rect 1068 19242 1078 19298
rect 1134 19242 1202 19298
rect 1258 19242 1326 19298
rect 1382 19242 1450 19298
rect 1506 19242 1574 19298
rect 1630 19242 1698 19298
rect 1754 19242 1822 19298
rect 1878 19242 1946 19298
rect 2002 19242 2070 19298
rect 2126 19242 2136 19298
rect 1068 19232 2136 19242
rect 4425 22150 6237 22160
rect 4425 22094 4435 22150
rect 4491 22094 4559 22150
rect 4615 22094 4683 22150
rect 4739 22094 4807 22150
rect 4863 22094 4931 22150
rect 4987 22094 5055 22150
rect 5111 22094 5179 22150
rect 5235 22094 5303 22150
rect 5359 22094 5427 22150
rect 5483 22094 5551 22150
rect 5607 22094 5675 22150
rect 5731 22094 5799 22150
rect 5855 22094 5923 22150
rect 5979 22094 6047 22150
rect 6103 22094 6171 22150
rect 6227 22094 6237 22150
rect 4425 22026 6237 22094
rect 4425 21970 4435 22026
rect 4491 21970 4559 22026
rect 4615 21970 4683 22026
rect 4739 21970 4807 22026
rect 4863 21970 4931 22026
rect 4987 21970 5055 22026
rect 5111 21970 5179 22026
rect 5235 21970 5303 22026
rect 5359 21970 5427 22026
rect 5483 21970 5551 22026
rect 5607 21970 5675 22026
rect 5731 21970 5799 22026
rect 5855 21970 5923 22026
rect 5979 21970 6047 22026
rect 6103 21970 6171 22026
rect 6227 21970 6237 22026
rect 4425 21902 6237 21970
rect 4425 21846 4435 21902
rect 4491 21846 4559 21902
rect 4615 21846 4683 21902
rect 4739 21846 4807 21902
rect 4863 21846 4931 21902
rect 4987 21846 5055 21902
rect 5111 21846 5179 21902
rect 5235 21846 5303 21902
rect 5359 21846 5427 21902
rect 5483 21846 5551 21902
rect 5607 21846 5675 21902
rect 5731 21846 5799 21902
rect 5855 21846 5923 21902
rect 5979 21846 6047 21902
rect 6103 21846 6171 21902
rect 6227 21846 6237 21902
rect 4425 21778 6237 21846
rect 4425 21722 4435 21778
rect 4491 21722 4559 21778
rect 4615 21722 4683 21778
rect 4739 21722 4807 21778
rect 4863 21722 4931 21778
rect 4987 21722 5055 21778
rect 5111 21722 5179 21778
rect 5235 21722 5303 21778
rect 5359 21722 5427 21778
rect 5483 21722 5551 21778
rect 5607 21722 5675 21778
rect 5731 21722 5799 21778
rect 5855 21722 5923 21778
rect 5979 21722 6047 21778
rect 6103 21722 6171 21778
rect 6227 21722 6237 21778
rect 4425 21654 6237 21722
rect 4425 21598 4435 21654
rect 4491 21598 4559 21654
rect 4615 21598 4683 21654
rect 4739 21598 4807 21654
rect 4863 21598 4931 21654
rect 4987 21598 5055 21654
rect 5111 21598 5179 21654
rect 5235 21598 5303 21654
rect 5359 21598 5427 21654
rect 5483 21598 5551 21654
rect 5607 21598 5675 21654
rect 5731 21598 5799 21654
rect 5855 21598 5923 21654
rect 5979 21598 6047 21654
rect 6103 21598 6171 21654
rect 6227 21598 6237 21654
rect 4425 21530 6237 21598
rect 4425 21474 4435 21530
rect 4491 21474 4559 21530
rect 4615 21474 4683 21530
rect 4739 21474 4807 21530
rect 4863 21474 4931 21530
rect 4987 21474 5055 21530
rect 5111 21474 5179 21530
rect 5235 21474 5303 21530
rect 5359 21474 5427 21530
rect 5483 21474 5551 21530
rect 5607 21474 5675 21530
rect 5731 21474 5799 21530
rect 5855 21474 5923 21530
rect 5979 21474 6047 21530
rect 6103 21474 6171 21530
rect 6227 21474 6237 21530
rect 4425 21406 6237 21474
rect 4425 21350 4435 21406
rect 4491 21350 4559 21406
rect 4615 21350 4683 21406
rect 4739 21350 4807 21406
rect 4863 21350 4931 21406
rect 4987 21350 5055 21406
rect 5111 21350 5179 21406
rect 5235 21350 5303 21406
rect 5359 21350 5427 21406
rect 5483 21350 5551 21406
rect 5607 21350 5675 21406
rect 5731 21350 5799 21406
rect 5855 21350 5923 21406
rect 5979 21350 6047 21406
rect 6103 21350 6171 21406
rect 6227 21350 6237 21406
rect 4425 21282 6237 21350
rect 4425 21226 4435 21282
rect 4491 21226 4559 21282
rect 4615 21226 4683 21282
rect 4739 21226 4807 21282
rect 4863 21226 4931 21282
rect 4987 21226 5055 21282
rect 5111 21226 5179 21282
rect 5235 21226 5303 21282
rect 5359 21226 5427 21282
rect 5483 21226 5551 21282
rect 5607 21226 5675 21282
rect 5731 21226 5799 21282
rect 5855 21226 5923 21282
rect 5979 21226 6047 21282
rect 6103 21226 6171 21282
rect 6227 21226 6237 21282
rect 4425 21158 6237 21226
rect 4425 21102 4435 21158
rect 4491 21102 4559 21158
rect 4615 21102 4683 21158
rect 4739 21102 4807 21158
rect 4863 21102 4931 21158
rect 4987 21102 5055 21158
rect 5111 21102 5179 21158
rect 5235 21102 5303 21158
rect 5359 21102 5427 21158
rect 5483 21102 5551 21158
rect 5607 21102 5675 21158
rect 5731 21102 5799 21158
rect 5855 21102 5923 21158
rect 5979 21102 6047 21158
rect 6103 21102 6171 21158
rect 6227 21102 6237 21158
rect 4425 21034 6237 21102
rect 4425 20978 4435 21034
rect 4491 20978 4559 21034
rect 4615 20978 4683 21034
rect 4739 20978 4807 21034
rect 4863 20978 4931 21034
rect 4987 20978 5055 21034
rect 5111 20978 5179 21034
rect 5235 20978 5303 21034
rect 5359 20978 5427 21034
rect 5483 20978 5551 21034
rect 5607 20978 5675 21034
rect 5731 20978 5799 21034
rect 5855 20978 5923 21034
rect 5979 20978 6047 21034
rect 6103 20978 6171 21034
rect 6227 20978 6237 21034
rect 4425 20910 6237 20978
rect 4425 20854 4435 20910
rect 4491 20854 4559 20910
rect 4615 20854 4683 20910
rect 4739 20854 4807 20910
rect 4863 20854 4931 20910
rect 4987 20854 5055 20910
rect 5111 20854 5179 20910
rect 5235 20854 5303 20910
rect 5359 20854 5427 20910
rect 5483 20854 5551 20910
rect 5607 20854 5675 20910
rect 5731 20854 5799 20910
rect 5855 20854 5923 20910
rect 5979 20854 6047 20910
rect 6103 20854 6171 20910
rect 6227 20854 6237 20910
rect 4425 20786 6237 20854
rect 4425 20730 4435 20786
rect 4491 20730 4559 20786
rect 4615 20730 4683 20786
rect 4739 20730 4807 20786
rect 4863 20730 4931 20786
rect 4987 20730 5055 20786
rect 5111 20730 5179 20786
rect 5235 20730 5303 20786
rect 5359 20730 5427 20786
rect 5483 20730 5551 20786
rect 5607 20730 5675 20786
rect 5731 20730 5799 20786
rect 5855 20730 5923 20786
rect 5979 20730 6047 20786
rect 6103 20730 6171 20786
rect 6227 20730 6237 20786
rect 4425 20662 6237 20730
rect 4425 20606 4435 20662
rect 4491 20606 4559 20662
rect 4615 20606 4683 20662
rect 4739 20606 4807 20662
rect 4863 20606 4931 20662
rect 4987 20606 5055 20662
rect 5111 20606 5179 20662
rect 5235 20606 5303 20662
rect 5359 20606 5427 20662
rect 5483 20606 5551 20662
rect 5607 20606 5675 20662
rect 5731 20606 5799 20662
rect 5855 20606 5923 20662
rect 5979 20606 6047 20662
rect 6103 20606 6171 20662
rect 6227 20606 6237 20662
rect 4425 20538 6237 20606
rect 4425 20482 4435 20538
rect 4491 20482 4559 20538
rect 4615 20482 4683 20538
rect 4739 20482 4807 20538
rect 4863 20482 4931 20538
rect 4987 20482 5055 20538
rect 5111 20482 5179 20538
rect 5235 20482 5303 20538
rect 5359 20482 5427 20538
rect 5483 20482 5551 20538
rect 5607 20482 5675 20538
rect 5731 20482 5799 20538
rect 5855 20482 5923 20538
rect 5979 20482 6047 20538
rect 6103 20482 6171 20538
rect 6227 20482 6237 20538
rect 4425 20414 6237 20482
rect 4425 20358 4435 20414
rect 4491 20358 4559 20414
rect 4615 20358 4683 20414
rect 4739 20358 4807 20414
rect 4863 20358 4931 20414
rect 4987 20358 5055 20414
rect 5111 20358 5179 20414
rect 5235 20358 5303 20414
rect 5359 20358 5427 20414
rect 5483 20358 5551 20414
rect 5607 20358 5675 20414
rect 5731 20358 5799 20414
rect 5855 20358 5923 20414
rect 5979 20358 6047 20414
rect 6103 20358 6171 20414
rect 6227 20358 6237 20414
rect 4425 20290 6237 20358
rect 4425 20234 4435 20290
rect 4491 20234 4559 20290
rect 4615 20234 4683 20290
rect 4739 20234 4807 20290
rect 4863 20234 4931 20290
rect 4987 20234 5055 20290
rect 5111 20234 5179 20290
rect 5235 20234 5303 20290
rect 5359 20234 5427 20290
rect 5483 20234 5551 20290
rect 5607 20234 5675 20290
rect 5731 20234 5799 20290
rect 5855 20234 5923 20290
rect 5979 20234 6047 20290
rect 6103 20234 6171 20290
rect 6227 20234 6237 20290
rect 4425 20166 6237 20234
rect 4425 20110 4435 20166
rect 4491 20110 4559 20166
rect 4615 20110 4683 20166
rect 4739 20110 4807 20166
rect 4863 20110 4931 20166
rect 4987 20110 5055 20166
rect 5111 20110 5179 20166
rect 5235 20110 5303 20166
rect 5359 20110 5427 20166
rect 5483 20110 5551 20166
rect 5607 20110 5675 20166
rect 5731 20110 5799 20166
rect 5855 20110 5923 20166
rect 5979 20110 6047 20166
rect 6103 20110 6171 20166
rect 6227 20110 6237 20166
rect 4425 20042 6237 20110
rect 4425 19986 4435 20042
rect 4491 19986 4559 20042
rect 4615 19986 4683 20042
rect 4739 19986 4807 20042
rect 4863 19986 4931 20042
rect 4987 19986 5055 20042
rect 5111 19986 5179 20042
rect 5235 19986 5303 20042
rect 5359 19986 5427 20042
rect 5483 19986 5551 20042
rect 5607 19986 5675 20042
rect 5731 19986 5799 20042
rect 5855 19986 5923 20042
rect 5979 19986 6047 20042
rect 6103 19986 6171 20042
rect 6227 19986 6237 20042
rect 4425 19918 6237 19986
rect 4425 19862 4435 19918
rect 4491 19862 4559 19918
rect 4615 19862 4683 19918
rect 4739 19862 4807 19918
rect 4863 19862 4931 19918
rect 4987 19862 5055 19918
rect 5111 19862 5179 19918
rect 5235 19862 5303 19918
rect 5359 19862 5427 19918
rect 5483 19862 5551 19918
rect 5607 19862 5675 19918
rect 5731 19862 5799 19918
rect 5855 19862 5923 19918
rect 5979 19862 6047 19918
rect 6103 19862 6171 19918
rect 6227 19862 6237 19918
rect 4425 19794 6237 19862
rect 4425 19738 4435 19794
rect 4491 19738 4559 19794
rect 4615 19738 4683 19794
rect 4739 19738 4807 19794
rect 4863 19738 4931 19794
rect 4987 19738 5055 19794
rect 5111 19738 5179 19794
rect 5235 19738 5303 19794
rect 5359 19738 5427 19794
rect 5483 19738 5551 19794
rect 5607 19738 5675 19794
rect 5731 19738 5799 19794
rect 5855 19738 5923 19794
rect 5979 19738 6047 19794
rect 6103 19738 6171 19794
rect 6227 19738 6237 19794
rect 4425 19670 6237 19738
rect 4425 19614 4435 19670
rect 4491 19614 4559 19670
rect 4615 19614 4683 19670
rect 4739 19614 4807 19670
rect 4863 19614 4931 19670
rect 4987 19614 5055 19670
rect 5111 19614 5179 19670
rect 5235 19614 5303 19670
rect 5359 19614 5427 19670
rect 5483 19614 5551 19670
rect 5607 19614 5675 19670
rect 5731 19614 5799 19670
rect 5855 19614 5923 19670
rect 5979 19614 6047 19670
rect 6103 19614 6171 19670
rect 6227 19614 6237 19670
rect 4425 19546 6237 19614
rect 4425 19490 4435 19546
rect 4491 19490 4559 19546
rect 4615 19490 4683 19546
rect 4739 19490 4807 19546
rect 4863 19490 4931 19546
rect 4987 19490 5055 19546
rect 5111 19490 5179 19546
rect 5235 19490 5303 19546
rect 5359 19490 5427 19546
rect 5483 19490 5551 19546
rect 5607 19490 5675 19546
rect 5731 19490 5799 19546
rect 5855 19490 5923 19546
rect 5979 19490 6047 19546
rect 6103 19490 6171 19546
rect 6227 19490 6237 19546
rect 4425 19422 6237 19490
rect 4425 19366 4435 19422
rect 4491 19366 4559 19422
rect 4615 19366 4683 19422
rect 4739 19366 4807 19422
rect 4863 19366 4931 19422
rect 4987 19366 5055 19422
rect 5111 19366 5179 19422
rect 5235 19366 5303 19422
rect 5359 19366 5427 19422
rect 5483 19366 5551 19422
rect 5607 19366 5675 19422
rect 5731 19366 5799 19422
rect 5855 19366 5923 19422
rect 5979 19366 6047 19422
rect 6103 19366 6171 19422
rect 6227 19366 6237 19422
rect 4425 19298 6237 19366
rect 4425 19242 4435 19298
rect 4491 19242 4559 19298
rect 4615 19242 4683 19298
rect 4739 19242 4807 19298
rect 4863 19242 4931 19298
rect 4987 19242 5055 19298
rect 5111 19242 5179 19298
rect 5235 19242 5303 19298
rect 5359 19242 5427 19298
rect 5483 19242 5551 19298
rect 5607 19242 5675 19298
rect 5731 19242 5799 19298
rect 5855 19242 5923 19298
rect 5979 19242 6047 19298
rect 6103 19242 6171 19298
rect 6227 19242 6237 19298
rect 4425 19232 6237 19242
rect 7552 22150 8620 22160
rect 7552 22094 7562 22150
rect 7618 22094 7686 22150
rect 7742 22094 7810 22150
rect 7866 22094 7934 22150
rect 7990 22094 8058 22150
rect 8114 22094 8182 22150
rect 8238 22094 8306 22150
rect 8362 22094 8430 22150
rect 8486 22094 8554 22150
rect 8610 22094 8620 22150
rect 7552 22026 8620 22094
rect 7552 21970 7562 22026
rect 7618 21970 7686 22026
rect 7742 21970 7810 22026
rect 7866 21970 7934 22026
rect 7990 21970 8058 22026
rect 8114 21970 8182 22026
rect 8238 21970 8306 22026
rect 8362 21970 8430 22026
rect 8486 21970 8554 22026
rect 8610 21970 8620 22026
rect 7552 21902 8620 21970
rect 7552 21846 7562 21902
rect 7618 21846 7686 21902
rect 7742 21846 7810 21902
rect 7866 21846 7934 21902
rect 7990 21846 8058 21902
rect 8114 21846 8182 21902
rect 8238 21846 8306 21902
rect 8362 21846 8430 21902
rect 8486 21846 8554 21902
rect 8610 21846 8620 21902
rect 7552 21778 8620 21846
rect 7552 21722 7562 21778
rect 7618 21722 7686 21778
rect 7742 21722 7810 21778
rect 7866 21722 7934 21778
rect 7990 21722 8058 21778
rect 8114 21722 8182 21778
rect 8238 21722 8306 21778
rect 8362 21722 8430 21778
rect 8486 21722 8554 21778
rect 8610 21722 8620 21778
rect 7552 21654 8620 21722
rect 7552 21598 7562 21654
rect 7618 21598 7686 21654
rect 7742 21598 7810 21654
rect 7866 21598 7934 21654
rect 7990 21598 8058 21654
rect 8114 21598 8182 21654
rect 8238 21598 8306 21654
rect 8362 21598 8430 21654
rect 8486 21598 8554 21654
rect 8610 21598 8620 21654
rect 7552 21530 8620 21598
rect 7552 21474 7562 21530
rect 7618 21474 7686 21530
rect 7742 21474 7810 21530
rect 7866 21474 7934 21530
rect 7990 21474 8058 21530
rect 8114 21474 8182 21530
rect 8238 21474 8306 21530
rect 8362 21474 8430 21530
rect 8486 21474 8554 21530
rect 8610 21474 8620 21530
rect 7552 21406 8620 21474
rect 7552 21350 7562 21406
rect 7618 21350 7686 21406
rect 7742 21350 7810 21406
rect 7866 21350 7934 21406
rect 7990 21350 8058 21406
rect 8114 21350 8182 21406
rect 8238 21350 8306 21406
rect 8362 21350 8430 21406
rect 8486 21350 8554 21406
rect 8610 21350 8620 21406
rect 7552 21282 8620 21350
rect 7552 21226 7562 21282
rect 7618 21226 7686 21282
rect 7742 21226 7810 21282
rect 7866 21226 7934 21282
rect 7990 21226 8058 21282
rect 8114 21226 8182 21282
rect 8238 21226 8306 21282
rect 8362 21226 8430 21282
rect 8486 21226 8554 21282
rect 8610 21226 8620 21282
rect 7552 21158 8620 21226
rect 7552 21102 7562 21158
rect 7618 21102 7686 21158
rect 7742 21102 7810 21158
rect 7866 21102 7934 21158
rect 7990 21102 8058 21158
rect 8114 21102 8182 21158
rect 8238 21102 8306 21158
rect 8362 21102 8430 21158
rect 8486 21102 8554 21158
rect 8610 21102 8620 21158
rect 7552 21034 8620 21102
rect 7552 20978 7562 21034
rect 7618 20978 7686 21034
rect 7742 20978 7810 21034
rect 7866 20978 7934 21034
rect 7990 20978 8058 21034
rect 8114 20978 8182 21034
rect 8238 20978 8306 21034
rect 8362 20978 8430 21034
rect 8486 20978 8554 21034
rect 8610 20978 8620 21034
rect 7552 20910 8620 20978
rect 7552 20854 7562 20910
rect 7618 20854 7686 20910
rect 7742 20854 7810 20910
rect 7866 20854 7934 20910
rect 7990 20854 8058 20910
rect 8114 20854 8182 20910
rect 8238 20854 8306 20910
rect 8362 20854 8430 20910
rect 8486 20854 8554 20910
rect 8610 20854 8620 20910
rect 7552 20786 8620 20854
rect 7552 20730 7562 20786
rect 7618 20730 7686 20786
rect 7742 20730 7810 20786
rect 7866 20730 7934 20786
rect 7990 20730 8058 20786
rect 8114 20730 8182 20786
rect 8238 20730 8306 20786
rect 8362 20730 8430 20786
rect 8486 20730 8554 20786
rect 8610 20730 8620 20786
rect 7552 20662 8620 20730
rect 7552 20606 7562 20662
rect 7618 20606 7686 20662
rect 7742 20606 7810 20662
rect 7866 20606 7934 20662
rect 7990 20606 8058 20662
rect 8114 20606 8182 20662
rect 8238 20606 8306 20662
rect 8362 20606 8430 20662
rect 8486 20606 8554 20662
rect 8610 20606 8620 20662
rect 7552 20538 8620 20606
rect 7552 20482 7562 20538
rect 7618 20482 7686 20538
rect 7742 20482 7810 20538
rect 7866 20482 7934 20538
rect 7990 20482 8058 20538
rect 8114 20482 8182 20538
rect 8238 20482 8306 20538
rect 8362 20482 8430 20538
rect 8486 20482 8554 20538
rect 8610 20482 8620 20538
rect 7552 20414 8620 20482
rect 7552 20358 7562 20414
rect 7618 20358 7686 20414
rect 7742 20358 7810 20414
rect 7866 20358 7934 20414
rect 7990 20358 8058 20414
rect 8114 20358 8182 20414
rect 8238 20358 8306 20414
rect 8362 20358 8430 20414
rect 8486 20358 8554 20414
rect 8610 20358 8620 20414
rect 7552 20290 8620 20358
rect 7552 20234 7562 20290
rect 7618 20234 7686 20290
rect 7742 20234 7810 20290
rect 7866 20234 7934 20290
rect 7990 20234 8058 20290
rect 8114 20234 8182 20290
rect 8238 20234 8306 20290
rect 8362 20234 8430 20290
rect 8486 20234 8554 20290
rect 8610 20234 8620 20290
rect 7552 20166 8620 20234
rect 7552 20110 7562 20166
rect 7618 20110 7686 20166
rect 7742 20110 7810 20166
rect 7866 20110 7934 20166
rect 7990 20110 8058 20166
rect 8114 20110 8182 20166
rect 8238 20110 8306 20166
rect 8362 20110 8430 20166
rect 8486 20110 8554 20166
rect 8610 20110 8620 20166
rect 7552 20042 8620 20110
rect 7552 19986 7562 20042
rect 7618 19986 7686 20042
rect 7742 19986 7810 20042
rect 7866 19986 7934 20042
rect 7990 19986 8058 20042
rect 8114 19986 8182 20042
rect 8238 19986 8306 20042
rect 8362 19986 8430 20042
rect 8486 19986 8554 20042
rect 8610 19986 8620 20042
rect 7552 19918 8620 19986
rect 7552 19862 7562 19918
rect 7618 19862 7686 19918
rect 7742 19862 7810 19918
rect 7866 19862 7934 19918
rect 7990 19862 8058 19918
rect 8114 19862 8182 19918
rect 8238 19862 8306 19918
rect 8362 19862 8430 19918
rect 8486 19862 8554 19918
rect 8610 19862 8620 19918
rect 7552 19794 8620 19862
rect 7552 19738 7562 19794
rect 7618 19738 7686 19794
rect 7742 19738 7810 19794
rect 7866 19738 7934 19794
rect 7990 19738 8058 19794
rect 8114 19738 8182 19794
rect 8238 19738 8306 19794
rect 8362 19738 8430 19794
rect 8486 19738 8554 19794
rect 8610 19738 8620 19794
rect 7552 19670 8620 19738
rect 7552 19614 7562 19670
rect 7618 19614 7686 19670
rect 7742 19614 7810 19670
rect 7866 19614 7934 19670
rect 7990 19614 8058 19670
rect 8114 19614 8182 19670
rect 8238 19614 8306 19670
rect 8362 19614 8430 19670
rect 8486 19614 8554 19670
rect 8610 19614 8620 19670
rect 7552 19546 8620 19614
rect 7552 19490 7562 19546
rect 7618 19490 7686 19546
rect 7742 19490 7810 19546
rect 7866 19490 7934 19546
rect 7990 19490 8058 19546
rect 8114 19490 8182 19546
rect 8238 19490 8306 19546
rect 8362 19490 8430 19546
rect 8486 19490 8554 19546
rect 8610 19490 8620 19546
rect 7552 19422 8620 19490
rect 7552 19366 7562 19422
rect 7618 19366 7686 19422
rect 7742 19366 7810 19422
rect 7866 19366 7934 19422
rect 7990 19366 8058 19422
rect 8114 19366 8182 19422
rect 8238 19366 8306 19422
rect 8362 19366 8430 19422
rect 8486 19366 8554 19422
rect 8610 19366 8620 19422
rect 7552 19298 8620 19366
rect 7552 19242 7562 19298
rect 7618 19242 7686 19298
rect 7742 19242 7810 19298
rect 7866 19242 7934 19298
rect 7990 19242 8058 19298
rect 8114 19242 8182 19298
rect 8238 19242 8306 19298
rect 8362 19242 8430 19298
rect 8486 19242 8554 19298
rect 8610 19242 8620 19298
rect 7552 19232 8620 19242
rect 10669 22150 12481 22160
rect 10669 22094 10679 22150
rect 10735 22094 10803 22150
rect 10859 22094 10927 22150
rect 10983 22094 11051 22150
rect 11107 22094 11175 22150
rect 11231 22094 11299 22150
rect 11355 22094 11423 22150
rect 11479 22094 11547 22150
rect 11603 22094 11671 22150
rect 11727 22094 11795 22150
rect 11851 22094 11919 22150
rect 11975 22094 12043 22150
rect 12099 22094 12167 22150
rect 12223 22094 12291 22150
rect 12347 22094 12415 22150
rect 12471 22094 12481 22150
rect 10669 22026 12481 22094
rect 10669 21970 10679 22026
rect 10735 21970 10803 22026
rect 10859 21970 10927 22026
rect 10983 21970 11051 22026
rect 11107 21970 11175 22026
rect 11231 21970 11299 22026
rect 11355 21970 11423 22026
rect 11479 21970 11547 22026
rect 11603 21970 11671 22026
rect 11727 21970 11795 22026
rect 11851 21970 11919 22026
rect 11975 21970 12043 22026
rect 12099 21970 12167 22026
rect 12223 21970 12291 22026
rect 12347 21970 12415 22026
rect 12471 21970 12481 22026
rect 10669 21902 12481 21970
rect 10669 21846 10679 21902
rect 10735 21846 10803 21902
rect 10859 21846 10927 21902
rect 10983 21846 11051 21902
rect 11107 21846 11175 21902
rect 11231 21846 11299 21902
rect 11355 21846 11423 21902
rect 11479 21846 11547 21902
rect 11603 21846 11671 21902
rect 11727 21846 11795 21902
rect 11851 21846 11919 21902
rect 11975 21846 12043 21902
rect 12099 21846 12167 21902
rect 12223 21846 12291 21902
rect 12347 21846 12415 21902
rect 12471 21846 12481 21902
rect 10669 21778 12481 21846
rect 10669 21722 10679 21778
rect 10735 21722 10803 21778
rect 10859 21722 10927 21778
rect 10983 21722 11051 21778
rect 11107 21722 11175 21778
rect 11231 21722 11299 21778
rect 11355 21722 11423 21778
rect 11479 21722 11547 21778
rect 11603 21722 11671 21778
rect 11727 21722 11795 21778
rect 11851 21722 11919 21778
rect 11975 21722 12043 21778
rect 12099 21722 12167 21778
rect 12223 21722 12291 21778
rect 12347 21722 12415 21778
rect 12471 21722 12481 21778
rect 10669 21654 12481 21722
rect 10669 21598 10679 21654
rect 10735 21598 10803 21654
rect 10859 21598 10927 21654
rect 10983 21598 11051 21654
rect 11107 21598 11175 21654
rect 11231 21598 11299 21654
rect 11355 21598 11423 21654
rect 11479 21598 11547 21654
rect 11603 21598 11671 21654
rect 11727 21598 11795 21654
rect 11851 21598 11919 21654
rect 11975 21598 12043 21654
rect 12099 21598 12167 21654
rect 12223 21598 12291 21654
rect 12347 21598 12415 21654
rect 12471 21598 12481 21654
rect 10669 21530 12481 21598
rect 10669 21474 10679 21530
rect 10735 21474 10803 21530
rect 10859 21474 10927 21530
rect 10983 21474 11051 21530
rect 11107 21474 11175 21530
rect 11231 21474 11299 21530
rect 11355 21474 11423 21530
rect 11479 21474 11547 21530
rect 11603 21474 11671 21530
rect 11727 21474 11795 21530
rect 11851 21474 11919 21530
rect 11975 21474 12043 21530
rect 12099 21474 12167 21530
rect 12223 21474 12291 21530
rect 12347 21474 12415 21530
rect 12471 21474 12481 21530
rect 10669 21406 12481 21474
rect 10669 21350 10679 21406
rect 10735 21350 10803 21406
rect 10859 21350 10927 21406
rect 10983 21350 11051 21406
rect 11107 21350 11175 21406
rect 11231 21350 11299 21406
rect 11355 21350 11423 21406
rect 11479 21350 11547 21406
rect 11603 21350 11671 21406
rect 11727 21350 11795 21406
rect 11851 21350 11919 21406
rect 11975 21350 12043 21406
rect 12099 21350 12167 21406
rect 12223 21350 12291 21406
rect 12347 21350 12415 21406
rect 12471 21350 12481 21406
rect 10669 21282 12481 21350
rect 10669 21226 10679 21282
rect 10735 21226 10803 21282
rect 10859 21226 10927 21282
rect 10983 21226 11051 21282
rect 11107 21226 11175 21282
rect 11231 21226 11299 21282
rect 11355 21226 11423 21282
rect 11479 21226 11547 21282
rect 11603 21226 11671 21282
rect 11727 21226 11795 21282
rect 11851 21226 11919 21282
rect 11975 21226 12043 21282
rect 12099 21226 12167 21282
rect 12223 21226 12291 21282
rect 12347 21226 12415 21282
rect 12471 21226 12481 21282
rect 10669 21158 12481 21226
rect 10669 21102 10679 21158
rect 10735 21102 10803 21158
rect 10859 21102 10927 21158
rect 10983 21102 11051 21158
rect 11107 21102 11175 21158
rect 11231 21102 11299 21158
rect 11355 21102 11423 21158
rect 11479 21102 11547 21158
rect 11603 21102 11671 21158
rect 11727 21102 11795 21158
rect 11851 21102 11919 21158
rect 11975 21102 12043 21158
rect 12099 21102 12167 21158
rect 12223 21102 12291 21158
rect 12347 21102 12415 21158
rect 12471 21102 12481 21158
rect 10669 21034 12481 21102
rect 10669 20978 10679 21034
rect 10735 20978 10803 21034
rect 10859 20978 10927 21034
rect 10983 20978 11051 21034
rect 11107 20978 11175 21034
rect 11231 20978 11299 21034
rect 11355 20978 11423 21034
rect 11479 20978 11547 21034
rect 11603 20978 11671 21034
rect 11727 20978 11795 21034
rect 11851 20978 11919 21034
rect 11975 20978 12043 21034
rect 12099 20978 12167 21034
rect 12223 20978 12291 21034
rect 12347 20978 12415 21034
rect 12471 20978 12481 21034
rect 10669 20910 12481 20978
rect 10669 20854 10679 20910
rect 10735 20854 10803 20910
rect 10859 20854 10927 20910
rect 10983 20854 11051 20910
rect 11107 20854 11175 20910
rect 11231 20854 11299 20910
rect 11355 20854 11423 20910
rect 11479 20854 11547 20910
rect 11603 20854 11671 20910
rect 11727 20854 11795 20910
rect 11851 20854 11919 20910
rect 11975 20854 12043 20910
rect 12099 20854 12167 20910
rect 12223 20854 12291 20910
rect 12347 20854 12415 20910
rect 12471 20854 12481 20910
rect 10669 20786 12481 20854
rect 10669 20730 10679 20786
rect 10735 20730 10803 20786
rect 10859 20730 10927 20786
rect 10983 20730 11051 20786
rect 11107 20730 11175 20786
rect 11231 20730 11299 20786
rect 11355 20730 11423 20786
rect 11479 20730 11547 20786
rect 11603 20730 11671 20786
rect 11727 20730 11795 20786
rect 11851 20730 11919 20786
rect 11975 20730 12043 20786
rect 12099 20730 12167 20786
rect 12223 20730 12291 20786
rect 12347 20730 12415 20786
rect 12471 20730 12481 20786
rect 10669 20662 12481 20730
rect 10669 20606 10679 20662
rect 10735 20606 10803 20662
rect 10859 20606 10927 20662
rect 10983 20606 11051 20662
rect 11107 20606 11175 20662
rect 11231 20606 11299 20662
rect 11355 20606 11423 20662
rect 11479 20606 11547 20662
rect 11603 20606 11671 20662
rect 11727 20606 11795 20662
rect 11851 20606 11919 20662
rect 11975 20606 12043 20662
rect 12099 20606 12167 20662
rect 12223 20606 12291 20662
rect 12347 20606 12415 20662
rect 12471 20606 12481 20662
rect 10669 20538 12481 20606
rect 10669 20482 10679 20538
rect 10735 20482 10803 20538
rect 10859 20482 10927 20538
rect 10983 20482 11051 20538
rect 11107 20482 11175 20538
rect 11231 20482 11299 20538
rect 11355 20482 11423 20538
rect 11479 20482 11547 20538
rect 11603 20482 11671 20538
rect 11727 20482 11795 20538
rect 11851 20482 11919 20538
rect 11975 20482 12043 20538
rect 12099 20482 12167 20538
rect 12223 20482 12291 20538
rect 12347 20482 12415 20538
rect 12471 20482 12481 20538
rect 10669 20414 12481 20482
rect 10669 20358 10679 20414
rect 10735 20358 10803 20414
rect 10859 20358 10927 20414
rect 10983 20358 11051 20414
rect 11107 20358 11175 20414
rect 11231 20358 11299 20414
rect 11355 20358 11423 20414
rect 11479 20358 11547 20414
rect 11603 20358 11671 20414
rect 11727 20358 11795 20414
rect 11851 20358 11919 20414
rect 11975 20358 12043 20414
rect 12099 20358 12167 20414
rect 12223 20358 12291 20414
rect 12347 20358 12415 20414
rect 12471 20358 12481 20414
rect 10669 20290 12481 20358
rect 10669 20234 10679 20290
rect 10735 20234 10803 20290
rect 10859 20234 10927 20290
rect 10983 20234 11051 20290
rect 11107 20234 11175 20290
rect 11231 20234 11299 20290
rect 11355 20234 11423 20290
rect 11479 20234 11547 20290
rect 11603 20234 11671 20290
rect 11727 20234 11795 20290
rect 11851 20234 11919 20290
rect 11975 20234 12043 20290
rect 12099 20234 12167 20290
rect 12223 20234 12291 20290
rect 12347 20234 12415 20290
rect 12471 20234 12481 20290
rect 10669 20166 12481 20234
rect 10669 20110 10679 20166
rect 10735 20110 10803 20166
rect 10859 20110 10927 20166
rect 10983 20110 11051 20166
rect 11107 20110 11175 20166
rect 11231 20110 11299 20166
rect 11355 20110 11423 20166
rect 11479 20110 11547 20166
rect 11603 20110 11671 20166
rect 11727 20110 11795 20166
rect 11851 20110 11919 20166
rect 11975 20110 12043 20166
rect 12099 20110 12167 20166
rect 12223 20110 12291 20166
rect 12347 20110 12415 20166
rect 12471 20110 12481 20166
rect 10669 20042 12481 20110
rect 10669 19986 10679 20042
rect 10735 19986 10803 20042
rect 10859 19986 10927 20042
rect 10983 19986 11051 20042
rect 11107 19986 11175 20042
rect 11231 19986 11299 20042
rect 11355 19986 11423 20042
rect 11479 19986 11547 20042
rect 11603 19986 11671 20042
rect 11727 19986 11795 20042
rect 11851 19986 11919 20042
rect 11975 19986 12043 20042
rect 12099 19986 12167 20042
rect 12223 19986 12291 20042
rect 12347 19986 12415 20042
rect 12471 19986 12481 20042
rect 10669 19918 12481 19986
rect 10669 19862 10679 19918
rect 10735 19862 10803 19918
rect 10859 19862 10927 19918
rect 10983 19862 11051 19918
rect 11107 19862 11175 19918
rect 11231 19862 11299 19918
rect 11355 19862 11423 19918
rect 11479 19862 11547 19918
rect 11603 19862 11671 19918
rect 11727 19862 11795 19918
rect 11851 19862 11919 19918
rect 11975 19862 12043 19918
rect 12099 19862 12167 19918
rect 12223 19862 12291 19918
rect 12347 19862 12415 19918
rect 12471 19862 12481 19918
rect 10669 19794 12481 19862
rect 10669 19738 10679 19794
rect 10735 19738 10803 19794
rect 10859 19738 10927 19794
rect 10983 19738 11051 19794
rect 11107 19738 11175 19794
rect 11231 19738 11299 19794
rect 11355 19738 11423 19794
rect 11479 19738 11547 19794
rect 11603 19738 11671 19794
rect 11727 19738 11795 19794
rect 11851 19738 11919 19794
rect 11975 19738 12043 19794
rect 12099 19738 12167 19794
rect 12223 19738 12291 19794
rect 12347 19738 12415 19794
rect 12471 19738 12481 19794
rect 10669 19670 12481 19738
rect 10669 19614 10679 19670
rect 10735 19614 10803 19670
rect 10859 19614 10927 19670
rect 10983 19614 11051 19670
rect 11107 19614 11175 19670
rect 11231 19614 11299 19670
rect 11355 19614 11423 19670
rect 11479 19614 11547 19670
rect 11603 19614 11671 19670
rect 11727 19614 11795 19670
rect 11851 19614 11919 19670
rect 11975 19614 12043 19670
rect 12099 19614 12167 19670
rect 12223 19614 12291 19670
rect 12347 19614 12415 19670
rect 12471 19614 12481 19670
rect 10669 19546 12481 19614
rect 10669 19490 10679 19546
rect 10735 19490 10803 19546
rect 10859 19490 10927 19546
rect 10983 19490 11051 19546
rect 11107 19490 11175 19546
rect 11231 19490 11299 19546
rect 11355 19490 11423 19546
rect 11479 19490 11547 19546
rect 11603 19490 11671 19546
rect 11727 19490 11795 19546
rect 11851 19490 11919 19546
rect 11975 19490 12043 19546
rect 12099 19490 12167 19546
rect 12223 19490 12291 19546
rect 12347 19490 12415 19546
rect 12471 19490 12481 19546
rect 10669 19422 12481 19490
rect 10669 19366 10679 19422
rect 10735 19366 10803 19422
rect 10859 19366 10927 19422
rect 10983 19366 11051 19422
rect 11107 19366 11175 19422
rect 11231 19366 11299 19422
rect 11355 19366 11423 19422
rect 11479 19366 11547 19422
rect 11603 19366 11671 19422
rect 11727 19366 11795 19422
rect 11851 19366 11919 19422
rect 11975 19366 12043 19422
rect 12099 19366 12167 19422
rect 12223 19366 12291 19422
rect 12347 19366 12415 19422
rect 12471 19366 12481 19422
rect 10669 19298 12481 19366
rect 10669 19242 10679 19298
rect 10735 19242 10803 19298
rect 10859 19242 10927 19298
rect 10983 19242 11051 19298
rect 11107 19242 11175 19298
rect 11231 19242 11299 19298
rect 11355 19242 11423 19298
rect 11479 19242 11547 19298
rect 11603 19242 11671 19298
rect 11727 19242 11795 19298
rect 11851 19242 11919 19298
rect 11975 19242 12043 19298
rect 12099 19242 12167 19298
rect 12223 19242 12291 19298
rect 12347 19242 12415 19298
rect 12471 19242 12481 19298
rect 10669 19232 12481 19242
rect 1068 18950 2136 18960
rect 1068 18894 1078 18950
rect 1134 18894 1202 18950
rect 1258 18894 1326 18950
rect 1382 18894 1450 18950
rect 1506 18894 1574 18950
rect 1630 18894 1698 18950
rect 1754 18894 1822 18950
rect 1878 18894 1946 18950
rect 2002 18894 2070 18950
rect 2126 18894 2136 18950
rect 1068 18826 2136 18894
rect 1068 18770 1078 18826
rect 1134 18770 1202 18826
rect 1258 18770 1326 18826
rect 1382 18770 1450 18826
rect 1506 18770 1574 18826
rect 1630 18770 1698 18826
rect 1754 18770 1822 18826
rect 1878 18770 1946 18826
rect 2002 18770 2070 18826
rect 2126 18770 2136 18826
rect 1068 18702 2136 18770
rect 1068 18646 1078 18702
rect 1134 18646 1202 18702
rect 1258 18646 1326 18702
rect 1382 18646 1450 18702
rect 1506 18646 1574 18702
rect 1630 18646 1698 18702
rect 1754 18646 1822 18702
rect 1878 18646 1946 18702
rect 2002 18646 2070 18702
rect 2126 18646 2136 18702
rect 1068 18578 2136 18646
rect 1068 18522 1078 18578
rect 1134 18522 1202 18578
rect 1258 18522 1326 18578
rect 1382 18522 1450 18578
rect 1506 18522 1574 18578
rect 1630 18522 1698 18578
rect 1754 18522 1822 18578
rect 1878 18522 1946 18578
rect 2002 18522 2070 18578
rect 2126 18522 2136 18578
rect 1068 18454 2136 18522
rect 1068 18398 1078 18454
rect 1134 18398 1202 18454
rect 1258 18398 1326 18454
rect 1382 18398 1450 18454
rect 1506 18398 1574 18454
rect 1630 18398 1698 18454
rect 1754 18398 1822 18454
rect 1878 18398 1946 18454
rect 2002 18398 2070 18454
rect 2126 18398 2136 18454
rect 1068 18330 2136 18398
rect 1068 18274 1078 18330
rect 1134 18274 1202 18330
rect 1258 18274 1326 18330
rect 1382 18274 1450 18330
rect 1506 18274 1574 18330
rect 1630 18274 1698 18330
rect 1754 18274 1822 18330
rect 1878 18274 1946 18330
rect 2002 18274 2070 18330
rect 2126 18274 2136 18330
rect 1068 18206 2136 18274
rect 1068 18150 1078 18206
rect 1134 18150 1202 18206
rect 1258 18150 1326 18206
rect 1382 18150 1450 18206
rect 1506 18150 1574 18206
rect 1630 18150 1698 18206
rect 1754 18150 1822 18206
rect 1878 18150 1946 18206
rect 2002 18150 2070 18206
rect 2126 18150 2136 18206
rect 1068 18082 2136 18150
rect 1068 18026 1078 18082
rect 1134 18026 1202 18082
rect 1258 18026 1326 18082
rect 1382 18026 1450 18082
rect 1506 18026 1574 18082
rect 1630 18026 1698 18082
rect 1754 18026 1822 18082
rect 1878 18026 1946 18082
rect 2002 18026 2070 18082
rect 2126 18026 2136 18082
rect 1068 17958 2136 18026
rect 1068 17902 1078 17958
rect 1134 17902 1202 17958
rect 1258 17902 1326 17958
rect 1382 17902 1450 17958
rect 1506 17902 1574 17958
rect 1630 17902 1698 17958
rect 1754 17902 1822 17958
rect 1878 17902 1946 17958
rect 2002 17902 2070 17958
rect 2126 17902 2136 17958
rect 1068 17834 2136 17902
rect 1068 17778 1078 17834
rect 1134 17778 1202 17834
rect 1258 17778 1326 17834
rect 1382 17778 1450 17834
rect 1506 17778 1574 17834
rect 1630 17778 1698 17834
rect 1754 17778 1822 17834
rect 1878 17778 1946 17834
rect 2002 17778 2070 17834
rect 2126 17778 2136 17834
rect 1068 17710 2136 17778
rect 1068 17654 1078 17710
rect 1134 17654 1202 17710
rect 1258 17654 1326 17710
rect 1382 17654 1450 17710
rect 1506 17654 1574 17710
rect 1630 17654 1698 17710
rect 1754 17654 1822 17710
rect 1878 17654 1946 17710
rect 2002 17654 2070 17710
rect 2126 17654 2136 17710
rect 1068 17586 2136 17654
rect 1068 17530 1078 17586
rect 1134 17530 1202 17586
rect 1258 17530 1326 17586
rect 1382 17530 1450 17586
rect 1506 17530 1574 17586
rect 1630 17530 1698 17586
rect 1754 17530 1822 17586
rect 1878 17530 1946 17586
rect 2002 17530 2070 17586
rect 2126 17530 2136 17586
rect 1068 17462 2136 17530
rect 1068 17406 1078 17462
rect 1134 17406 1202 17462
rect 1258 17406 1326 17462
rect 1382 17406 1450 17462
rect 1506 17406 1574 17462
rect 1630 17406 1698 17462
rect 1754 17406 1822 17462
rect 1878 17406 1946 17462
rect 2002 17406 2070 17462
rect 2126 17406 2136 17462
rect 1068 17338 2136 17406
rect 1068 17282 1078 17338
rect 1134 17282 1202 17338
rect 1258 17282 1326 17338
rect 1382 17282 1450 17338
rect 1506 17282 1574 17338
rect 1630 17282 1698 17338
rect 1754 17282 1822 17338
rect 1878 17282 1946 17338
rect 2002 17282 2070 17338
rect 2126 17282 2136 17338
rect 1068 17214 2136 17282
rect 1068 17158 1078 17214
rect 1134 17158 1202 17214
rect 1258 17158 1326 17214
rect 1382 17158 1450 17214
rect 1506 17158 1574 17214
rect 1630 17158 1698 17214
rect 1754 17158 1822 17214
rect 1878 17158 1946 17214
rect 2002 17158 2070 17214
rect 2126 17158 2136 17214
rect 1068 17090 2136 17158
rect 1068 17034 1078 17090
rect 1134 17034 1202 17090
rect 1258 17034 1326 17090
rect 1382 17034 1450 17090
rect 1506 17034 1574 17090
rect 1630 17034 1698 17090
rect 1754 17034 1822 17090
rect 1878 17034 1946 17090
rect 2002 17034 2070 17090
rect 2126 17034 2136 17090
rect 1068 16966 2136 17034
rect 1068 16910 1078 16966
rect 1134 16910 1202 16966
rect 1258 16910 1326 16966
rect 1382 16910 1450 16966
rect 1506 16910 1574 16966
rect 1630 16910 1698 16966
rect 1754 16910 1822 16966
rect 1878 16910 1946 16966
rect 2002 16910 2070 16966
rect 2126 16910 2136 16966
rect 1068 16842 2136 16910
rect 1068 16786 1078 16842
rect 1134 16786 1202 16842
rect 1258 16786 1326 16842
rect 1382 16786 1450 16842
rect 1506 16786 1574 16842
rect 1630 16786 1698 16842
rect 1754 16786 1822 16842
rect 1878 16786 1946 16842
rect 2002 16786 2070 16842
rect 2126 16786 2136 16842
rect 1068 16718 2136 16786
rect 1068 16662 1078 16718
rect 1134 16662 1202 16718
rect 1258 16662 1326 16718
rect 1382 16662 1450 16718
rect 1506 16662 1574 16718
rect 1630 16662 1698 16718
rect 1754 16662 1822 16718
rect 1878 16662 1946 16718
rect 2002 16662 2070 16718
rect 2126 16662 2136 16718
rect 1068 16594 2136 16662
rect 1068 16538 1078 16594
rect 1134 16538 1202 16594
rect 1258 16538 1326 16594
rect 1382 16538 1450 16594
rect 1506 16538 1574 16594
rect 1630 16538 1698 16594
rect 1754 16538 1822 16594
rect 1878 16538 1946 16594
rect 2002 16538 2070 16594
rect 2126 16538 2136 16594
rect 1068 16470 2136 16538
rect 1068 16414 1078 16470
rect 1134 16414 1202 16470
rect 1258 16414 1326 16470
rect 1382 16414 1450 16470
rect 1506 16414 1574 16470
rect 1630 16414 1698 16470
rect 1754 16414 1822 16470
rect 1878 16414 1946 16470
rect 2002 16414 2070 16470
rect 2126 16414 2136 16470
rect 1068 16346 2136 16414
rect 1068 16290 1078 16346
rect 1134 16290 1202 16346
rect 1258 16290 1326 16346
rect 1382 16290 1450 16346
rect 1506 16290 1574 16346
rect 1630 16290 1698 16346
rect 1754 16290 1822 16346
rect 1878 16290 1946 16346
rect 2002 16290 2070 16346
rect 2126 16290 2136 16346
rect 1068 16222 2136 16290
rect 1068 16166 1078 16222
rect 1134 16166 1202 16222
rect 1258 16166 1326 16222
rect 1382 16166 1450 16222
rect 1506 16166 1574 16222
rect 1630 16166 1698 16222
rect 1754 16166 1822 16222
rect 1878 16166 1946 16222
rect 2002 16166 2070 16222
rect 2126 16166 2136 16222
rect 1068 16098 2136 16166
rect 1068 16042 1078 16098
rect 1134 16042 1202 16098
rect 1258 16042 1326 16098
rect 1382 16042 1450 16098
rect 1506 16042 1574 16098
rect 1630 16042 1698 16098
rect 1754 16042 1822 16098
rect 1878 16042 1946 16098
rect 2002 16042 2070 16098
rect 2126 16042 2136 16098
rect 1068 16032 2136 16042
rect 4425 18950 6237 18960
rect 4425 18894 4435 18950
rect 4491 18894 4559 18950
rect 4615 18894 4683 18950
rect 4739 18894 4807 18950
rect 4863 18894 4931 18950
rect 4987 18894 5055 18950
rect 5111 18894 5179 18950
rect 5235 18894 5303 18950
rect 5359 18894 5427 18950
rect 5483 18894 5551 18950
rect 5607 18894 5675 18950
rect 5731 18894 5799 18950
rect 5855 18894 5923 18950
rect 5979 18894 6047 18950
rect 6103 18894 6171 18950
rect 6227 18894 6237 18950
rect 4425 18826 6237 18894
rect 4425 18770 4435 18826
rect 4491 18770 4559 18826
rect 4615 18770 4683 18826
rect 4739 18770 4807 18826
rect 4863 18770 4931 18826
rect 4987 18770 5055 18826
rect 5111 18770 5179 18826
rect 5235 18770 5303 18826
rect 5359 18770 5427 18826
rect 5483 18770 5551 18826
rect 5607 18770 5675 18826
rect 5731 18770 5799 18826
rect 5855 18770 5923 18826
rect 5979 18770 6047 18826
rect 6103 18770 6171 18826
rect 6227 18770 6237 18826
rect 4425 18702 6237 18770
rect 4425 18646 4435 18702
rect 4491 18646 4559 18702
rect 4615 18646 4683 18702
rect 4739 18646 4807 18702
rect 4863 18646 4931 18702
rect 4987 18646 5055 18702
rect 5111 18646 5179 18702
rect 5235 18646 5303 18702
rect 5359 18646 5427 18702
rect 5483 18646 5551 18702
rect 5607 18646 5675 18702
rect 5731 18646 5799 18702
rect 5855 18646 5923 18702
rect 5979 18646 6047 18702
rect 6103 18646 6171 18702
rect 6227 18646 6237 18702
rect 4425 18578 6237 18646
rect 4425 18522 4435 18578
rect 4491 18522 4559 18578
rect 4615 18522 4683 18578
rect 4739 18522 4807 18578
rect 4863 18522 4931 18578
rect 4987 18522 5055 18578
rect 5111 18522 5179 18578
rect 5235 18522 5303 18578
rect 5359 18522 5427 18578
rect 5483 18522 5551 18578
rect 5607 18522 5675 18578
rect 5731 18522 5799 18578
rect 5855 18522 5923 18578
rect 5979 18522 6047 18578
rect 6103 18522 6171 18578
rect 6227 18522 6237 18578
rect 4425 18454 6237 18522
rect 4425 18398 4435 18454
rect 4491 18398 4559 18454
rect 4615 18398 4683 18454
rect 4739 18398 4807 18454
rect 4863 18398 4931 18454
rect 4987 18398 5055 18454
rect 5111 18398 5179 18454
rect 5235 18398 5303 18454
rect 5359 18398 5427 18454
rect 5483 18398 5551 18454
rect 5607 18398 5675 18454
rect 5731 18398 5799 18454
rect 5855 18398 5923 18454
rect 5979 18398 6047 18454
rect 6103 18398 6171 18454
rect 6227 18398 6237 18454
rect 4425 18330 6237 18398
rect 4425 18274 4435 18330
rect 4491 18274 4559 18330
rect 4615 18274 4683 18330
rect 4739 18274 4807 18330
rect 4863 18274 4931 18330
rect 4987 18274 5055 18330
rect 5111 18274 5179 18330
rect 5235 18274 5303 18330
rect 5359 18274 5427 18330
rect 5483 18274 5551 18330
rect 5607 18274 5675 18330
rect 5731 18274 5799 18330
rect 5855 18274 5923 18330
rect 5979 18274 6047 18330
rect 6103 18274 6171 18330
rect 6227 18274 6237 18330
rect 4425 18206 6237 18274
rect 4425 18150 4435 18206
rect 4491 18150 4559 18206
rect 4615 18150 4683 18206
rect 4739 18150 4807 18206
rect 4863 18150 4931 18206
rect 4987 18150 5055 18206
rect 5111 18150 5179 18206
rect 5235 18150 5303 18206
rect 5359 18150 5427 18206
rect 5483 18150 5551 18206
rect 5607 18150 5675 18206
rect 5731 18150 5799 18206
rect 5855 18150 5923 18206
rect 5979 18150 6047 18206
rect 6103 18150 6171 18206
rect 6227 18150 6237 18206
rect 4425 18082 6237 18150
rect 4425 18026 4435 18082
rect 4491 18026 4559 18082
rect 4615 18026 4683 18082
rect 4739 18026 4807 18082
rect 4863 18026 4931 18082
rect 4987 18026 5055 18082
rect 5111 18026 5179 18082
rect 5235 18026 5303 18082
rect 5359 18026 5427 18082
rect 5483 18026 5551 18082
rect 5607 18026 5675 18082
rect 5731 18026 5799 18082
rect 5855 18026 5923 18082
rect 5979 18026 6047 18082
rect 6103 18026 6171 18082
rect 6227 18026 6237 18082
rect 4425 17958 6237 18026
rect 4425 17902 4435 17958
rect 4491 17902 4559 17958
rect 4615 17902 4683 17958
rect 4739 17902 4807 17958
rect 4863 17902 4931 17958
rect 4987 17902 5055 17958
rect 5111 17902 5179 17958
rect 5235 17902 5303 17958
rect 5359 17902 5427 17958
rect 5483 17902 5551 17958
rect 5607 17902 5675 17958
rect 5731 17902 5799 17958
rect 5855 17902 5923 17958
rect 5979 17902 6047 17958
rect 6103 17902 6171 17958
rect 6227 17902 6237 17958
rect 4425 17834 6237 17902
rect 4425 17778 4435 17834
rect 4491 17778 4559 17834
rect 4615 17778 4683 17834
rect 4739 17778 4807 17834
rect 4863 17778 4931 17834
rect 4987 17778 5055 17834
rect 5111 17778 5179 17834
rect 5235 17778 5303 17834
rect 5359 17778 5427 17834
rect 5483 17778 5551 17834
rect 5607 17778 5675 17834
rect 5731 17778 5799 17834
rect 5855 17778 5923 17834
rect 5979 17778 6047 17834
rect 6103 17778 6171 17834
rect 6227 17778 6237 17834
rect 4425 17710 6237 17778
rect 4425 17654 4435 17710
rect 4491 17654 4559 17710
rect 4615 17654 4683 17710
rect 4739 17654 4807 17710
rect 4863 17654 4931 17710
rect 4987 17654 5055 17710
rect 5111 17654 5179 17710
rect 5235 17654 5303 17710
rect 5359 17654 5427 17710
rect 5483 17654 5551 17710
rect 5607 17654 5675 17710
rect 5731 17654 5799 17710
rect 5855 17654 5923 17710
rect 5979 17654 6047 17710
rect 6103 17654 6171 17710
rect 6227 17654 6237 17710
rect 4425 17586 6237 17654
rect 4425 17530 4435 17586
rect 4491 17530 4559 17586
rect 4615 17530 4683 17586
rect 4739 17530 4807 17586
rect 4863 17530 4931 17586
rect 4987 17530 5055 17586
rect 5111 17530 5179 17586
rect 5235 17530 5303 17586
rect 5359 17530 5427 17586
rect 5483 17530 5551 17586
rect 5607 17530 5675 17586
rect 5731 17530 5799 17586
rect 5855 17530 5923 17586
rect 5979 17530 6047 17586
rect 6103 17530 6171 17586
rect 6227 17530 6237 17586
rect 4425 17462 6237 17530
rect 4425 17406 4435 17462
rect 4491 17406 4559 17462
rect 4615 17406 4683 17462
rect 4739 17406 4807 17462
rect 4863 17406 4931 17462
rect 4987 17406 5055 17462
rect 5111 17406 5179 17462
rect 5235 17406 5303 17462
rect 5359 17406 5427 17462
rect 5483 17406 5551 17462
rect 5607 17406 5675 17462
rect 5731 17406 5799 17462
rect 5855 17406 5923 17462
rect 5979 17406 6047 17462
rect 6103 17406 6171 17462
rect 6227 17406 6237 17462
rect 4425 17338 6237 17406
rect 4425 17282 4435 17338
rect 4491 17282 4559 17338
rect 4615 17282 4683 17338
rect 4739 17282 4807 17338
rect 4863 17282 4931 17338
rect 4987 17282 5055 17338
rect 5111 17282 5179 17338
rect 5235 17282 5303 17338
rect 5359 17282 5427 17338
rect 5483 17282 5551 17338
rect 5607 17282 5675 17338
rect 5731 17282 5799 17338
rect 5855 17282 5923 17338
rect 5979 17282 6047 17338
rect 6103 17282 6171 17338
rect 6227 17282 6237 17338
rect 4425 17214 6237 17282
rect 4425 17158 4435 17214
rect 4491 17158 4559 17214
rect 4615 17158 4683 17214
rect 4739 17158 4807 17214
rect 4863 17158 4931 17214
rect 4987 17158 5055 17214
rect 5111 17158 5179 17214
rect 5235 17158 5303 17214
rect 5359 17158 5427 17214
rect 5483 17158 5551 17214
rect 5607 17158 5675 17214
rect 5731 17158 5799 17214
rect 5855 17158 5923 17214
rect 5979 17158 6047 17214
rect 6103 17158 6171 17214
rect 6227 17158 6237 17214
rect 4425 17090 6237 17158
rect 4425 17034 4435 17090
rect 4491 17034 4559 17090
rect 4615 17034 4683 17090
rect 4739 17034 4807 17090
rect 4863 17034 4931 17090
rect 4987 17034 5055 17090
rect 5111 17034 5179 17090
rect 5235 17034 5303 17090
rect 5359 17034 5427 17090
rect 5483 17034 5551 17090
rect 5607 17034 5675 17090
rect 5731 17034 5799 17090
rect 5855 17034 5923 17090
rect 5979 17034 6047 17090
rect 6103 17034 6171 17090
rect 6227 17034 6237 17090
rect 4425 16966 6237 17034
rect 4425 16910 4435 16966
rect 4491 16910 4559 16966
rect 4615 16910 4683 16966
rect 4739 16910 4807 16966
rect 4863 16910 4931 16966
rect 4987 16910 5055 16966
rect 5111 16910 5179 16966
rect 5235 16910 5303 16966
rect 5359 16910 5427 16966
rect 5483 16910 5551 16966
rect 5607 16910 5675 16966
rect 5731 16910 5799 16966
rect 5855 16910 5923 16966
rect 5979 16910 6047 16966
rect 6103 16910 6171 16966
rect 6227 16910 6237 16966
rect 4425 16842 6237 16910
rect 4425 16786 4435 16842
rect 4491 16786 4559 16842
rect 4615 16786 4683 16842
rect 4739 16786 4807 16842
rect 4863 16786 4931 16842
rect 4987 16786 5055 16842
rect 5111 16786 5179 16842
rect 5235 16786 5303 16842
rect 5359 16786 5427 16842
rect 5483 16786 5551 16842
rect 5607 16786 5675 16842
rect 5731 16786 5799 16842
rect 5855 16786 5923 16842
rect 5979 16786 6047 16842
rect 6103 16786 6171 16842
rect 6227 16786 6237 16842
rect 4425 16718 6237 16786
rect 4425 16662 4435 16718
rect 4491 16662 4559 16718
rect 4615 16662 4683 16718
rect 4739 16662 4807 16718
rect 4863 16662 4931 16718
rect 4987 16662 5055 16718
rect 5111 16662 5179 16718
rect 5235 16662 5303 16718
rect 5359 16662 5427 16718
rect 5483 16662 5551 16718
rect 5607 16662 5675 16718
rect 5731 16662 5799 16718
rect 5855 16662 5923 16718
rect 5979 16662 6047 16718
rect 6103 16662 6171 16718
rect 6227 16662 6237 16718
rect 4425 16594 6237 16662
rect 4425 16538 4435 16594
rect 4491 16538 4559 16594
rect 4615 16538 4683 16594
rect 4739 16538 4807 16594
rect 4863 16538 4931 16594
rect 4987 16538 5055 16594
rect 5111 16538 5179 16594
rect 5235 16538 5303 16594
rect 5359 16538 5427 16594
rect 5483 16538 5551 16594
rect 5607 16538 5675 16594
rect 5731 16538 5799 16594
rect 5855 16538 5923 16594
rect 5979 16538 6047 16594
rect 6103 16538 6171 16594
rect 6227 16538 6237 16594
rect 4425 16470 6237 16538
rect 4425 16414 4435 16470
rect 4491 16414 4559 16470
rect 4615 16414 4683 16470
rect 4739 16414 4807 16470
rect 4863 16414 4931 16470
rect 4987 16414 5055 16470
rect 5111 16414 5179 16470
rect 5235 16414 5303 16470
rect 5359 16414 5427 16470
rect 5483 16414 5551 16470
rect 5607 16414 5675 16470
rect 5731 16414 5799 16470
rect 5855 16414 5923 16470
rect 5979 16414 6047 16470
rect 6103 16414 6171 16470
rect 6227 16414 6237 16470
rect 4425 16346 6237 16414
rect 4425 16290 4435 16346
rect 4491 16290 4559 16346
rect 4615 16290 4683 16346
rect 4739 16290 4807 16346
rect 4863 16290 4931 16346
rect 4987 16290 5055 16346
rect 5111 16290 5179 16346
rect 5235 16290 5303 16346
rect 5359 16290 5427 16346
rect 5483 16290 5551 16346
rect 5607 16290 5675 16346
rect 5731 16290 5799 16346
rect 5855 16290 5923 16346
rect 5979 16290 6047 16346
rect 6103 16290 6171 16346
rect 6227 16290 6237 16346
rect 4425 16222 6237 16290
rect 4425 16166 4435 16222
rect 4491 16166 4559 16222
rect 4615 16166 4683 16222
rect 4739 16166 4807 16222
rect 4863 16166 4931 16222
rect 4987 16166 5055 16222
rect 5111 16166 5179 16222
rect 5235 16166 5303 16222
rect 5359 16166 5427 16222
rect 5483 16166 5551 16222
rect 5607 16166 5675 16222
rect 5731 16166 5799 16222
rect 5855 16166 5923 16222
rect 5979 16166 6047 16222
rect 6103 16166 6171 16222
rect 6227 16166 6237 16222
rect 4425 16098 6237 16166
rect 4425 16042 4435 16098
rect 4491 16042 4559 16098
rect 4615 16042 4683 16098
rect 4739 16042 4807 16098
rect 4863 16042 4931 16098
rect 4987 16042 5055 16098
rect 5111 16042 5179 16098
rect 5235 16042 5303 16098
rect 5359 16042 5427 16098
rect 5483 16042 5551 16098
rect 5607 16042 5675 16098
rect 5731 16042 5799 16098
rect 5855 16042 5923 16098
rect 5979 16042 6047 16098
rect 6103 16042 6171 16098
rect 6227 16042 6237 16098
rect 4425 16032 6237 16042
rect 7552 18950 8620 18960
rect 7552 18894 7562 18950
rect 7618 18894 7686 18950
rect 7742 18894 7810 18950
rect 7866 18894 7934 18950
rect 7990 18894 8058 18950
rect 8114 18894 8182 18950
rect 8238 18894 8306 18950
rect 8362 18894 8430 18950
rect 8486 18894 8554 18950
rect 8610 18894 8620 18950
rect 7552 18826 8620 18894
rect 7552 18770 7562 18826
rect 7618 18770 7686 18826
rect 7742 18770 7810 18826
rect 7866 18770 7934 18826
rect 7990 18770 8058 18826
rect 8114 18770 8182 18826
rect 8238 18770 8306 18826
rect 8362 18770 8430 18826
rect 8486 18770 8554 18826
rect 8610 18770 8620 18826
rect 7552 18702 8620 18770
rect 7552 18646 7562 18702
rect 7618 18646 7686 18702
rect 7742 18646 7810 18702
rect 7866 18646 7934 18702
rect 7990 18646 8058 18702
rect 8114 18646 8182 18702
rect 8238 18646 8306 18702
rect 8362 18646 8430 18702
rect 8486 18646 8554 18702
rect 8610 18646 8620 18702
rect 7552 18578 8620 18646
rect 7552 18522 7562 18578
rect 7618 18522 7686 18578
rect 7742 18522 7810 18578
rect 7866 18522 7934 18578
rect 7990 18522 8058 18578
rect 8114 18522 8182 18578
rect 8238 18522 8306 18578
rect 8362 18522 8430 18578
rect 8486 18522 8554 18578
rect 8610 18522 8620 18578
rect 7552 18454 8620 18522
rect 7552 18398 7562 18454
rect 7618 18398 7686 18454
rect 7742 18398 7810 18454
rect 7866 18398 7934 18454
rect 7990 18398 8058 18454
rect 8114 18398 8182 18454
rect 8238 18398 8306 18454
rect 8362 18398 8430 18454
rect 8486 18398 8554 18454
rect 8610 18398 8620 18454
rect 7552 18330 8620 18398
rect 7552 18274 7562 18330
rect 7618 18274 7686 18330
rect 7742 18274 7810 18330
rect 7866 18274 7934 18330
rect 7990 18274 8058 18330
rect 8114 18274 8182 18330
rect 8238 18274 8306 18330
rect 8362 18274 8430 18330
rect 8486 18274 8554 18330
rect 8610 18274 8620 18330
rect 7552 18206 8620 18274
rect 7552 18150 7562 18206
rect 7618 18150 7686 18206
rect 7742 18150 7810 18206
rect 7866 18150 7934 18206
rect 7990 18150 8058 18206
rect 8114 18150 8182 18206
rect 8238 18150 8306 18206
rect 8362 18150 8430 18206
rect 8486 18150 8554 18206
rect 8610 18150 8620 18206
rect 7552 18082 8620 18150
rect 7552 18026 7562 18082
rect 7618 18026 7686 18082
rect 7742 18026 7810 18082
rect 7866 18026 7934 18082
rect 7990 18026 8058 18082
rect 8114 18026 8182 18082
rect 8238 18026 8306 18082
rect 8362 18026 8430 18082
rect 8486 18026 8554 18082
rect 8610 18026 8620 18082
rect 7552 17958 8620 18026
rect 7552 17902 7562 17958
rect 7618 17902 7686 17958
rect 7742 17902 7810 17958
rect 7866 17902 7934 17958
rect 7990 17902 8058 17958
rect 8114 17902 8182 17958
rect 8238 17902 8306 17958
rect 8362 17902 8430 17958
rect 8486 17902 8554 17958
rect 8610 17902 8620 17958
rect 7552 17834 8620 17902
rect 7552 17778 7562 17834
rect 7618 17778 7686 17834
rect 7742 17778 7810 17834
rect 7866 17778 7934 17834
rect 7990 17778 8058 17834
rect 8114 17778 8182 17834
rect 8238 17778 8306 17834
rect 8362 17778 8430 17834
rect 8486 17778 8554 17834
rect 8610 17778 8620 17834
rect 7552 17710 8620 17778
rect 7552 17654 7562 17710
rect 7618 17654 7686 17710
rect 7742 17654 7810 17710
rect 7866 17654 7934 17710
rect 7990 17654 8058 17710
rect 8114 17654 8182 17710
rect 8238 17654 8306 17710
rect 8362 17654 8430 17710
rect 8486 17654 8554 17710
rect 8610 17654 8620 17710
rect 7552 17586 8620 17654
rect 7552 17530 7562 17586
rect 7618 17530 7686 17586
rect 7742 17530 7810 17586
rect 7866 17530 7934 17586
rect 7990 17530 8058 17586
rect 8114 17530 8182 17586
rect 8238 17530 8306 17586
rect 8362 17530 8430 17586
rect 8486 17530 8554 17586
rect 8610 17530 8620 17586
rect 7552 17462 8620 17530
rect 7552 17406 7562 17462
rect 7618 17406 7686 17462
rect 7742 17406 7810 17462
rect 7866 17406 7934 17462
rect 7990 17406 8058 17462
rect 8114 17406 8182 17462
rect 8238 17406 8306 17462
rect 8362 17406 8430 17462
rect 8486 17406 8554 17462
rect 8610 17406 8620 17462
rect 7552 17338 8620 17406
rect 7552 17282 7562 17338
rect 7618 17282 7686 17338
rect 7742 17282 7810 17338
rect 7866 17282 7934 17338
rect 7990 17282 8058 17338
rect 8114 17282 8182 17338
rect 8238 17282 8306 17338
rect 8362 17282 8430 17338
rect 8486 17282 8554 17338
rect 8610 17282 8620 17338
rect 7552 17214 8620 17282
rect 7552 17158 7562 17214
rect 7618 17158 7686 17214
rect 7742 17158 7810 17214
rect 7866 17158 7934 17214
rect 7990 17158 8058 17214
rect 8114 17158 8182 17214
rect 8238 17158 8306 17214
rect 8362 17158 8430 17214
rect 8486 17158 8554 17214
rect 8610 17158 8620 17214
rect 7552 17090 8620 17158
rect 7552 17034 7562 17090
rect 7618 17034 7686 17090
rect 7742 17034 7810 17090
rect 7866 17034 7934 17090
rect 7990 17034 8058 17090
rect 8114 17034 8182 17090
rect 8238 17034 8306 17090
rect 8362 17034 8430 17090
rect 8486 17034 8554 17090
rect 8610 17034 8620 17090
rect 7552 16966 8620 17034
rect 7552 16910 7562 16966
rect 7618 16910 7686 16966
rect 7742 16910 7810 16966
rect 7866 16910 7934 16966
rect 7990 16910 8058 16966
rect 8114 16910 8182 16966
rect 8238 16910 8306 16966
rect 8362 16910 8430 16966
rect 8486 16910 8554 16966
rect 8610 16910 8620 16966
rect 7552 16842 8620 16910
rect 7552 16786 7562 16842
rect 7618 16786 7686 16842
rect 7742 16786 7810 16842
rect 7866 16786 7934 16842
rect 7990 16786 8058 16842
rect 8114 16786 8182 16842
rect 8238 16786 8306 16842
rect 8362 16786 8430 16842
rect 8486 16786 8554 16842
rect 8610 16786 8620 16842
rect 7552 16718 8620 16786
rect 7552 16662 7562 16718
rect 7618 16662 7686 16718
rect 7742 16662 7810 16718
rect 7866 16662 7934 16718
rect 7990 16662 8058 16718
rect 8114 16662 8182 16718
rect 8238 16662 8306 16718
rect 8362 16662 8430 16718
rect 8486 16662 8554 16718
rect 8610 16662 8620 16718
rect 7552 16594 8620 16662
rect 7552 16538 7562 16594
rect 7618 16538 7686 16594
rect 7742 16538 7810 16594
rect 7866 16538 7934 16594
rect 7990 16538 8058 16594
rect 8114 16538 8182 16594
rect 8238 16538 8306 16594
rect 8362 16538 8430 16594
rect 8486 16538 8554 16594
rect 8610 16538 8620 16594
rect 7552 16470 8620 16538
rect 7552 16414 7562 16470
rect 7618 16414 7686 16470
rect 7742 16414 7810 16470
rect 7866 16414 7934 16470
rect 7990 16414 8058 16470
rect 8114 16414 8182 16470
rect 8238 16414 8306 16470
rect 8362 16414 8430 16470
rect 8486 16414 8554 16470
rect 8610 16414 8620 16470
rect 7552 16346 8620 16414
rect 7552 16290 7562 16346
rect 7618 16290 7686 16346
rect 7742 16290 7810 16346
rect 7866 16290 7934 16346
rect 7990 16290 8058 16346
rect 8114 16290 8182 16346
rect 8238 16290 8306 16346
rect 8362 16290 8430 16346
rect 8486 16290 8554 16346
rect 8610 16290 8620 16346
rect 7552 16222 8620 16290
rect 7552 16166 7562 16222
rect 7618 16166 7686 16222
rect 7742 16166 7810 16222
rect 7866 16166 7934 16222
rect 7990 16166 8058 16222
rect 8114 16166 8182 16222
rect 8238 16166 8306 16222
rect 8362 16166 8430 16222
rect 8486 16166 8554 16222
rect 8610 16166 8620 16222
rect 7552 16098 8620 16166
rect 7552 16042 7562 16098
rect 7618 16042 7686 16098
rect 7742 16042 7810 16098
rect 7866 16042 7934 16098
rect 7990 16042 8058 16098
rect 8114 16042 8182 16098
rect 8238 16042 8306 16098
rect 8362 16042 8430 16098
rect 8486 16042 8554 16098
rect 8610 16042 8620 16098
rect 7552 16032 8620 16042
rect 10669 18950 12481 18960
rect 10669 18894 10679 18950
rect 10735 18894 10803 18950
rect 10859 18894 10927 18950
rect 10983 18894 11051 18950
rect 11107 18894 11175 18950
rect 11231 18894 11299 18950
rect 11355 18894 11423 18950
rect 11479 18894 11547 18950
rect 11603 18894 11671 18950
rect 11727 18894 11795 18950
rect 11851 18894 11919 18950
rect 11975 18894 12043 18950
rect 12099 18894 12167 18950
rect 12223 18894 12291 18950
rect 12347 18894 12415 18950
rect 12471 18894 12481 18950
rect 10669 18826 12481 18894
rect 10669 18770 10679 18826
rect 10735 18770 10803 18826
rect 10859 18770 10927 18826
rect 10983 18770 11051 18826
rect 11107 18770 11175 18826
rect 11231 18770 11299 18826
rect 11355 18770 11423 18826
rect 11479 18770 11547 18826
rect 11603 18770 11671 18826
rect 11727 18770 11795 18826
rect 11851 18770 11919 18826
rect 11975 18770 12043 18826
rect 12099 18770 12167 18826
rect 12223 18770 12291 18826
rect 12347 18770 12415 18826
rect 12471 18770 12481 18826
rect 10669 18702 12481 18770
rect 10669 18646 10679 18702
rect 10735 18646 10803 18702
rect 10859 18646 10927 18702
rect 10983 18646 11051 18702
rect 11107 18646 11175 18702
rect 11231 18646 11299 18702
rect 11355 18646 11423 18702
rect 11479 18646 11547 18702
rect 11603 18646 11671 18702
rect 11727 18646 11795 18702
rect 11851 18646 11919 18702
rect 11975 18646 12043 18702
rect 12099 18646 12167 18702
rect 12223 18646 12291 18702
rect 12347 18646 12415 18702
rect 12471 18646 12481 18702
rect 10669 18578 12481 18646
rect 10669 18522 10679 18578
rect 10735 18522 10803 18578
rect 10859 18522 10927 18578
rect 10983 18522 11051 18578
rect 11107 18522 11175 18578
rect 11231 18522 11299 18578
rect 11355 18522 11423 18578
rect 11479 18522 11547 18578
rect 11603 18522 11671 18578
rect 11727 18522 11795 18578
rect 11851 18522 11919 18578
rect 11975 18522 12043 18578
rect 12099 18522 12167 18578
rect 12223 18522 12291 18578
rect 12347 18522 12415 18578
rect 12471 18522 12481 18578
rect 10669 18454 12481 18522
rect 10669 18398 10679 18454
rect 10735 18398 10803 18454
rect 10859 18398 10927 18454
rect 10983 18398 11051 18454
rect 11107 18398 11175 18454
rect 11231 18398 11299 18454
rect 11355 18398 11423 18454
rect 11479 18398 11547 18454
rect 11603 18398 11671 18454
rect 11727 18398 11795 18454
rect 11851 18398 11919 18454
rect 11975 18398 12043 18454
rect 12099 18398 12167 18454
rect 12223 18398 12291 18454
rect 12347 18398 12415 18454
rect 12471 18398 12481 18454
rect 10669 18330 12481 18398
rect 10669 18274 10679 18330
rect 10735 18274 10803 18330
rect 10859 18274 10927 18330
rect 10983 18274 11051 18330
rect 11107 18274 11175 18330
rect 11231 18274 11299 18330
rect 11355 18274 11423 18330
rect 11479 18274 11547 18330
rect 11603 18274 11671 18330
rect 11727 18274 11795 18330
rect 11851 18274 11919 18330
rect 11975 18274 12043 18330
rect 12099 18274 12167 18330
rect 12223 18274 12291 18330
rect 12347 18274 12415 18330
rect 12471 18274 12481 18330
rect 10669 18206 12481 18274
rect 10669 18150 10679 18206
rect 10735 18150 10803 18206
rect 10859 18150 10927 18206
rect 10983 18150 11051 18206
rect 11107 18150 11175 18206
rect 11231 18150 11299 18206
rect 11355 18150 11423 18206
rect 11479 18150 11547 18206
rect 11603 18150 11671 18206
rect 11727 18150 11795 18206
rect 11851 18150 11919 18206
rect 11975 18150 12043 18206
rect 12099 18150 12167 18206
rect 12223 18150 12291 18206
rect 12347 18150 12415 18206
rect 12471 18150 12481 18206
rect 10669 18082 12481 18150
rect 10669 18026 10679 18082
rect 10735 18026 10803 18082
rect 10859 18026 10927 18082
rect 10983 18026 11051 18082
rect 11107 18026 11175 18082
rect 11231 18026 11299 18082
rect 11355 18026 11423 18082
rect 11479 18026 11547 18082
rect 11603 18026 11671 18082
rect 11727 18026 11795 18082
rect 11851 18026 11919 18082
rect 11975 18026 12043 18082
rect 12099 18026 12167 18082
rect 12223 18026 12291 18082
rect 12347 18026 12415 18082
rect 12471 18026 12481 18082
rect 10669 17958 12481 18026
rect 10669 17902 10679 17958
rect 10735 17902 10803 17958
rect 10859 17902 10927 17958
rect 10983 17902 11051 17958
rect 11107 17902 11175 17958
rect 11231 17902 11299 17958
rect 11355 17902 11423 17958
rect 11479 17902 11547 17958
rect 11603 17902 11671 17958
rect 11727 17902 11795 17958
rect 11851 17902 11919 17958
rect 11975 17902 12043 17958
rect 12099 17902 12167 17958
rect 12223 17902 12291 17958
rect 12347 17902 12415 17958
rect 12471 17902 12481 17958
rect 10669 17834 12481 17902
rect 10669 17778 10679 17834
rect 10735 17778 10803 17834
rect 10859 17778 10927 17834
rect 10983 17778 11051 17834
rect 11107 17778 11175 17834
rect 11231 17778 11299 17834
rect 11355 17778 11423 17834
rect 11479 17778 11547 17834
rect 11603 17778 11671 17834
rect 11727 17778 11795 17834
rect 11851 17778 11919 17834
rect 11975 17778 12043 17834
rect 12099 17778 12167 17834
rect 12223 17778 12291 17834
rect 12347 17778 12415 17834
rect 12471 17778 12481 17834
rect 10669 17710 12481 17778
rect 10669 17654 10679 17710
rect 10735 17654 10803 17710
rect 10859 17654 10927 17710
rect 10983 17654 11051 17710
rect 11107 17654 11175 17710
rect 11231 17654 11299 17710
rect 11355 17654 11423 17710
rect 11479 17654 11547 17710
rect 11603 17654 11671 17710
rect 11727 17654 11795 17710
rect 11851 17654 11919 17710
rect 11975 17654 12043 17710
rect 12099 17654 12167 17710
rect 12223 17654 12291 17710
rect 12347 17654 12415 17710
rect 12471 17654 12481 17710
rect 10669 17586 12481 17654
rect 10669 17530 10679 17586
rect 10735 17530 10803 17586
rect 10859 17530 10927 17586
rect 10983 17530 11051 17586
rect 11107 17530 11175 17586
rect 11231 17530 11299 17586
rect 11355 17530 11423 17586
rect 11479 17530 11547 17586
rect 11603 17530 11671 17586
rect 11727 17530 11795 17586
rect 11851 17530 11919 17586
rect 11975 17530 12043 17586
rect 12099 17530 12167 17586
rect 12223 17530 12291 17586
rect 12347 17530 12415 17586
rect 12471 17530 12481 17586
rect 10669 17462 12481 17530
rect 10669 17406 10679 17462
rect 10735 17406 10803 17462
rect 10859 17406 10927 17462
rect 10983 17406 11051 17462
rect 11107 17406 11175 17462
rect 11231 17406 11299 17462
rect 11355 17406 11423 17462
rect 11479 17406 11547 17462
rect 11603 17406 11671 17462
rect 11727 17406 11795 17462
rect 11851 17406 11919 17462
rect 11975 17406 12043 17462
rect 12099 17406 12167 17462
rect 12223 17406 12291 17462
rect 12347 17406 12415 17462
rect 12471 17406 12481 17462
rect 10669 17338 12481 17406
rect 10669 17282 10679 17338
rect 10735 17282 10803 17338
rect 10859 17282 10927 17338
rect 10983 17282 11051 17338
rect 11107 17282 11175 17338
rect 11231 17282 11299 17338
rect 11355 17282 11423 17338
rect 11479 17282 11547 17338
rect 11603 17282 11671 17338
rect 11727 17282 11795 17338
rect 11851 17282 11919 17338
rect 11975 17282 12043 17338
rect 12099 17282 12167 17338
rect 12223 17282 12291 17338
rect 12347 17282 12415 17338
rect 12471 17282 12481 17338
rect 10669 17214 12481 17282
rect 10669 17158 10679 17214
rect 10735 17158 10803 17214
rect 10859 17158 10927 17214
rect 10983 17158 11051 17214
rect 11107 17158 11175 17214
rect 11231 17158 11299 17214
rect 11355 17158 11423 17214
rect 11479 17158 11547 17214
rect 11603 17158 11671 17214
rect 11727 17158 11795 17214
rect 11851 17158 11919 17214
rect 11975 17158 12043 17214
rect 12099 17158 12167 17214
rect 12223 17158 12291 17214
rect 12347 17158 12415 17214
rect 12471 17158 12481 17214
rect 10669 17090 12481 17158
rect 10669 17034 10679 17090
rect 10735 17034 10803 17090
rect 10859 17034 10927 17090
rect 10983 17034 11051 17090
rect 11107 17034 11175 17090
rect 11231 17034 11299 17090
rect 11355 17034 11423 17090
rect 11479 17034 11547 17090
rect 11603 17034 11671 17090
rect 11727 17034 11795 17090
rect 11851 17034 11919 17090
rect 11975 17034 12043 17090
rect 12099 17034 12167 17090
rect 12223 17034 12291 17090
rect 12347 17034 12415 17090
rect 12471 17034 12481 17090
rect 10669 16966 12481 17034
rect 10669 16910 10679 16966
rect 10735 16910 10803 16966
rect 10859 16910 10927 16966
rect 10983 16910 11051 16966
rect 11107 16910 11175 16966
rect 11231 16910 11299 16966
rect 11355 16910 11423 16966
rect 11479 16910 11547 16966
rect 11603 16910 11671 16966
rect 11727 16910 11795 16966
rect 11851 16910 11919 16966
rect 11975 16910 12043 16966
rect 12099 16910 12167 16966
rect 12223 16910 12291 16966
rect 12347 16910 12415 16966
rect 12471 16910 12481 16966
rect 10669 16842 12481 16910
rect 10669 16786 10679 16842
rect 10735 16786 10803 16842
rect 10859 16786 10927 16842
rect 10983 16786 11051 16842
rect 11107 16786 11175 16842
rect 11231 16786 11299 16842
rect 11355 16786 11423 16842
rect 11479 16786 11547 16842
rect 11603 16786 11671 16842
rect 11727 16786 11795 16842
rect 11851 16786 11919 16842
rect 11975 16786 12043 16842
rect 12099 16786 12167 16842
rect 12223 16786 12291 16842
rect 12347 16786 12415 16842
rect 12471 16786 12481 16842
rect 10669 16718 12481 16786
rect 10669 16662 10679 16718
rect 10735 16662 10803 16718
rect 10859 16662 10927 16718
rect 10983 16662 11051 16718
rect 11107 16662 11175 16718
rect 11231 16662 11299 16718
rect 11355 16662 11423 16718
rect 11479 16662 11547 16718
rect 11603 16662 11671 16718
rect 11727 16662 11795 16718
rect 11851 16662 11919 16718
rect 11975 16662 12043 16718
rect 12099 16662 12167 16718
rect 12223 16662 12291 16718
rect 12347 16662 12415 16718
rect 12471 16662 12481 16718
rect 10669 16594 12481 16662
rect 10669 16538 10679 16594
rect 10735 16538 10803 16594
rect 10859 16538 10927 16594
rect 10983 16538 11051 16594
rect 11107 16538 11175 16594
rect 11231 16538 11299 16594
rect 11355 16538 11423 16594
rect 11479 16538 11547 16594
rect 11603 16538 11671 16594
rect 11727 16538 11795 16594
rect 11851 16538 11919 16594
rect 11975 16538 12043 16594
rect 12099 16538 12167 16594
rect 12223 16538 12291 16594
rect 12347 16538 12415 16594
rect 12471 16538 12481 16594
rect 10669 16470 12481 16538
rect 10669 16414 10679 16470
rect 10735 16414 10803 16470
rect 10859 16414 10927 16470
rect 10983 16414 11051 16470
rect 11107 16414 11175 16470
rect 11231 16414 11299 16470
rect 11355 16414 11423 16470
rect 11479 16414 11547 16470
rect 11603 16414 11671 16470
rect 11727 16414 11795 16470
rect 11851 16414 11919 16470
rect 11975 16414 12043 16470
rect 12099 16414 12167 16470
rect 12223 16414 12291 16470
rect 12347 16414 12415 16470
rect 12471 16414 12481 16470
rect 10669 16346 12481 16414
rect 10669 16290 10679 16346
rect 10735 16290 10803 16346
rect 10859 16290 10927 16346
rect 10983 16290 11051 16346
rect 11107 16290 11175 16346
rect 11231 16290 11299 16346
rect 11355 16290 11423 16346
rect 11479 16290 11547 16346
rect 11603 16290 11671 16346
rect 11727 16290 11795 16346
rect 11851 16290 11919 16346
rect 11975 16290 12043 16346
rect 12099 16290 12167 16346
rect 12223 16290 12291 16346
rect 12347 16290 12415 16346
rect 12471 16290 12481 16346
rect 10669 16222 12481 16290
rect 10669 16166 10679 16222
rect 10735 16166 10803 16222
rect 10859 16166 10927 16222
rect 10983 16166 11051 16222
rect 11107 16166 11175 16222
rect 11231 16166 11299 16222
rect 11355 16166 11423 16222
rect 11479 16166 11547 16222
rect 11603 16166 11671 16222
rect 11727 16166 11795 16222
rect 11851 16166 11919 16222
rect 11975 16166 12043 16222
rect 12099 16166 12167 16222
rect 12223 16166 12291 16222
rect 12347 16166 12415 16222
rect 12471 16166 12481 16222
rect 10669 16098 12481 16166
rect 10669 16042 10679 16098
rect 10735 16042 10803 16098
rect 10859 16042 10927 16098
rect 10983 16042 11051 16098
rect 11107 16042 11175 16098
rect 11231 16042 11299 16098
rect 11355 16042 11423 16098
rect 11479 16042 11547 16098
rect 11603 16042 11671 16098
rect 11727 16042 11795 16098
rect 11851 16042 11919 16098
rect 11975 16042 12043 16098
rect 12099 16042 12167 16098
rect 12223 16042 12291 16098
rect 12347 16042 12415 16098
rect 12471 16042 12481 16098
rect 10669 16032 12481 16042
rect 1068 15750 2136 15760
rect 1068 15694 1078 15750
rect 1134 15694 1202 15750
rect 1258 15694 1326 15750
rect 1382 15694 1450 15750
rect 1506 15694 1574 15750
rect 1630 15694 1698 15750
rect 1754 15694 1822 15750
rect 1878 15694 1946 15750
rect 2002 15694 2070 15750
rect 2126 15694 2136 15750
rect 1068 15626 2136 15694
rect 1068 15570 1078 15626
rect 1134 15570 1202 15626
rect 1258 15570 1326 15626
rect 1382 15570 1450 15626
rect 1506 15570 1574 15626
rect 1630 15570 1698 15626
rect 1754 15570 1822 15626
rect 1878 15570 1946 15626
rect 2002 15570 2070 15626
rect 2126 15570 2136 15626
rect 1068 15502 2136 15570
rect 1068 15446 1078 15502
rect 1134 15446 1202 15502
rect 1258 15446 1326 15502
rect 1382 15446 1450 15502
rect 1506 15446 1574 15502
rect 1630 15446 1698 15502
rect 1754 15446 1822 15502
rect 1878 15446 1946 15502
rect 2002 15446 2070 15502
rect 2126 15446 2136 15502
rect 1068 15378 2136 15446
rect 1068 15322 1078 15378
rect 1134 15322 1202 15378
rect 1258 15322 1326 15378
rect 1382 15322 1450 15378
rect 1506 15322 1574 15378
rect 1630 15322 1698 15378
rect 1754 15322 1822 15378
rect 1878 15322 1946 15378
rect 2002 15322 2070 15378
rect 2126 15322 2136 15378
rect 1068 15254 2136 15322
rect 1068 15198 1078 15254
rect 1134 15198 1202 15254
rect 1258 15198 1326 15254
rect 1382 15198 1450 15254
rect 1506 15198 1574 15254
rect 1630 15198 1698 15254
rect 1754 15198 1822 15254
rect 1878 15198 1946 15254
rect 2002 15198 2070 15254
rect 2126 15198 2136 15254
rect 1068 15130 2136 15198
rect 1068 15074 1078 15130
rect 1134 15074 1202 15130
rect 1258 15074 1326 15130
rect 1382 15074 1450 15130
rect 1506 15074 1574 15130
rect 1630 15074 1698 15130
rect 1754 15074 1822 15130
rect 1878 15074 1946 15130
rect 2002 15074 2070 15130
rect 2126 15074 2136 15130
rect 1068 15006 2136 15074
rect 1068 14950 1078 15006
rect 1134 14950 1202 15006
rect 1258 14950 1326 15006
rect 1382 14950 1450 15006
rect 1506 14950 1574 15006
rect 1630 14950 1698 15006
rect 1754 14950 1822 15006
rect 1878 14950 1946 15006
rect 2002 14950 2070 15006
rect 2126 14950 2136 15006
rect 1068 14882 2136 14950
rect 1068 14826 1078 14882
rect 1134 14826 1202 14882
rect 1258 14826 1326 14882
rect 1382 14826 1450 14882
rect 1506 14826 1574 14882
rect 1630 14826 1698 14882
rect 1754 14826 1822 14882
rect 1878 14826 1946 14882
rect 2002 14826 2070 14882
rect 2126 14826 2136 14882
rect 1068 14758 2136 14826
rect 1068 14702 1078 14758
rect 1134 14702 1202 14758
rect 1258 14702 1326 14758
rect 1382 14702 1450 14758
rect 1506 14702 1574 14758
rect 1630 14702 1698 14758
rect 1754 14702 1822 14758
rect 1878 14702 1946 14758
rect 2002 14702 2070 14758
rect 2126 14702 2136 14758
rect 1068 14634 2136 14702
rect 1068 14578 1078 14634
rect 1134 14578 1202 14634
rect 1258 14578 1326 14634
rect 1382 14578 1450 14634
rect 1506 14578 1574 14634
rect 1630 14578 1698 14634
rect 1754 14578 1822 14634
rect 1878 14578 1946 14634
rect 2002 14578 2070 14634
rect 2126 14578 2136 14634
rect 1068 14510 2136 14578
rect 1068 14454 1078 14510
rect 1134 14454 1202 14510
rect 1258 14454 1326 14510
rect 1382 14454 1450 14510
rect 1506 14454 1574 14510
rect 1630 14454 1698 14510
rect 1754 14454 1822 14510
rect 1878 14454 1946 14510
rect 2002 14454 2070 14510
rect 2126 14454 2136 14510
rect 1068 14386 2136 14454
rect 1068 14330 1078 14386
rect 1134 14330 1202 14386
rect 1258 14330 1326 14386
rect 1382 14330 1450 14386
rect 1506 14330 1574 14386
rect 1630 14330 1698 14386
rect 1754 14330 1822 14386
rect 1878 14330 1946 14386
rect 2002 14330 2070 14386
rect 2126 14330 2136 14386
rect 1068 14262 2136 14330
rect 1068 14206 1078 14262
rect 1134 14206 1202 14262
rect 1258 14206 1326 14262
rect 1382 14206 1450 14262
rect 1506 14206 1574 14262
rect 1630 14206 1698 14262
rect 1754 14206 1822 14262
rect 1878 14206 1946 14262
rect 2002 14206 2070 14262
rect 2126 14206 2136 14262
rect 1068 14138 2136 14206
rect 1068 14082 1078 14138
rect 1134 14082 1202 14138
rect 1258 14082 1326 14138
rect 1382 14082 1450 14138
rect 1506 14082 1574 14138
rect 1630 14082 1698 14138
rect 1754 14082 1822 14138
rect 1878 14082 1946 14138
rect 2002 14082 2070 14138
rect 2126 14082 2136 14138
rect 1068 14014 2136 14082
rect 1068 13958 1078 14014
rect 1134 13958 1202 14014
rect 1258 13958 1326 14014
rect 1382 13958 1450 14014
rect 1506 13958 1574 14014
rect 1630 13958 1698 14014
rect 1754 13958 1822 14014
rect 1878 13958 1946 14014
rect 2002 13958 2070 14014
rect 2126 13958 2136 14014
rect 1068 13890 2136 13958
rect 1068 13834 1078 13890
rect 1134 13834 1202 13890
rect 1258 13834 1326 13890
rect 1382 13834 1450 13890
rect 1506 13834 1574 13890
rect 1630 13834 1698 13890
rect 1754 13834 1822 13890
rect 1878 13834 1946 13890
rect 2002 13834 2070 13890
rect 2126 13834 2136 13890
rect 1068 13766 2136 13834
rect 1068 13710 1078 13766
rect 1134 13710 1202 13766
rect 1258 13710 1326 13766
rect 1382 13710 1450 13766
rect 1506 13710 1574 13766
rect 1630 13710 1698 13766
rect 1754 13710 1822 13766
rect 1878 13710 1946 13766
rect 2002 13710 2070 13766
rect 2126 13710 2136 13766
rect 1068 13642 2136 13710
rect 1068 13586 1078 13642
rect 1134 13586 1202 13642
rect 1258 13586 1326 13642
rect 1382 13586 1450 13642
rect 1506 13586 1574 13642
rect 1630 13586 1698 13642
rect 1754 13586 1822 13642
rect 1878 13586 1946 13642
rect 2002 13586 2070 13642
rect 2126 13586 2136 13642
rect 1068 13518 2136 13586
rect 1068 13462 1078 13518
rect 1134 13462 1202 13518
rect 1258 13462 1326 13518
rect 1382 13462 1450 13518
rect 1506 13462 1574 13518
rect 1630 13462 1698 13518
rect 1754 13462 1822 13518
rect 1878 13462 1946 13518
rect 2002 13462 2070 13518
rect 2126 13462 2136 13518
rect 1068 13394 2136 13462
rect 1068 13338 1078 13394
rect 1134 13338 1202 13394
rect 1258 13338 1326 13394
rect 1382 13338 1450 13394
rect 1506 13338 1574 13394
rect 1630 13338 1698 13394
rect 1754 13338 1822 13394
rect 1878 13338 1946 13394
rect 2002 13338 2070 13394
rect 2126 13338 2136 13394
rect 1068 13270 2136 13338
rect 1068 13214 1078 13270
rect 1134 13214 1202 13270
rect 1258 13214 1326 13270
rect 1382 13214 1450 13270
rect 1506 13214 1574 13270
rect 1630 13214 1698 13270
rect 1754 13214 1822 13270
rect 1878 13214 1946 13270
rect 2002 13214 2070 13270
rect 2126 13214 2136 13270
rect 1068 13146 2136 13214
rect 1068 13090 1078 13146
rect 1134 13090 1202 13146
rect 1258 13090 1326 13146
rect 1382 13090 1450 13146
rect 1506 13090 1574 13146
rect 1630 13090 1698 13146
rect 1754 13090 1822 13146
rect 1878 13090 1946 13146
rect 2002 13090 2070 13146
rect 2126 13090 2136 13146
rect 1068 13022 2136 13090
rect 1068 12966 1078 13022
rect 1134 12966 1202 13022
rect 1258 12966 1326 13022
rect 1382 12966 1450 13022
rect 1506 12966 1574 13022
rect 1630 12966 1698 13022
rect 1754 12966 1822 13022
rect 1878 12966 1946 13022
rect 2002 12966 2070 13022
rect 2126 12966 2136 13022
rect 1068 12898 2136 12966
rect 1068 12842 1078 12898
rect 1134 12842 1202 12898
rect 1258 12842 1326 12898
rect 1382 12842 1450 12898
rect 1506 12842 1574 12898
rect 1630 12842 1698 12898
rect 1754 12842 1822 12898
rect 1878 12842 1946 12898
rect 2002 12842 2070 12898
rect 2126 12842 2136 12898
rect 1068 12832 2136 12842
rect 4425 15750 6237 15760
rect 4425 15694 4435 15750
rect 4491 15694 4559 15750
rect 4615 15694 4683 15750
rect 4739 15694 4807 15750
rect 4863 15694 4931 15750
rect 4987 15694 5055 15750
rect 5111 15694 5179 15750
rect 5235 15694 5303 15750
rect 5359 15694 5427 15750
rect 5483 15694 5551 15750
rect 5607 15694 5675 15750
rect 5731 15694 5799 15750
rect 5855 15694 5923 15750
rect 5979 15694 6047 15750
rect 6103 15694 6171 15750
rect 6227 15694 6237 15750
rect 4425 15626 6237 15694
rect 4425 15570 4435 15626
rect 4491 15570 4559 15626
rect 4615 15570 4683 15626
rect 4739 15570 4807 15626
rect 4863 15570 4931 15626
rect 4987 15570 5055 15626
rect 5111 15570 5179 15626
rect 5235 15570 5303 15626
rect 5359 15570 5427 15626
rect 5483 15570 5551 15626
rect 5607 15570 5675 15626
rect 5731 15570 5799 15626
rect 5855 15570 5923 15626
rect 5979 15570 6047 15626
rect 6103 15570 6171 15626
rect 6227 15570 6237 15626
rect 4425 15502 6237 15570
rect 4425 15446 4435 15502
rect 4491 15446 4559 15502
rect 4615 15446 4683 15502
rect 4739 15446 4807 15502
rect 4863 15446 4931 15502
rect 4987 15446 5055 15502
rect 5111 15446 5179 15502
rect 5235 15446 5303 15502
rect 5359 15446 5427 15502
rect 5483 15446 5551 15502
rect 5607 15446 5675 15502
rect 5731 15446 5799 15502
rect 5855 15446 5923 15502
rect 5979 15446 6047 15502
rect 6103 15446 6171 15502
rect 6227 15446 6237 15502
rect 4425 15378 6237 15446
rect 4425 15322 4435 15378
rect 4491 15322 4559 15378
rect 4615 15322 4683 15378
rect 4739 15322 4807 15378
rect 4863 15322 4931 15378
rect 4987 15322 5055 15378
rect 5111 15322 5179 15378
rect 5235 15322 5303 15378
rect 5359 15322 5427 15378
rect 5483 15322 5551 15378
rect 5607 15322 5675 15378
rect 5731 15322 5799 15378
rect 5855 15322 5923 15378
rect 5979 15322 6047 15378
rect 6103 15322 6171 15378
rect 6227 15322 6237 15378
rect 4425 15254 6237 15322
rect 4425 15198 4435 15254
rect 4491 15198 4559 15254
rect 4615 15198 4683 15254
rect 4739 15198 4807 15254
rect 4863 15198 4931 15254
rect 4987 15198 5055 15254
rect 5111 15198 5179 15254
rect 5235 15198 5303 15254
rect 5359 15198 5427 15254
rect 5483 15198 5551 15254
rect 5607 15198 5675 15254
rect 5731 15198 5799 15254
rect 5855 15198 5923 15254
rect 5979 15198 6047 15254
rect 6103 15198 6171 15254
rect 6227 15198 6237 15254
rect 4425 15130 6237 15198
rect 4425 15074 4435 15130
rect 4491 15074 4559 15130
rect 4615 15074 4683 15130
rect 4739 15074 4807 15130
rect 4863 15074 4931 15130
rect 4987 15074 5055 15130
rect 5111 15074 5179 15130
rect 5235 15074 5303 15130
rect 5359 15074 5427 15130
rect 5483 15074 5551 15130
rect 5607 15074 5675 15130
rect 5731 15074 5799 15130
rect 5855 15074 5923 15130
rect 5979 15074 6047 15130
rect 6103 15074 6171 15130
rect 6227 15074 6237 15130
rect 4425 15006 6237 15074
rect 4425 14950 4435 15006
rect 4491 14950 4559 15006
rect 4615 14950 4683 15006
rect 4739 14950 4807 15006
rect 4863 14950 4931 15006
rect 4987 14950 5055 15006
rect 5111 14950 5179 15006
rect 5235 14950 5303 15006
rect 5359 14950 5427 15006
rect 5483 14950 5551 15006
rect 5607 14950 5675 15006
rect 5731 14950 5799 15006
rect 5855 14950 5923 15006
rect 5979 14950 6047 15006
rect 6103 14950 6171 15006
rect 6227 14950 6237 15006
rect 4425 14882 6237 14950
rect 4425 14826 4435 14882
rect 4491 14826 4559 14882
rect 4615 14826 4683 14882
rect 4739 14826 4807 14882
rect 4863 14826 4931 14882
rect 4987 14826 5055 14882
rect 5111 14826 5179 14882
rect 5235 14826 5303 14882
rect 5359 14826 5427 14882
rect 5483 14826 5551 14882
rect 5607 14826 5675 14882
rect 5731 14826 5799 14882
rect 5855 14826 5923 14882
rect 5979 14826 6047 14882
rect 6103 14826 6171 14882
rect 6227 14826 6237 14882
rect 4425 14758 6237 14826
rect 4425 14702 4435 14758
rect 4491 14702 4559 14758
rect 4615 14702 4683 14758
rect 4739 14702 4807 14758
rect 4863 14702 4931 14758
rect 4987 14702 5055 14758
rect 5111 14702 5179 14758
rect 5235 14702 5303 14758
rect 5359 14702 5427 14758
rect 5483 14702 5551 14758
rect 5607 14702 5675 14758
rect 5731 14702 5799 14758
rect 5855 14702 5923 14758
rect 5979 14702 6047 14758
rect 6103 14702 6171 14758
rect 6227 14702 6237 14758
rect 4425 14634 6237 14702
rect 4425 14578 4435 14634
rect 4491 14578 4559 14634
rect 4615 14578 4683 14634
rect 4739 14578 4807 14634
rect 4863 14578 4931 14634
rect 4987 14578 5055 14634
rect 5111 14578 5179 14634
rect 5235 14578 5303 14634
rect 5359 14578 5427 14634
rect 5483 14578 5551 14634
rect 5607 14578 5675 14634
rect 5731 14578 5799 14634
rect 5855 14578 5923 14634
rect 5979 14578 6047 14634
rect 6103 14578 6171 14634
rect 6227 14578 6237 14634
rect 4425 14510 6237 14578
rect 4425 14454 4435 14510
rect 4491 14454 4559 14510
rect 4615 14454 4683 14510
rect 4739 14454 4807 14510
rect 4863 14454 4931 14510
rect 4987 14454 5055 14510
rect 5111 14454 5179 14510
rect 5235 14454 5303 14510
rect 5359 14454 5427 14510
rect 5483 14454 5551 14510
rect 5607 14454 5675 14510
rect 5731 14454 5799 14510
rect 5855 14454 5923 14510
rect 5979 14454 6047 14510
rect 6103 14454 6171 14510
rect 6227 14454 6237 14510
rect 4425 14386 6237 14454
rect 4425 14330 4435 14386
rect 4491 14330 4559 14386
rect 4615 14330 4683 14386
rect 4739 14330 4807 14386
rect 4863 14330 4931 14386
rect 4987 14330 5055 14386
rect 5111 14330 5179 14386
rect 5235 14330 5303 14386
rect 5359 14330 5427 14386
rect 5483 14330 5551 14386
rect 5607 14330 5675 14386
rect 5731 14330 5799 14386
rect 5855 14330 5923 14386
rect 5979 14330 6047 14386
rect 6103 14330 6171 14386
rect 6227 14330 6237 14386
rect 4425 14262 6237 14330
rect 4425 14206 4435 14262
rect 4491 14206 4559 14262
rect 4615 14206 4683 14262
rect 4739 14206 4807 14262
rect 4863 14206 4931 14262
rect 4987 14206 5055 14262
rect 5111 14206 5179 14262
rect 5235 14206 5303 14262
rect 5359 14206 5427 14262
rect 5483 14206 5551 14262
rect 5607 14206 5675 14262
rect 5731 14206 5799 14262
rect 5855 14206 5923 14262
rect 5979 14206 6047 14262
rect 6103 14206 6171 14262
rect 6227 14206 6237 14262
rect 4425 14138 6237 14206
rect 4425 14082 4435 14138
rect 4491 14082 4559 14138
rect 4615 14082 4683 14138
rect 4739 14082 4807 14138
rect 4863 14082 4931 14138
rect 4987 14082 5055 14138
rect 5111 14082 5179 14138
rect 5235 14082 5303 14138
rect 5359 14082 5427 14138
rect 5483 14082 5551 14138
rect 5607 14082 5675 14138
rect 5731 14082 5799 14138
rect 5855 14082 5923 14138
rect 5979 14082 6047 14138
rect 6103 14082 6171 14138
rect 6227 14082 6237 14138
rect 4425 14014 6237 14082
rect 4425 13958 4435 14014
rect 4491 13958 4559 14014
rect 4615 13958 4683 14014
rect 4739 13958 4807 14014
rect 4863 13958 4931 14014
rect 4987 13958 5055 14014
rect 5111 13958 5179 14014
rect 5235 13958 5303 14014
rect 5359 13958 5427 14014
rect 5483 13958 5551 14014
rect 5607 13958 5675 14014
rect 5731 13958 5799 14014
rect 5855 13958 5923 14014
rect 5979 13958 6047 14014
rect 6103 13958 6171 14014
rect 6227 13958 6237 14014
rect 4425 13890 6237 13958
rect 4425 13834 4435 13890
rect 4491 13834 4559 13890
rect 4615 13834 4683 13890
rect 4739 13834 4807 13890
rect 4863 13834 4931 13890
rect 4987 13834 5055 13890
rect 5111 13834 5179 13890
rect 5235 13834 5303 13890
rect 5359 13834 5427 13890
rect 5483 13834 5551 13890
rect 5607 13834 5675 13890
rect 5731 13834 5799 13890
rect 5855 13834 5923 13890
rect 5979 13834 6047 13890
rect 6103 13834 6171 13890
rect 6227 13834 6237 13890
rect 4425 13766 6237 13834
rect 4425 13710 4435 13766
rect 4491 13710 4559 13766
rect 4615 13710 4683 13766
rect 4739 13710 4807 13766
rect 4863 13710 4931 13766
rect 4987 13710 5055 13766
rect 5111 13710 5179 13766
rect 5235 13710 5303 13766
rect 5359 13710 5427 13766
rect 5483 13710 5551 13766
rect 5607 13710 5675 13766
rect 5731 13710 5799 13766
rect 5855 13710 5923 13766
rect 5979 13710 6047 13766
rect 6103 13710 6171 13766
rect 6227 13710 6237 13766
rect 4425 13642 6237 13710
rect 4425 13586 4435 13642
rect 4491 13586 4559 13642
rect 4615 13586 4683 13642
rect 4739 13586 4807 13642
rect 4863 13586 4931 13642
rect 4987 13586 5055 13642
rect 5111 13586 5179 13642
rect 5235 13586 5303 13642
rect 5359 13586 5427 13642
rect 5483 13586 5551 13642
rect 5607 13586 5675 13642
rect 5731 13586 5799 13642
rect 5855 13586 5923 13642
rect 5979 13586 6047 13642
rect 6103 13586 6171 13642
rect 6227 13586 6237 13642
rect 4425 13518 6237 13586
rect 4425 13462 4435 13518
rect 4491 13462 4559 13518
rect 4615 13462 4683 13518
rect 4739 13462 4807 13518
rect 4863 13462 4931 13518
rect 4987 13462 5055 13518
rect 5111 13462 5179 13518
rect 5235 13462 5303 13518
rect 5359 13462 5427 13518
rect 5483 13462 5551 13518
rect 5607 13462 5675 13518
rect 5731 13462 5799 13518
rect 5855 13462 5923 13518
rect 5979 13462 6047 13518
rect 6103 13462 6171 13518
rect 6227 13462 6237 13518
rect 4425 13394 6237 13462
rect 4425 13338 4435 13394
rect 4491 13338 4559 13394
rect 4615 13338 4683 13394
rect 4739 13338 4807 13394
rect 4863 13338 4931 13394
rect 4987 13338 5055 13394
rect 5111 13338 5179 13394
rect 5235 13338 5303 13394
rect 5359 13338 5427 13394
rect 5483 13338 5551 13394
rect 5607 13338 5675 13394
rect 5731 13338 5799 13394
rect 5855 13338 5923 13394
rect 5979 13338 6047 13394
rect 6103 13338 6171 13394
rect 6227 13338 6237 13394
rect 4425 13270 6237 13338
rect 4425 13214 4435 13270
rect 4491 13214 4559 13270
rect 4615 13214 4683 13270
rect 4739 13214 4807 13270
rect 4863 13214 4931 13270
rect 4987 13214 5055 13270
rect 5111 13214 5179 13270
rect 5235 13214 5303 13270
rect 5359 13214 5427 13270
rect 5483 13214 5551 13270
rect 5607 13214 5675 13270
rect 5731 13214 5799 13270
rect 5855 13214 5923 13270
rect 5979 13214 6047 13270
rect 6103 13214 6171 13270
rect 6227 13214 6237 13270
rect 4425 13146 6237 13214
rect 4425 13090 4435 13146
rect 4491 13090 4559 13146
rect 4615 13090 4683 13146
rect 4739 13090 4807 13146
rect 4863 13090 4931 13146
rect 4987 13090 5055 13146
rect 5111 13090 5179 13146
rect 5235 13090 5303 13146
rect 5359 13090 5427 13146
rect 5483 13090 5551 13146
rect 5607 13090 5675 13146
rect 5731 13090 5799 13146
rect 5855 13090 5923 13146
rect 5979 13090 6047 13146
rect 6103 13090 6171 13146
rect 6227 13090 6237 13146
rect 4425 13022 6237 13090
rect 4425 12966 4435 13022
rect 4491 12966 4559 13022
rect 4615 12966 4683 13022
rect 4739 12966 4807 13022
rect 4863 12966 4931 13022
rect 4987 12966 5055 13022
rect 5111 12966 5179 13022
rect 5235 12966 5303 13022
rect 5359 12966 5427 13022
rect 5483 12966 5551 13022
rect 5607 12966 5675 13022
rect 5731 12966 5799 13022
rect 5855 12966 5923 13022
rect 5979 12966 6047 13022
rect 6103 12966 6171 13022
rect 6227 12966 6237 13022
rect 4425 12898 6237 12966
rect 4425 12842 4435 12898
rect 4491 12842 4559 12898
rect 4615 12842 4683 12898
rect 4739 12842 4807 12898
rect 4863 12842 4931 12898
rect 4987 12842 5055 12898
rect 5111 12842 5179 12898
rect 5235 12842 5303 12898
rect 5359 12842 5427 12898
rect 5483 12842 5551 12898
rect 5607 12842 5675 12898
rect 5731 12842 5799 12898
rect 5855 12842 5923 12898
rect 5979 12842 6047 12898
rect 6103 12842 6171 12898
rect 6227 12842 6237 12898
rect 4425 12832 6237 12842
rect 7552 15750 8620 15760
rect 7552 15694 7562 15750
rect 7618 15694 7686 15750
rect 7742 15694 7810 15750
rect 7866 15694 7934 15750
rect 7990 15694 8058 15750
rect 8114 15694 8182 15750
rect 8238 15694 8306 15750
rect 8362 15694 8430 15750
rect 8486 15694 8554 15750
rect 8610 15694 8620 15750
rect 7552 15626 8620 15694
rect 7552 15570 7562 15626
rect 7618 15570 7686 15626
rect 7742 15570 7810 15626
rect 7866 15570 7934 15626
rect 7990 15570 8058 15626
rect 8114 15570 8182 15626
rect 8238 15570 8306 15626
rect 8362 15570 8430 15626
rect 8486 15570 8554 15626
rect 8610 15570 8620 15626
rect 7552 15502 8620 15570
rect 7552 15446 7562 15502
rect 7618 15446 7686 15502
rect 7742 15446 7810 15502
rect 7866 15446 7934 15502
rect 7990 15446 8058 15502
rect 8114 15446 8182 15502
rect 8238 15446 8306 15502
rect 8362 15446 8430 15502
rect 8486 15446 8554 15502
rect 8610 15446 8620 15502
rect 7552 15378 8620 15446
rect 7552 15322 7562 15378
rect 7618 15322 7686 15378
rect 7742 15322 7810 15378
rect 7866 15322 7934 15378
rect 7990 15322 8058 15378
rect 8114 15322 8182 15378
rect 8238 15322 8306 15378
rect 8362 15322 8430 15378
rect 8486 15322 8554 15378
rect 8610 15322 8620 15378
rect 7552 15254 8620 15322
rect 7552 15198 7562 15254
rect 7618 15198 7686 15254
rect 7742 15198 7810 15254
rect 7866 15198 7934 15254
rect 7990 15198 8058 15254
rect 8114 15198 8182 15254
rect 8238 15198 8306 15254
rect 8362 15198 8430 15254
rect 8486 15198 8554 15254
rect 8610 15198 8620 15254
rect 7552 15130 8620 15198
rect 7552 15074 7562 15130
rect 7618 15074 7686 15130
rect 7742 15074 7810 15130
rect 7866 15074 7934 15130
rect 7990 15074 8058 15130
rect 8114 15074 8182 15130
rect 8238 15074 8306 15130
rect 8362 15074 8430 15130
rect 8486 15074 8554 15130
rect 8610 15074 8620 15130
rect 7552 15006 8620 15074
rect 7552 14950 7562 15006
rect 7618 14950 7686 15006
rect 7742 14950 7810 15006
rect 7866 14950 7934 15006
rect 7990 14950 8058 15006
rect 8114 14950 8182 15006
rect 8238 14950 8306 15006
rect 8362 14950 8430 15006
rect 8486 14950 8554 15006
rect 8610 14950 8620 15006
rect 7552 14882 8620 14950
rect 7552 14826 7562 14882
rect 7618 14826 7686 14882
rect 7742 14826 7810 14882
rect 7866 14826 7934 14882
rect 7990 14826 8058 14882
rect 8114 14826 8182 14882
rect 8238 14826 8306 14882
rect 8362 14826 8430 14882
rect 8486 14826 8554 14882
rect 8610 14826 8620 14882
rect 7552 14758 8620 14826
rect 7552 14702 7562 14758
rect 7618 14702 7686 14758
rect 7742 14702 7810 14758
rect 7866 14702 7934 14758
rect 7990 14702 8058 14758
rect 8114 14702 8182 14758
rect 8238 14702 8306 14758
rect 8362 14702 8430 14758
rect 8486 14702 8554 14758
rect 8610 14702 8620 14758
rect 7552 14634 8620 14702
rect 7552 14578 7562 14634
rect 7618 14578 7686 14634
rect 7742 14578 7810 14634
rect 7866 14578 7934 14634
rect 7990 14578 8058 14634
rect 8114 14578 8182 14634
rect 8238 14578 8306 14634
rect 8362 14578 8430 14634
rect 8486 14578 8554 14634
rect 8610 14578 8620 14634
rect 7552 14510 8620 14578
rect 7552 14454 7562 14510
rect 7618 14454 7686 14510
rect 7742 14454 7810 14510
rect 7866 14454 7934 14510
rect 7990 14454 8058 14510
rect 8114 14454 8182 14510
rect 8238 14454 8306 14510
rect 8362 14454 8430 14510
rect 8486 14454 8554 14510
rect 8610 14454 8620 14510
rect 7552 14386 8620 14454
rect 7552 14330 7562 14386
rect 7618 14330 7686 14386
rect 7742 14330 7810 14386
rect 7866 14330 7934 14386
rect 7990 14330 8058 14386
rect 8114 14330 8182 14386
rect 8238 14330 8306 14386
rect 8362 14330 8430 14386
rect 8486 14330 8554 14386
rect 8610 14330 8620 14386
rect 7552 14262 8620 14330
rect 7552 14206 7562 14262
rect 7618 14206 7686 14262
rect 7742 14206 7810 14262
rect 7866 14206 7934 14262
rect 7990 14206 8058 14262
rect 8114 14206 8182 14262
rect 8238 14206 8306 14262
rect 8362 14206 8430 14262
rect 8486 14206 8554 14262
rect 8610 14206 8620 14262
rect 7552 14138 8620 14206
rect 7552 14082 7562 14138
rect 7618 14082 7686 14138
rect 7742 14082 7810 14138
rect 7866 14082 7934 14138
rect 7990 14082 8058 14138
rect 8114 14082 8182 14138
rect 8238 14082 8306 14138
rect 8362 14082 8430 14138
rect 8486 14082 8554 14138
rect 8610 14082 8620 14138
rect 7552 14014 8620 14082
rect 7552 13958 7562 14014
rect 7618 13958 7686 14014
rect 7742 13958 7810 14014
rect 7866 13958 7934 14014
rect 7990 13958 8058 14014
rect 8114 13958 8182 14014
rect 8238 13958 8306 14014
rect 8362 13958 8430 14014
rect 8486 13958 8554 14014
rect 8610 13958 8620 14014
rect 7552 13890 8620 13958
rect 7552 13834 7562 13890
rect 7618 13834 7686 13890
rect 7742 13834 7810 13890
rect 7866 13834 7934 13890
rect 7990 13834 8058 13890
rect 8114 13834 8182 13890
rect 8238 13834 8306 13890
rect 8362 13834 8430 13890
rect 8486 13834 8554 13890
rect 8610 13834 8620 13890
rect 7552 13766 8620 13834
rect 7552 13710 7562 13766
rect 7618 13710 7686 13766
rect 7742 13710 7810 13766
rect 7866 13710 7934 13766
rect 7990 13710 8058 13766
rect 8114 13710 8182 13766
rect 8238 13710 8306 13766
rect 8362 13710 8430 13766
rect 8486 13710 8554 13766
rect 8610 13710 8620 13766
rect 7552 13642 8620 13710
rect 7552 13586 7562 13642
rect 7618 13586 7686 13642
rect 7742 13586 7810 13642
rect 7866 13586 7934 13642
rect 7990 13586 8058 13642
rect 8114 13586 8182 13642
rect 8238 13586 8306 13642
rect 8362 13586 8430 13642
rect 8486 13586 8554 13642
rect 8610 13586 8620 13642
rect 7552 13518 8620 13586
rect 7552 13462 7562 13518
rect 7618 13462 7686 13518
rect 7742 13462 7810 13518
rect 7866 13462 7934 13518
rect 7990 13462 8058 13518
rect 8114 13462 8182 13518
rect 8238 13462 8306 13518
rect 8362 13462 8430 13518
rect 8486 13462 8554 13518
rect 8610 13462 8620 13518
rect 7552 13394 8620 13462
rect 7552 13338 7562 13394
rect 7618 13338 7686 13394
rect 7742 13338 7810 13394
rect 7866 13338 7934 13394
rect 7990 13338 8058 13394
rect 8114 13338 8182 13394
rect 8238 13338 8306 13394
rect 8362 13338 8430 13394
rect 8486 13338 8554 13394
rect 8610 13338 8620 13394
rect 7552 13270 8620 13338
rect 7552 13214 7562 13270
rect 7618 13214 7686 13270
rect 7742 13214 7810 13270
rect 7866 13214 7934 13270
rect 7990 13214 8058 13270
rect 8114 13214 8182 13270
rect 8238 13214 8306 13270
rect 8362 13214 8430 13270
rect 8486 13214 8554 13270
rect 8610 13214 8620 13270
rect 7552 13146 8620 13214
rect 7552 13090 7562 13146
rect 7618 13090 7686 13146
rect 7742 13090 7810 13146
rect 7866 13090 7934 13146
rect 7990 13090 8058 13146
rect 8114 13090 8182 13146
rect 8238 13090 8306 13146
rect 8362 13090 8430 13146
rect 8486 13090 8554 13146
rect 8610 13090 8620 13146
rect 7552 13022 8620 13090
rect 7552 12966 7562 13022
rect 7618 12966 7686 13022
rect 7742 12966 7810 13022
rect 7866 12966 7934 13022
rect 7990 12966 8058 13022
rect 8114 12966 8182 13022
rect 8238 12966 8306 13022
rect 8362 12966 8430 13022
rect 8486 12966 8554 13022
rect 8610 12966 8620 13022
rect 7552 12898 8620 12966
rect 7552 12842 7562 12898
rect 7618 12842 7686 12898
rect 7742 12842 7810 12898
rect 7866 12842 7934 12898
rect 7990 12842 8058 12898
rect 8114 12842 8182 12898
rect 8238 12842 8306 12898
rect 8362 12842 8430 12898
rect 8486 12842 8554 12898
rect 8610 12842 8620 12898
rect 7552 12832 8620 12842
rect 10669 15750 12481 15760
rect 10669 15694 10679 15750
rect 10735 15694 10803 15750
rect 10859 15694 10927 15750
rect 10983 15694 11051 15750
rect 11107 15694 11175 15750
rect 11231 15694 11299 15750
rect 11355 15694 11423 15750
rect 11479 15694 11547 15750
rect 11603 15694 11671 15750
rect 11727 15694 11795 15750
rect 11851 15694 11919 15750
rect 11975 15694 12043 15750
rect 12099 15694 12167 15750
rect 12223 15694 12291 15750
rect 12347 15694 12415 15750
rect 12471 15694 12481 15750
rect 10669 15626 12481 15694
rect 10669 15570 10679 15626
rect 10735 15570 10803 15626
rect 10859 15570 10927 15626
rect 10983 15570 11051 15626
rect 11107 15570 11175 15626
rect 11231 15570 11299 15626
rect 11355 15570 11423 15626
rect 11479 15570 11547 15626
rect 11603 15570 11671 15626
rect 11727 15570 11795 15626
rect 11851 15570 11919 15626
rect 11975 15570 12043 15626
rect 12099 15570 12167 15626
rect 12223 15570 12291 15626
rect 12347 15570 12415 15626
rect 12471 15570 12481 15626
rect 10669 15502 12481 15570
rect 10669 15446 10679 15502
rect 10735 15446 10803 15502
rect 10859 15446 10927 15502
rect 10983 15446 11051 15502
rect 11107 15446 11175 15502
rect 11231 15446 11299 15502
rect 11355 15446 11423 15502
rect 11479 15446 11547 15502
rect 11603 15446 11671 15502
rect 11727 15446 11795 15502
rect 11851 15446 11919 15502
rect 11975 15446 12043 15502
rect 12099 15446 12167 15502
rect 12223 15446 12291 15502
rect 12347 15446 12415 15502
rect 12471 15446 12481 15502
rect 10669 15378 12481 15446
rect 10669 15322 10679 15378
rect 10735 15322 10803 15378
rect 10859 15322 10927 15378
rect 10983 15322 11051 15378
rect 11107 15322 11175 15378
rect 11231 15322 11299 15378
rect 11355 15322 11423 15378
rect 11479 15322 11547 15378
rect 11603 15322 11671 15378
rect 11727 15322 11795 15378
rect 11851 15322 11919 15378
rect 11975 15322 12043 15378
rect 12099 15322 12167 15378
rect 12223 15322 12291 15378
rect 12347 15322 12415 15378
rect 12471 15322 12481 15378
rect 10669 15254 12481 15322
rect 10669 15198 10679 15254
rect 10735 15198 10803 15254
rect 10859 15198 10927 15254
rect 10983 15198 11051 15254
rect 11107 15198 11175 15254
rect 11231 15198 11299 15254
rect 11355 15198 11423 15254
rect 11479 15198 11547 15254
rect 11603 15198 11671 15254
rect 11727 15198 11795 15254
rect 11851 15198 11919 15254
rect 11975 15198 12043 15254
rect 12099 15198 12167 15254
rect 12223 15198 12291 15254
rect 12347 15198 12415 15254
rect 12471 15198 12481 15254
rect 10669 15130 12481 15198
rect 10669 15074 10679 15130
rect 10735 15074 10803 15130
rect 10859 15074 10927 15130
rect 10983 15074 11051 15130
rect 11107 15074 11175 15130
rect 11231 15074 11299 15130
rect 11355 15074 11423 15130
rect 11479 15074 11547 15130
rect 11603 15074 11671 15130
rect 11727 15074 11795 15130
rect 11851 15074 11919 15130
rect 11975 15074 12043 15130
rect 12099 15074 12167 15130
rect 12223 15074 12291 15130
rect 12347 15074 12415 15130
rect 12471 15074 12481 15130
rect 10669 15006 12481 15074
rect 10669 14950 10679 15006
rect 10735 14950 10803 15006
rect 10859 14950 10927 15006
rect 10983 14950 11051 15006
rect 11107 14950 11175 15006
rect 11231 14950 11299 15006
rect 11355 14950 11423 15006
rect 11479 14950 11547 15006
rect 11603 14950 11671 15006
rect 11727 14950 11795 15006
rect 11851 14950 11919 15006
rect 11975 14950 12043 15006
rect 12099 14950 12167 15006
rect 12223 14950 12291 15006
rect 12347 14950 12415 15006
rect 12471 14950 12481 15006
rect 10669 14882 12481 14950
rect 10669 14826 10679 14882
rect 10735 14826 10803 14882
rect 10859 14826 10927 14882
rect 10983 14826 11051 14882
rect 11107 14826 11175 14882
rect 11231 14826 11299 14882
rect 11355 14826 11423 14882
rect 11479 14826 11547 14882
rect 11603 14826 11671 14882
rect 11727 14826 11795 14882
rect 11851 14826 11919 14882
rect 11975 14826 12043 14882
rect 12099 14826 12167 14882
rect 12223 14826 12291 14882
rect 12347 14826 12415 14882
rect 12471 14826 12481 14882
rect 10669 14758 12481 14826
rect 10669 14702 10679 14758
rect 10735 14702 10803 14758
rect 10859 14702 10927 14758
rect 10983 14702 11051 14758
rect 11107 14702 11175 14758
rect 11231 14702 11299 14758
rect 11355 14702 11423 14758
rect 11479 14702 11547 14758
rect 11603 14702 11671 14758
rect 11727 14702 11795 14758
rect 11851 14702 11919 14758
rect 11975 14702 12043 14758
rect 12099 14702 12167 14758
rect 12223 14702 12291 14758
rect 12347 14702 12415 14758
rect 12471 14702 12481 14758
rect 10669 14634 12481 14702
rect 10669 14578 10679 14634
rect 10735 14578 10803 14634
rect 10859 14578 10927 14634
rect 10983 14578 11051 14634
rect 11107 14578 11175 14634
rect 11231 14578 11299 14634
rect 11355 14578 11423 14634
rect 11479 14578 11547 14634
rect 11603 14578 11671 14634
rect 11727 14578 11795 14634
rect 11851 14578 11919 14634
rect 11975 14578 12043 14634
rect 12099 14578 12167 14634
rect 12223 14578 12291 14634
rect 12347 14578 12415 14634
rect 12471 14578 12481 14634
rect 10669 14510 12481 14578
rect 10669 14454 10679 14510
rect 10735 14454 10803 14510
rect 10859 14454 10927 14510
rect 10983 14454 11051 14510
rect 11107 14454 11175 14510
rect 11231 14454 11299 14510
rect 11355 14454 11423 14510
rect 11479 14454 11547 14510
rect 11603 14454 11671 14510
rect 11727 14454 11795 14510
rect 11851 14454 11919 14510
rect 11975 14454 12043 14510
rect 12099 14454 12167 14510
rect 12223 14454 12291 14510
rect 12347 14454 12415 14510
rect 12471 14454 12481 14510
rect 10669 14386 12481 14454
rect 10669 14330 10679 14386
rect 10735 14330 10803 14386
rect 10859 14330 10927 14386
rect 10983 14330 11051 14386
rect 11107 14330 11175 14386
rect 11231 14330 11299 14386
rect 11355 14330 11423 14386
rect 11479 14330 11547 14386
rect 11603 14330 11671 14386
rect 11727 14330 11795 14386
rect 11851 14330 11919 14386
rect 11975 14330 12043 14386
rect 12099 14330 12167 14386
rect 12223 14330 12291 14386
rect 12347 14330 12415 14386
rect 12471 14330 12481 14386
rect 10669 14262 12481 14330
rect 10669 14206 10679 14262
rect 10735 14206 10803 14262
rect 10859 14206 10927 14262
rect 10983 14206 11051 14262
rect 11107 14206 11175 14262
rect 11231 14206 11299 14262
rect 11355 14206 11423 14262
rect 11479 14206 11547 14262
rect 11603 14206 11671 14262
rect 11727 14206 11795 14262
rect 11851 14206 11919 14262
rect 11975 14206 12043 14262
rect 12099 14206 12167 14262
rect 12223 14206 12291 14262
rect 12347 14206 12415 14262
rect 12471 14206 12481 14262
rect 10669 14138 12481 14206
rect 10669 14082 10679 14138
rect 10735 14082 10803 14138
rect 10859 14082 10927 14138
rect 10983 14082 11051 14138
rect 11107 14082 11175 14138
rect 11231 14082 11299 14138
rect 11355 14082 11423 14138
rect 11479 14082 11547 14138
rect 11603 14082 11671 14138
rect 11727 14082 11795 14138
rect 11851 14082 11919 14138
rect 11975 14082 12043 14138
rect 12099 14082 12167 14138
rect 12223 14082 12291 14138
rect 12347 14082 12415 14138
rect 12471 14082 12481 14138
rect 10669 14014 12481 14082
rect 10669 13958 10679 14014
rect 10735 13958 10803 14014
rect 10859 13958 10927 14014
rect 10983 13958 11051 14014
rect 11107 13958 11175 14014
rect 11231 13958 11299 14014
rect 11355 13958 11423 14014
rect 11479 13958 11547 14014
rect 11603 13958 11671 14014
rect 11727 13958 11795 14014
rect 11851 13958 11919 14014
rect 11975 13958 12043 14014
rect 12099 13958 12167 14014
rect 12223 13958 12291 14014
rect 12347 13958 12415 14014
rect 12471 13958 12481 14014
rect 10669 13890 12481 13958
rect 10669 13834 10679 13890
rect 10735 13834 10803 13890
rect 10859 13834 10927 13890
rect 10983 13834 11051 13890
rect 11107 13834 11175 13890
rect 11231 13834 11299 13890
rect 11355 13834 11423 13890
rect 11479 13834 11547 13890
rect 11603 13834 11671 13890
rect 11727 13834 11795 13890
rect 11851 13834 11919 13890
rect 11975 13834 12043 13890
rect 12099 13834 12167 13890
rect 12223 13834 12291 13890
rect 12347 13834 12415 13890
rect 12471 13834 12481 13890
rect 10669 13766 12481 13834
rect 10669 13710 10679 13766
rect 10735 13710 10803 13766
rect 10859 13710 10927 13766
rect 10983 13710 11051 13766
rect 11107 13710 11175 13766
rect 11231 13710 11299 13766
rect 11355 13710 11423 13766
rect 11479 13710 11547 13766
rect 11603 13710 11671 13766
rect 11727 13710 11795 13766
rect 11851 13710 11919 13766
rect 11975 13710 12043 13766
rect 12099 13710 12167 13766
rect 12223 13710 12291 13766
rect 12347 13710 12415 13766
rect 12471 13710 12481 13766
rect 10669 13642 12481 13710
rect 10669 13586 10679 13642
rect 10735 13586 10803 13642
rect 10859 13586 10927 13642
rect 10983 13586 11051 13642
rect 11107 13586 11175 13642
rect 11231 13586 11299 13642
rect 11355 13586 11423 13642
rect 11479 13586 11547 13642
rect 11603 13586 11671 13642
rect 11727 13586 11795 13642
rect 11851 13586 11919 13642
rect 11975 13586 12043 13642
rect 12099 13586 12167 13642
rect 12223 13586 12291 13642
rect 12347 13586 12415 13642
rect 12471 13586 12481 13642
rect 10669 13518 12481 13586
rect 10669 13462 10679 13518
rect 10735 13462 10803 13518
rect 10859 13462 10927 13518
rect 10983 13462 11051 13518
rect 11107 13462 11175 13518
rect 11231 13462 11299 13518
rect 11355 13462 11423 13518
rect 11479 13462 11547 13518
rect 11603 13462 11671 13518
rect 11727 13462 11795 13518
rect 11851 13462 11919 13518
rect 11975 13462 12043 13518
rect 12099 13462 12167 13518
rect 12223 13462 12291 13518
rect 12347 13462 12415 13518
rect 12471 13462 12481 13518
rect 10669 13394 12481 13462
rect 10669 13338 10679 13394
rect 10735 13338 10803 13394
rect 10859 13338 10927 13394
rect 10983 13338 11051 13394
rect 11107 13338 11175 13394
rect 11231 13338 11299 13394
rect 11355 13338 11423 13394
rect 11479 13338 11547 13394
rect 11603 13338 11671 13394
rect 11727 13338 11795 13394
rect 11851 13338 11919 13394
rect 11975 13338 12043 13394
rect 12099 13338 12167 13394
rect 12223 13338 12291 13394
rect 12347 13338 12415 13394
rect 12471 13338 12481 13394
rect 10669 13270 12481 13338
rect 10669 13214 10679 13270
rect 10735 13214 10803 13270
rect 10859 13214 10927 13270
rect 10983 13214 11051 13270
rect 11107 13214 11175 13270
rect 11231 13214 11299 13270
rect 11355 13214 11423 13270
rect 11479 13214 11547 13270
rect 11603 13214 11671 13270
rect 11727 13214 11795 13270
rect 11851 13214 11919 13270
rect 11975 13214 12043 13270
rect 12099 13214 12167 13270
rect 12223 13214 12291 13270
rect 12347 13214 12415 13270
rect 12471 13214 12481 13270
rect 10669 13146 12481 13214
rect 10669 13090 10679 13146
rect 10735 13090 10803 13146
rect 10859 13090 10927 13146
rect 10983 13090 11051 13146
rect 11107 13090 11175 13146
rect 11231 13090 11299 13146
rect 11355 13090 11423 13146
rect 11479 13090 11547 13146
rect 11603 13090 11671 13146
rect 11727 13090 11795 13146
rect 11851 13090 11919 13146
rect 11975 13090 12043 13146
rect 12099 13090 12167 13146
rect 12223 13090 12291 13146
rect 12347 13090 12415 13146
rect 12471 13090 12481 13146
rect 10669 13022 12481 13090
rect 10669 12966 10679 13022
rect 10735 12966 10803 13022
rect 10859 12966 10927 13022
rect 10983 12966 11051 13022
rect 11107 12966 11175 13022
rect 11231 12966 11299 13022
rect 11355 12966 11423 13022
rect 11479 12966 11547 13022
rect 11603 12966 11671 13022
rect 11727 12966 11795 13022
rect 11851 12966 11919 13022
rect 11975 12966 12043 13022
rect 12099 12966 12167 13022
rect 12223 12966 12291 13022
rect 12347 12966 12415 13022
rect 12471 12966 12481 13022
rect 10669 12898 12481 12966
rect 10669 12842 10679 12898
rect 10735 12842 10803 12898
rect 10859 12842 10927 12898
rect 10983 12842 11051 12898
rect 11107 12842 11175 12898
rect 11231 12842 11299 12898
rect 11355 12842 11423 12898
rect 11479 12842 11547 12898
rect 11603 12842 11671 12898
rect 11727 12842 11795 12898
rect 11851 12842 11919 12898
rect 11975 12842 12043 12898
rect 12099 12842 12167 12898
rect 12223 12842 12291 12898
rect 12347 12842 12415 12898
rect 12471 12842 12481 12898
rect 10669 12832 12481 12842
rect 2497 12544 4309 12554
rect 2497 12488 2507 12544
rect 2563 12488 2631 12544
rect 2687 12488 2755 12544
rect 2811 12488 2879 12544
rect 2935 12488 3003 12544
rect 3059 12488 3127 12544
rect 3183 12488 3251 12544
rect 3307 12488 3375 12544
rect 3431 12488 3499 12544
rect 3555 12488 3623 12544
rect 3679 12488 3747 12544
rect 3803 12488 3871 12544
rect 3927 12488 3995 12544
rect 4051 12488 4119 12544
rect 4175 12488 4243 12544
rect 4299 12488 4309 12544
rect 2497 12420 4309 12488
rect 2497 12364 2507 12420
rect 2563 12364 2631 12420
rect 2687 12364 2755 12420
rect 2811 12364 2879 12420
rect 2935 12364 3003 12420
rect 3059 12364 3127 12420
rect 3183 12364 3251 12420
rect 3307 12364 3375 12420
rect 3431 12364 3499 12420
rect 3555 12364 3623 12420
rect 3679 12364 3747 12420
rect 3803 12364 3871 12420
rect 3927 12364 3995 12420
rect 4051 12364 4119 12420
rect 4175 12364 4243 12420
rect 4299 12364 4309 12420
rect 2497 12296 4309 12364
rect 2497 12240 2507 12296
rect 2563 12240 2631 12296
rect 2687 12240 2755 12296
rect 2811 12240 2879 12296
rect 2935 12240 3003 12296
rect 3059 12240 3127 12296
rect 3183 12240 3251 12296
rect 3307 12240 3375 12296
rect 3431 12240 3499 12296
rect 3555 12240 3623 12296
rect 3679 12240 3747 12296
rect 3803 12240 3871 12296
rect 3927 12240 3995 12296
rect 4051 12240 4119 12296
rect 4175 12240 4243 12296
rect 4299 12240 4309 12296
rect 2497 12172 4309 12240
rect 2497 12116 2507 12172
rect 2563 12116 2631 12172
rect 2687 12116 2755 12172
rect 2811 12116 2879 12172
rect 2935 12116 3003 12172
rect 3059 12116 3127 12172
rect 3183 12116 3251 12172
rect 3307 12116 3375 12172
rect 3431 12116 3499 12172
rect 3555 12116 3623 12172
rect 3679 12116 3747 12172
rect 3803 12116 3871 12172
rect 3927 12116 3995 12172
rect 4051 12116 4119 12172
rect 4175 12116 4243 12172
rect 4299 12116 4309 12172
rect 2497 12048 4309 12116
rect 2497 11992 2507 12048
rect 2563 11992 2631 12048
rect 2687 11992 2755 12048
rect 2811 11992 2879 12048
rect 2935 11992 3003 12048
rect 3059 11992 3127 12048
rect 3183 11992 3251 12048
rect 3307 11992 3375 12048
rect 3431 11992 3499 12048
rect 3555 11992 3623 12048
rect 3679 11992 3747 12048
rect 3803 11992 3871 12048
rect 3927 11992 3995 12048
rect 4051 11992 4119 12048
rect 4175 11992 4243 12048
rect 4299 11992 4309 12048
rect 2497 11924 4309 11992
rect 2497 11868 2507 11924
rect 2563 11868 2631 11924
rect 2687 11868 2755 11924
rect 2811 11868 2879 11924
rect 2935 11868 3003 11924
rect 3059 11868 3127 11924
rect 3183 11868 3251 11924
rect 3307 11868 3375 11924
rect 3431 11868 3499 11924
rect 3555 11868 3623 11924
rect 3679 11868 3747 11924
rect 3803 11868 3871 11924
rect 3927 11868 3995 11924
rect 4051 11868 4119 11924
rect 4175 11868 4243 11924
rect 4299 11868 4309 11924
rect 2497 11800 4309 11868
rect 2497 11744 2507 11800
rect 2563 11744 2631 11800
rect 2687 11744 2755 11800
rect 2811 11744 2879 11800
rect 2935 11744 3003 11800
rect 3059 11744 3127 11800
rect 3183 11744 3251 11800
rect 3307 11744 3375 11800
rect 3431 11744 3499 11800
rect 3555 11744 3623 11800
rect 3679 11744 3747 11800
rect 3803 11744 3871 11800
rect 3927 11744 3995 11800
rect 4051 11744 4119 11800
rect 4175 11744 4243 11800
rect 4299 11744 4309 11800
rect 2497 11676 4309 11744
rect 2497 11620 2507 11676
rect 2563 11620 2631 11676
rect 2687 11620 2755 11676
rect 2811 11620 2879 11676
rect 2935 11620 3003 11676
rect 3059 11620 3127 11676
rect 3183 11620 3251 11676
rect 3307 11620 3375 11676
rect 3431 11620 3499 11676
rect 3555 11620 3623 11676
rect 3679 11620 3747 11676
rect 3803 11620 3871 11676
rect 3927 11620 3995 11676
rect 4051 11620 4119 11676
rect 4175 11620 4243 11676
rect 4299 11620 4309 11676
rect 2497 11552 4309 11620
rect 2497 11496 2507 11552
rect 2563 11496 2631 11552
rect 2687 11496 2755 11552
rect 2811 11496 2879 11552
rect 2935 11496 3003 11552
rect 3059 11496 3127 11552
rect 3183 11496 3251 11552
rect 3307 11496 3375 11552
rect 3431 11496 3499 11552
rect 3555 11496 3623 11552
rect 3679 11496 3747 11552
rect 3803 11496 3871 11552
rect 3927 11496 3995 11552
rect 4051 11496 4119 11552
rect 4175 11496 4243 11552
rect 4299 11496 4309 11552
rect 2497 11428 4309 11496
rect 2497 11372 2507 11428
rect 2563 11372 2631 11428
rect 2687 11372 2755 11428
rect 2811 11372 2879 11428
rect 2935 11372 3003 11428
rect 3059 11372 3127 11428
rect 3183 11372 3251 11428
rect 3307 11372 3375 11428
rect 3431 11372 3499 11428
rect 3555 11372 3623 11428
rect 3679 11372 3747 11428
rect 3803 11372 3871 11428
rect 3927 11372 3995 11428
rect 4051 11372 4119 11428
rect 4175 11372 4243 11428
rect 4299 11372 4309 11428
rect 2497 11304 4309 11372
rect 2497 11248 2507 11304
rect 2563 11248 2631 11304
rect 2687 11248 2755 11304
rect 2811 11248 2879 11304
rect 2935 11248 3003 11304
rect 3059 11248 3127 11304
rect 3183 11248 3251 11304
rect 3307 11248 3375 11304
rect 3431 11248 3499 11304
rect 3555 11248 3623 11304
rect 3679 11248 3747 11304
rect 3803 11248 3871 11304
rect 3927 11248 3995 11304
rect 4051 11248 4119 11304
rect 4175 11248 4243 11304
rect 4299 11248 4309 11304
rect 2497 11238 4309 11248
rect 6358 12544 7426 12554
rect 6358 12488 6368 12544
rect 6424 12488 6492 12544
rect 6548 12488 6616 12544
rect 6672 12488 6740 12544
rect 6796 12488 6864 12544
rect 6920 12488 6988 12544
rect 7044 12488 7112 12544
rect 7168 12488 7236 12544
rect 7292 12488 7360 12544
rect 7416 12488 7426 12544
rect 6358 12420 7426 12488
rect 6358 12364 6368 12420
rect 6424 12364 6492 12420
rect 6548 12364 6616 12420
rect 6672 12364 6740 12420
rect 6796 12364 6864 12420
rect 6920 12364 6988 12420
rect 7044 12364 7112 12420
rect 7168 12364 7236 12420
rect 7292 12364 7360 12420
rect 7416 12364 7426 12420
rect 6358 12296 7426 12364
rect 6358 12240 6368 12296
rect 6424 12240 6492 12296
rect 6548 12240 6616 12296
rect 6672 12240 6740 12296
rect 6796 12240 6864 12296
rect 6920 12240 6988 12296
rect 7044 12240 7112 12296
rect 7168 12240 7236 12296
rect 7292 12240 7360 12296
rect 7416 12240 7426 12296
rect 6358 12172 7426 12240
rect 6358 12116 6368 12172
rect 6424 12116 6492 12172
rect 6548 12116 6616 12172
rect 6672 12116 6740 12172
rect 6796 12116 6864 12172
rect 6920 12116 6988 12172
rect 7044 12116 7112 12172
rect 7168 12116 7236 12172
rect 7292 12116 7360 12172
rect 7416 12116 7426 12172
rect 6358 12048 7426 12116
rect 6358 11992 6368 12048
rect 6424 11992 6492 12048
rect 6548 11992 6616 12048
rect 6672 11992 6740 12048
rect 6796 11992 6864 12048
rect 6920 11992 6988 12048
rect 7044 11992 7112 12048
rect 7168 11992 7236 12048
rect 7292 11992 7360 12048
rect 7416 11992 7426 12048
rect 6358 11924 7426 11992
rect 6358 11868 6368 11924
rect 6424 11868 6492 11924
rect 6548 11868 6616 11924
rect 6672 11868 6740 11924
rect 6796 11868 6864 11924
rect 6920 11868 6988 11924
rect 7044 11868 7112 11924
rect 7168 11868 7236 11924
rect 7292 11868 7360 11924
rect 7416 11868 7426 11924
rect 6358 11800 7426 11868
rect 6358 11744 6368 11800
rect 6424 11744 6492 11800
rect 6548 11744 6616 11800
rect 6672 11744 6740 11800
rect 6796 11744 6864 11800
rect 6920 11744 6988 11800
rect 7044 11744 7112 11800
rect 7168 11744 7236 11800
rect 7292 11744 7360 11800
rect 7416 11744 7426 11800
rect 6358 11676 7426 11744
rect 6358 11620 6368 11676
rect 6424 11620 6492 11676
rect 6548 11620 6616 11676
rect 6672 11620 6740 11676
rect 6796 11620 6864 11676
rect 6920 11620 6988 11676
rect 7044 11620 7112 11676
rect 7168 11620 7236 11676
rect 7292 11620 7360 11676
rect 7416 11620 7426 11676
rect 6358 11552 7426 11620
rect 6358 11496 6368 11552
rect 6424 11496 6492 11552
rect 6548 11496 6616 11552
rect 6672 11496 6740 11552
rect 6796 11496 6864 11552
rect 6920 11496 6988 11552
rect 7044 11496 7112 11552
rect 7168 11496 7236 11552
rect 7292 11496 7360 11552
rect 7416 11496 7426 11552
rect 6358 11428 7426 11496
rect 6358 11372 6368 11428
rect 6424 11372 6492 11428
rect 6548 11372 6616 11428
rect 6672 11372 6740 11428
rect 6796 11372 6864 11428
rect 6920 11372 6988 11428
rect 7044 11372 7112 11428
rect 7168 11372 7236 11428
rect 7292 11372 7360 11428
rect 7416 11372 7426 11428
rect 6358 11304 7426 11372
rect 6358 11248 6368 11304
rect 6424 11248 6492 11304
rect 6548 11248 6616 11304
rect 6672 11248 6740 11304
rect 6796 11248 6864 11304
rect 6920 11248 6988 11304
rect 7044 11248 7112 11304
rect 7168 11248 7236 11304
rect 7292 11248 7360 11304
rect 7416 11248 7426 11304
rect 6358 11238 7426 11248
rect 8741 12544 10553 12554
rect 8741 12488 8751 12544
rect 8807 12488 8875 12544
rect 8931 12488 8999 12544
rect 9055 12488 9123 12544
rect 9179 12488 9247 12544
rect 9303 12488 9371 12544
rect 9427 12488 9495 12544
rect 9551 12488 9619 12544
rect 9675 12488 9743 12544
rect 9799 12488 9867 12544
rect 9923 12488 9991 12544
rect 10047 12488 10115 12544
rect 10171 12488 10239 12544
rect 10295 12488 10363 12544
rect 10419 12488 10487 12544
rect 10543 12488 10553 12544
rect 8741 12420 10553 12488
rect 8741 12364 8751 12420
rect 8807 12364 8875 12420
rect 8931 12364 8999 12420
rect 9055 12364 9123 12420
rect 9179 12364 9247 12420
rect 9303 12364 9371 12420
rect 9427 12364 9495 12420
rect 9551 12364 9619 12420
rect 9675 12364 9743 12420
rect 9799 12364 9867 12420
rect 9923 12364 9991 12420
rect 10047 12364 10115 12420
rect 10171 12364 10239 12420
rect 10295 12364 10363 12420
rect 10419 12364 10487 12420
rect 10543 12364 10553 12420
rect 8741 12296 10553 12364
rect 8741 12240 8751 12296
rect 8807 12240 8875 12296
rect 8931 12240 8999 12296
rect 9055 12240 9123 12296
rect 9179 12240 9247 12296
rect 9303 12240 9371 12296
rect 9427 12240 9495 12296
rect 9551 12240 9619 12296
rect 9675 12240 9743 12296
rect 9799 12240 9867 12296
rect 9923 12240 9991 12296
rect 10047 12240 10115 12296
rect 10171 12240 10239 12296
rect 10295 12240 10363 12296
rect 10419 12240 10487 12296
rect 10543 12240 10553 12296
rect 8741 12172 10553 12240
rect 8741 12116 8751 12172
rect 8807 12116 8875 12172
rect 8931 12116 8999 12172
rect 9055 12116 9123 12172
rect 9179 12116 9247 12172
rect 9303 12116 9371 12172
rect 9427 12116 9495 12172
rect 9551 12116 9619 12172
rect 9675 12116 9743 12172
rect 9799 12116 9867 12172
rect 9923 12116 9991 12172
rect 10047 12116 10115 12172
rect 10171 12116 10239 12172
rect 10295 12116 10363 12172
rect 10419 12116 10487 12172
rect 10543 12116 10553 12172
rect 8741 12048 10553 12116
rect 8741 11992 8751 12048
rect 8807 11992 8875 12048
rect 8931 11992 8999 12048
rect 9055 11992 9123 12048
rect 9179 11992 9247 12048
rect 9303 11992 9371 12048
rect 9427 11992 9495 12048
rect 9551 11992 9619 12048
rect 9675 11992 9743 12048
rect 9799 11992 9867 12048
rect 9923 11992 9991 12048
rect 10047 11992 10115 12048
rect 10171 11992 10239 12048
rect 10295 11992 10363 12048
rect 10419 11992 10487 12048
rect 10543 11992 10553 12048
rect 8741 11924 10553 11992
rect 8741 11868 8751 11924
rect 8807 11868 8875 11924
rect 8931 11868 8999 11924
rect 9055 11868 9123 11924
rect 9179 11868 9247 11924
rect 9303 11868 9371 11924
rect 9427 11868 9495 11924
rect 9551 11868 9619 11924
rect 9675 11868 9743 11924
rect 9799 11868 9867 11924
rect 9923 11868 9991 11924
rect 10047 11868 10115 11924
rect 10171 11868 10239 11924
rect 10295 11868 10363 11924
rect 10419 11868 10487 11924
rect 10543 11868 10553 11924
rect 8741 11800 10553 11868
rect 8741 11744 8751 11800
rect 8807 11744 8875 11800
rect 8931 11744 8999 11800
rect 9055 11744 9123 11800
rect 9179 11744 9247 11800
rect 9303 11744 9371 11800
rect 9427 11744 9495 11800
rect 9551 11744 9619 11800
rect 9675 11744 9743 11800
rect 9799 11744 9867 11800
rect 9923 11744 9991 11800
rect 10047 11744 10115 11800
rect 10171 11744 10239 11800
rect 10295 11744 10363 11800
rect 10419 11744 10487 11800
rect 10543 11744 10553 11800
rect 8741 11676 10553 11744
rect 8741 11620 8751 11676
rect 8807 11620 8875 11676
rect 8931 11620 8999 11676
rect 9055 11620 9123 11676
rect 9179 11620 9247 11676
rect 9303 11620 9371 11676
rect 9427 11620 9495 11676
rect 9551 11620 9619 11676
rect 9675 11620 9743 11676
rect 9799 11620 9867 11676
rect 9923 11620 9991 11676
rect 10047 11620 10115 11676
rect 10171 11620 10239 11676
rect 10295 11620 10363 11676
rect 10419 11620 10487 11676
rect 10543 11620 10553 11676
rect 8741 11552 10553 11620
rect 8741 11496 8751 11552
rect 8807 11496 8875 11552
rect 8931 11496 8999 11552
rect 9055 11496 9123 11552
rect 9179 11496 9247 11552
rect 9303 11496 9371 11552
rect 9427 11496 9495 11552
rect 9551 11496 9619 11552
rect 9675 11496 9743 11552
rect 9799 11496 9867 11552
rect 9923 11496 9991 11552
rect 10047 11496 10115 11552
rect 10171 11496 10239 11552
rect 10295 11496 10363 11552
rect 10419 11496 10487 11552
rect 10543 11496 10553 11552
rect 8741 11428 10553 11496
rect 8741 11372 8751 11428
rect 8807 11372 8875 11428
rect 8931 11372 8999 11428
rect 9055 11372 9123 11428
rect 9179 11372 9247 11428
rect 9303 11372 9371 11428
rect 9427 11372 9495 11428
rect 9551 11372 9619 11428
rect 9675 11372 9743 11428
rect 9799 11372 9867 11428
rect 9923 11372 9991 11428
rect 10047 11372 10115 11428
rect 10171 11372 10239 11428
rect 10295 11372 10363 11428
rect 10419 11372 10487 11428
rect 10543 11372 10553 11428
rect 8741 11304 10553 11372
rect 8741 11248 8751 11304
rect 8807 11248 8875 11304
rect 8931 11248 8999 11304
rect 9055 11248 9123 11304
rect 9179 11248 9247 11304
rect 9303 11248 9371 11304
rect 9427 11248 9495 11304
rect 9551 11248 9619 11304
rect 9675 11248 9743 11304
rect 9799 11248 9867 11304
rect 9923 11248 9991 11304
rect 10047 11248 10115 11304
rect 10171 11248 10239 11304
rect 10295 11248 10363 11304
rect 10419 11248 10487 11304
rect 10543 11248 10553 11304
rect 8741 11238 10553 11248
rect 12842 12544 13910 12554
rect 12842 12488 12852 12544
rect 12908 12488 12976 12544
rect 13032 12488 13100 12544
rect 13156 12488 13224 12544
rect 13280 12488 13348 12544
rect 13404 12488 13472 12544
rect 13528 12488 13596 12544
rect 13652 12488 13720 12544
rect 13776 12488 13844 12544
rect 13900 12488 13910 12544
rect 12842 12420 13910 12488
rect 12842 12364 12852 12420
rect 12908 12364 12976 12420
rect 13032 12364 13100 12420
rect 13156 12364 13224 12420
rect 13280 12364 13348 12420
rect 13404 12364 13472 12420
rect 13528 12364 13596 12420
rect 13652 12364 13720 12420
rect 13776 12364 13844 12420
rect 13900 12364 13910 12420
rect 12842 12296 13910 12364
rect 12842 12240 12852 12296
rect 12908 12240 12976 12296
rect 13032 12240 13100 12296
rect 13156 12240 13224 12296
rect 13280 12240 13348 12296
rect 13404 12240 13472 12296
rect 13528 12240 13596 12296
rect 13652 12240 13720 12296
rect 13776 12240 13844 12296
rect 13900 12240 13910 12296
rect 12842 12172 13910 12240
rect 12842 12116 12852 12172
rect 12908 12116 12976 12172
rect 13032 12116 13100 12172
rect 13156 12116 13224 12172
rect 13280 12116 13348 12172
rect 13404 12116 13472 12172
rect 13528 12116 13596 12172
rect 13652 12116 13720 12172
rect 13776 12116 13844 12172
rect 13900 12116 13910 12172
rect 12842 12048 13910 12116
rect 12842 11992 12852 12048
rect 12908 11992 12976 12048
rect 13032 11992 13100 12048
rect 13156 11992 13224 12048
rect 13280 11992 13348 12048
rect 13404 11992 13472 12048
rect 13528 11992 13596 12048
rect 13652 11992 13720 12048
rect 13776 11992 13844 12048
rect 13900 11992 13910 12048
rect 12842 11924 13910 11992
rect 12842 11868 12852 11924
rect 12908 11868 12976 11924
rect 13032 11868 13100 11924
rect 13156 11868 13224 11924
rect 13280 11868 13348 11924
rect 13404 11868 13472 11924
rect 13528 11868 13596 11924
rect 13652 11868 13720 11924
rect 13776 11868 13844 11924
rect 13900 11868 13910 11924
rect 12842 11800 13910 11868
rect 12842 11744 12852 11800
rect 12908 11744 12976 11800
rect 13032 11744 13100 11800
rect 13156 11744 13224 11800
rect 13280 11744 13348 11800
rect 13404 11744 13472 11800
rect 13528 11744 13596 11800
rect 13652 11744 13720 11800
rect 13776 11744 13844 11800
rect 13900 11744 13910 11800
rect 12842 11676 13910 11744
rect 12842 11620 12852 11676
rect 12908 11620 12976 11676
rect 13032 11620 13100 11676
rect 13156 11620 13224 11676
rect 13280 11620 13348 11676
rect 13404 11620 13472 11676
rect 13528 11620 13596 11676
rect 13652 11620 13720 11676
rect 13776 11620 13844 11676
rect 13900 11620 13910 11676
rect 12842 11552 13910 11620
rect 12842 11496 12852 11552
rect 12908 11496 12976 11552
rect 13032 11496 13100 11552
rect 13156 11496 13224 11552
rect 13280 11496 13348 11552
rect 13404 11496 13472 11552
rect 13528 11496 13596 11552
rect 13652 11496 13720 11552
rect 13776 11496 13844 11552
rect 13900 11496 13910 11552
rect 12842 11428 13910 11496
rect 12842 11372 12852 11428
rect 12908 11372 12976 11428
rect 13032 11372 13100 11428
rect 13156 11372 13224 11428
rect 13280 11372 13348 11428
rect 13404 11372 13472 11428
rect 13528 11372 13596 11428
rect 13652 11372 13720 11428
rect 13776 11372 13844 11428
rect 13900 11372 13910 11428
rect 12842 11304 13910 11372
rect 12842 11248 12852 11304
rect 12908 11248 12976 11304
rect 13032 11248 13100 11304
rect 13156 11248 13224 11304
rect 13280 11248 13348 11304
rect 13404 11248 13472 11304
rect 13528 11248 13596 11304
rect 13652 11248 13720 11304
rect 13776 11248 13844 11304
rect 13900 11248 13910 11304
rect 12842 11238 13910 11248
rect 1068 10944 2136 10954
rect 1068 10888 1078 10944
rect 1134 10888 1202 10944
rect 1258 10888 1326 10944
rect 1382 10888 1450 10944
rect 1506 10888 1574 10944
rect 1630 10888 1698 10944
rect 1754 10888 1822 10944
rect 1878 10888 1946 10944
rect 2002 10888 2070 10944
rect 2126 10888 2136 10944
rect 1068 10820 2136 10888
rect 1068 10764 1078 10820
rect 1134 10764 1202 10820
rect 1258 10764 1326 10820
rect 1382 10764 1450 10820
rect 1506 10764 1574 10820
rect 1630 10764 1698 10820
rect 1754 10764 1822 10820
rect 1878 10764 1946 10820
rect 2002 10764 2070 10820
rect 2126 10764 2136 10820
rect 1068 10696 2136 10764
rect 1068 10640 1078 10696
rect 1134 10640 1202 10696
rect 1258 10640 1326 10696
rect 1382 10640 1450 10696
rect 1506 10640 1574 10696
rect 1630 10640 1698 10696
rect 1754 10640 1822 10696
rect 1878 10640 1946 10696
rect 2002 10640 2070 10696
rect 2126 10640 2136 10696
rect 1068 10572 2136 10640
rect 1068 10516 1078 10572
rect 1134 10516 1202 10572
rect 1258 10516 1326 10572
rect 1382 10516 1450 10572
rect 1506 10516 1574 10572
rect 1630 10516 1698 10572
rect 1754 10516 1822 10572
rect 1878 10516 1946 10572
rect 2002 10516 2070 10572
rect 2126 10516 2136 10572
rect 1068 10448 2136 10516
rect 1068 10392 1078 10448
rect 1134 10392 1202 10448
rect 1258 10392 1326 10448
rect 1382 10392 1450 10448
rect 1506 10392 1574 10448
rect 1630 10392 1698 10448
rect 1754 10392 1822 10448
rect 1878 10392 1946 10448
rect 2002 10392 2070 10448
rect 2126 10392 2136 10448
rect 1068 10324 2136 10392
rect 1068 10268 1078 10324
rect 1134 10268 1202 10324
rect 1258 10268 1326 10324
rect 1382 10268 1450 10324
rect 1506 10268 1574 10324
rect 1630 10268 1698 10324
rect 1754 10268 1822 10324
rect 1878 10268 1946 10324
rect 2002 10268 2070 10324
rect 2126 10268 2136 10324
rect 1068 10200 2136 10268
rect 1068 10144 1078 10200
rect 1134 10144 1202 10200
rect 1258 10144 1326 10200
rect 1382 10144 1450 10200
rect 1506 10144 1574 10200
rect 1630 10144 1698 10200
rect 1754 10144 1822 10200
rect 1878 10144 1946 10200
rect 2002 10144 2070 10200
rect 2126 10144 2136 10200
rect 1068 10076 2136 10144
rect 1068 10020 1078 10076
rect 1134 10020 1202 10076
rect 1258 10020 1326 10076
rect 1382 10020 1450 10076
rect 1506 10020 1574 10076
rect 1630 10020 1698 10076
rect 1754 10020 1822 10076
rect 1878 10020 1946 10076
rect 2002 10020 2070 10076
rect 2126 10020 2136 10076
rect 1068 9952 2136 10020
rect 1068 9896 1078 9952
rect 1134 9896 1202 9952
rect 1258 9896 1326 9952
rect 1382 9896 1450 9952
rect 1506 9896 1574 9952
rect 1630 9896 1698 9952
rect 1754 9896 1822 9952
rect 1878 9896 1946 9952
rect 2002 9896 2070 9952
rect 2126 9896 2136 9952
rect 1068 9828 2136 9896
rect 1068 9772 1078 9828
rect 1134 9772 1202 9828
rect 1258 9772 1326 9828
rect 1382 9772 1450 9828
rect 1506 9772 1574 9828
rect 1630 9772 1698 9828
rect 1754 9772 1822 9828
rect 1878 9772 1946 9828
rect 2002 9772 2070 9828
rect 2126 9772 2136 9828
rect 1068 9704 2136 9772
rect 1068 9648 1078 9704
rect 1134 9648 1202 9704
rect 1258 9648 1326 9704
rect 1382 9648 1450 9704
rect 1506 9648 1574 9704
rect 1630 9648 1698 9704
rect 1754 9648 1822 9704
rect 1878 9648 1946 9704
rect 2002 9648 2070 9704
rect 2126 9648 2136 9704
rect 1068 9638 2136 9648
rect 4425 10944 6237 10954
rect 4425 10888 4435 10944
rect 4491 10888 4559 10944
rect 4615 10888 4683 10944
rect 4739 10888 4807 10944
rect 4863 10888 4931 10944
rect 4987 10888 5055 10944
rect 5111 10888 5179 10944
rect 5235 10888 5303 10944
rect 5359 10888 5427 10944
rect 5483 10888 5551 10944
rect 5607 10888 5675 10944
rect 5731 10888 5799 10944
rect 5855 10888 5923 10944
rect 5979 10888 6047 10944
rect 6103 10888 6171 10944
rect 6227 10888 6237 10944
rect 4425 10820 6237 10888
rect 4425 10764 4435 10820
rect 4491 10764 4559 10820
rect 4615 10764 4683 10820
rect 4739 10764 4807 10820
rect 4863 10764 4931 10820
rect 4987 10764 5055 10820
rect 5111 10764 5179 10820
rect 5235 10764 5303 10820
rect 5359 10764 5427 10820
rect 5483 10764 5551 10820
rect 5607 10764 5675 10820
rect 5731 10764 5799 10820
rect 5855 10764 5923 10820
rect 5979 10764 6047 10820
rect 6103 10764 6171 10820
rect 6227 10764 6237 10820
rect 4425 10696 6237 10764
rect 4425 10640 4435 10696
rect 4491 10640 4559 10696
rect 4615 10640 4683 10696
rect 4739 10640 4807 10696
rect 4863 10640 4931 10696
rect 4987 10640 5055 10696
rect 5111 10640 5179 10696
rect 5235 10640 5303 10696
rect 5359 10640 5427 10696
rect 5483 10640 5551 10696
rect 5607 10640 5675 10696
rect 5731 10640 5799 10696
rect 5855 10640 5923 10696
rect 5979 10640 6047 10696
rect 6103 10640 6171 10696
rect 6227 10640 6237 10696
rect 4425 10572 6237 10640
rect 4425 10516 4435 10572
rect 4491 10516 4559 10572
rect 4615 10516 4683 10572
rect 4739 10516 4807 10572
rect 4863 10516 4931 10572
rect 4987 10516 5055 10572
rect 5111 10516 5179 10572
rect 5235 10516 5303 10572
rect 5359 10516 5427 10572
rect 5483 10516 5551 10572
rect 5607 10516 5675 10572
rect 5731 10516 5799 10572
rect 5855 10516 5923 10572
rect 5979 10516 6047 10572
rect 6103 10516 6171 10572
rect 6227 10516 6237 10572
rect 4425 10448 6237 10516
rect 4425 10392 4435 10448
rect 4491 10392 4559 10448
rect 4615 10392 4683 10448
rect 4739 10392 4807 10448
rect 4863 10392 4931 10448
rect 4987 10392 5055 10448
rect 5111 10392 5179 10448
rect 5235 10392 5303 10448
rect 5359 10392 5427 10448
rect 5483 10392 5551 10448
rect 5607 10392 5675 10448
rect 5731 10392 5799 10448
rect 5855 10392 5923 10448
rect 5979 10392 6047 10448
rect 6103 10392 6171 10448
rect 6227 10392 6237 10448
rect 4425 10324 6237 10392
rect 4425 10268 4435 10324
rect 4491 10268 4559 10324
rect 4615 10268 4683 10324
rect 4739 10268 4807 10324
rect 4863 10268 4931 10324
rect 4987 10268 5055 10324
rect 5111 10268 5179 10324
rect 5235 10268 5303 10324
rect 5359 10268 5427 10324
rect 5483 10268 5551 10324
rect 5607 10268 5675 10324
rect 5731 10268 5799 10324
rect 5855 10268 5923 10324
rect 5979 10268 6047 10324
rect 6103 10268 6171 10324
rect 6227 10268 6237 10324
rect 4425 10200 6237 10268
rect 4425 10144 4435 10200
rect 4491 10144 4559 10200
rect 4615 10144 4683 10200
rect 4739 10144 4807 10200
rect 4863 10144 4931 10200
rect 4987 10144 5055 10200
rect 5111 10144 5179 10200
rect 5235 10144 5303 10200
rect 5359 10144 5427 10200
rect 5483 10144 5551 10200
rect 5607 10144 5675 10200
rect 5731 10144 5799 10200
rect 5855 10144 5923 10200
rect 5979 10144 6047 10200
rect 6103 10144 6171 10200
rect 6227 10144 6237 10200
rect 4425 10076 6237 10144
rect 4425 10020 4435 10076
rect 4491 10020 4559 10076
rect 4615 10020 4683 10076
rect 4739 10020 4807 10076
rect 4863 10020 4931 10076
rect 4987 10020 5055 10076
rect 5111 10020 5179 10076
rect 5235 10020 5303 10076
rect 5359 10020 5427 10076
rect 5483 10020 5551 10076
rect 5607 10020 5675 10076
rect 5731 10020 5799 10076
rect 5855 10020 5923 10076
rect 5979 10020 6047 10076
rect 6103 10020 6171 10076
rect 6227 10020 6237 10076
rect 4425 9952 6237 10020
rect 4425 9896 4435 9952
rect 4491 9896 4559 9952
rect 4615 9896 4683 9952
rect 4739 9896 4807 9952
rect 4863 9896 4931 9952
rect 4987 9896 5055 9952
rect 5111 9896 5179 9952
rect 5235 9896 5303 9952
rect 5359 9896 5427 9952
rect 5483 9896 5551 9952
rect 5607 9896 5675 9952
rect 5731 9896 5799 9952
rect 5855 9896 5923 9952
rect 5979 9896 6047 9952
rect 6103 9896 6171 9952
rect 6227 9896 6237 9952
rect 4425 9828 6237 9896
rect 4425 9772 4435 9828
rect 4491 9772 4559 9828
rect 4615 9772 4683 9828
rect 4739 9772 4807 9828
rect 4863 9772 4931 9828
rect 4987 9772 5055 9828
rect 5111 9772 5179 9828
rect 5235 9772 5303 9828
rect 5359 9772 5427 9828
rect 5483 9772 5551 9828
rect 5607 9772 5675 9828
rect 5731 9772 5799 9828
rect 5855 9772 5923 9828
rect 5979 9772 6047 9828
rect 6103 9772 6171 9828
rect 6227 9772 6237 9828
rect 4425 9704 6237 9772
rect 4425 9648 4435 9704
rect 4491 9648 4559 9704
rect 4615 9648 4683 9704
rect 4739 9648 4807 9704
rect 4863 9648 4931 9704
rect 4987 9648 5055 9704
rect 5111 9648 5179 9704
rect 5235 9648 5303 9704
rect 5359 9648 5427 9704
rect 5483 9648 5551 9704
rect 5607 9648 5675 9704
rect 5731 9648 5799 9704
rect 5855 9648 5923 9704
rect 5979 9648 6047 9704
rect 6103 9648 6171 9704
rect 6227 9648 6237 9704
rect 4425 9638 6237 9648
rect 7552 10944 8620 10954
rect 7552 10888 7562 10944
rect 7618 10888 7686 10944
rect 7742 10888 7810 10944
rect 7866 10888 7934 10944
rect 7990 10888 8058 10944
rect 8114 10888 8182 10944
rect 8238 10888 8306 10944
rect 8362 10888 8430 10944
rect 8486 10888 8554 10944
rect 8610 10888 8620 10944
rect 7552 10820 8620 10888
rect 7552 10764 7562 10820
rect 7618 10764 7686 10820
rect 7742 10764 7810 10820
rect 7866 10764 7934 10820
rect 7990 10764 8058 10820
rect 8114 10764 8182 10820
rect 8238 10764 8306 10820
rect 8362 10764 8430 10820
rect 8486 10764 8554 10820
rect 8610 10764 8620 10820
rect 7552 10696 8620 10764
rect 7552 10640 7562 10696
rect 7618 10640 7686 10696
rect 7742 10640 7810 10696
rect 7866 10640 7934 10696
rect 7990 10640 8058 10696
rect 8114 10640 8182 10696
rect 8238 10640 8306 10696
rect 8362 10640 8430 10696
rect 8486 10640 8554 10696
rect 8610 10640 8620 10696
rect 7552 10572 8620 10640
rect 7552 10516 7562 10572
rect 7618 10516 7686 10572
rect 7742 10516 7810 10572
rect 7866 10516 7934 10572
rect 7990 10516 8058 10572
rect 8114 10516 8182 10572
rect 8238 10516 8306 10572
rect 8362 10516 8430 10572
rect 8486 10516 8554 10572
rect 8610 10516 8620 10572
rect 7552 10448 8620 10516
rect 7552 10392 7562 10448
rect 7618 10392 7686 10448
rect 7742 10392 7810 10448
rect 7866 10392 7934 10448
rect 7990 10392 8058 10448
rect 8114 10392 8182 10448
rect 8238 10392 8306 10448
rect 8362 10392 8430 10448
rect 8486 10392 8554 10448
rect 8610 10392 8620 10448
rect 7552 10324 8620 10392
rect 7552 10268 7562 10324
rect 7618 10268 7686 10324
rect 7742 10268 7810 10324
rect 7866 10268 7934 10324
rect 7990 10268 8058 10324
rect 8114 10268 8182 10324
rect 8238 10268 8306 10324
rect 8362 10268 8430 10324
rect 8486 10268 8554 10324
rect 8610 10268 8620 10324
rect 7552 10200 8620 10268
rect 7552 10144 7562 10200
rect 7618 10144 7686 10200
rect 7742 10144 7810 10200
rect 7866 10144 7934 10200
rect 7990 10144 8058 10200
rect 8114 10144 8182 10200
rect 8238 10144 8306 10200
rect 8362 10144 8430 10200
rect 8486 10144 8554 10200
rect 8610 10144 8620 10200
rect 7552 10076 8620 10144
rect 7552 10020 7562 10076
rect 7618 10020 7686 10076
rect 7742 10020 7810 10076
rect 7866 10020 7934 10076
rect 7990 10020 8058 10076
rect 8114 10020 8182 10076
rect 8238 10020 8306 10076
rect 8362 10020 8430 10076
rect 8486 10020 8554 10076
rect 8610 10020 8620 10076
rect 7552 9952 8620 10020
rect 7552 9896 7562 9952
rect 7618 9896 7686 9952
rect 7742 9896 7810 9952
rect 7866 9896 7934 9952
rect 7990 9896 8058 9952
rect 8114 9896 8182 9952
rect 8238 9896 8306 9952
rect 8362 9896 8430 9952
rect 8486 9896 8554 9952
rect 8610 9896 8620 9952
rect 7552 9828 8620 9896
rect 7552 9772 7562 9828
rect 7618 9772 7686 9828
rect 7742 9772 7810 9828
rect 7866 9772 7934 9828
rect 7990 9772 8058 9828
rect 8114 9772 8182 9828
rect 8238 9772 8306 9828
rect 8362 9772 8430 9828
rect 8486 9772 8554 9828
rect 8610 9772 8620 9828
rect 7552 9704 8620 9772
rect 7552 9648 7562 9704
rect 7618 9648 7686 9704
rect 7742 9648 7810 9704
rect 7866 9648 7934 9704
rect 7990 9648 8058 9704
rect 8114 9648 8182 9704
rect 8238 9648 8306 9704
rect 8362 9648 8430 9704
rect 8486 9648 8554 9704
rect 8610 9648 8620 9704
rect 7552 9638 8620 9648
rect 10669 10944 12481 10954
rect 10669 10888 10679 10944
rect 10735 10888 10803 10944
rect 10859 10888 10927 10944
rect 10983 10888 11051 10944
rect 11107 10888 11175 10944
rect 11231 10888 11299 10944
rect 11355 10888 11423 10944
rect 11479 10888 11547 10944
rect 11603 10888 11671 10944
rect 11727 10888 11795 10944
rect 11851 10888 11919 10944
rect 11975 10888 12043 10944
rect 12099 10888 12167 10944
rect 12223 10888 12291 10944
rect 12347 10888 12415 10944
rect 12471 10888 12481 10944
rect 10669 10820 12481 10888
rect 10669 10764 10679 10820
rect 10735 10764 10803 10820
rect 10859 10764 10927 10820
rect 10983 10764 11051 10820
rect 11107 10764 11175 10820
rect 11231 10764 11299 10820
rect 11355 10764 11423 10820
rect 11479 10764 11547 10820
rect 11603 10764 11671 10820
rect 11727 10764 11795 10820
rect 11851 10764 11919 10820
rect 11975 10764 12043 10820
rect 12099 10764 12167 10820
rect 12223 10764 12291 10820
rect 12347 10764 12415 10820
rect 12471 10764 12481 10820
rect 10669 10696 12481 10764
rect 10669 10640 10679 10696
rect 10735 10640 10803 10696
rect 10859 10640 10927 10696
rect 10983 10640 11051 10696
rect 11107 10640 11175 10696
rect 11231 10640 11299 10696
rect 11355 10640 11423 10696
rect 11479 10640 11547 10696
rect 11603 10640 11671 10696
rect 11727 10640 11795 10696
rect 11851 10640 11919 10696
rect 11975 10640 12043 10696
rect 12099 10640 12167 10696
rect 12223 10640 12291 10696
rect 12347 10640 12415 10696
rect 12471 10640 12481 10696
rect 10669 10572 12481 10640
rect 10669 10516 10679 10572
rect 10735 10516 10803 10572
rect 10859 10516 10927 10572
rect 10983 10516 11051 10572
rect 11107 10516 11175 10572
rect 11231 10516 11299 10572
rect 11355 10516 11423 10572
rect 11479 10516 11547 10572
rect 11603 10516 11671 10572
rect 11727 10516 11795 10572
rect 11851 10516 11919 10572
rect 11975 10516 12043 10572
rect 12099 10516 12167 10572
rect 12223 10516 12291 10572
rect 12347 10516 12415 10572
rect 12471 10516 12481 10572
rect 10669 10448 12481 10516
rect 10669 10392 10679 10448
rect 10735 10392 10803 10448
rect 10859 10392 10927 10448
rect 10983 10392 11051 10448
rect 11107 10392 11175 10448
rect 11231 10392 11299 10448
rect 11355 10392 11423 10448
rect 11479 10392 11547 10448
rect 11603 10392 11671 10448
rect 11727 10392 11795 10448
rect 11851 10392 11919 10448
rect 11975 10392 12043 10448
rect 12099 10392 12167 10448
rect 12223 10392 12291 10448
rect 12347 10392 12415 10448
rect 12471 10392 12481 10448
rect 10669 10324 12481 10392
rect 10669 10268 10679 10324
rect 10735 10268 10803 10324
rect 10859 10268 10927 10324
rect 10983 10268 11051 10324
rect 11107 10268 11175 10324
rect 11231 10268 11299 10324
rect 11355 10268 11423 10324
rect 11479 10268 11547 10324
rect 11603 10268 11671 10324
rect 11727 10268 11795 10324
rect 11851 10268 11919 10324
rect 11975 10268 12043 10324
rect 12099 10268 12167 10324
rect 12223 10268 12291 10324
rect 12347 10268 12415 10324
rect 12471 10268 12481 10324
rect 10669 10200 12481 10268
rect 10669 10144 10679 10200
rect 10735 10144 10803 10200
rect 10859 10144 10927 10200
rect 10983 10144 11051 10200
rect 11107 10144 11175 10200
rect 11231 10144 11299 10200
rect 11355 10144 11423 10200
rect 11479 10144 11547 10200
rect 11603 10144 11671 10200
rect 11727 10144 11795 10200
rect 11851 10144 11919 10200
rect 11975 10144 12043 10200
rect 12099 10144 12167 10200
rect 12223 10144 12291 10200
rect 12347 10144 12415 10200
rect 12471 10144 12481 10200
rect 10669 10076 12481 10144
rect 10669 10020 10679 10076
rect 10735 10020 10803 10076
rect 10859 10020 10927 10076
rect 10983 10020 11051 10076
rect 11107 10020 11175 10076
rect 11231 10020 11299 10076
rect 11355 10020 11423 10076
rect 11479 10020 11547 10076
rect 11603 10020 11671 10076
rect 11727 10020 11795 10076
rect 11851 10020 11919 10076
rect 11975 10020 12043 10076
rect 12099 10020 12167 10076
rect 12223 10020 12291 10076
rect 12347 10020 12415 10076
rect 12471 10020 12481 10076
rect 10669 9952 12481 10020
rect 10669 9896 10679 9952
rect 10735 9896 10803 9952
rect 10859 9896 10927 9952
rect 10983 9896 11051 9952
rect 11107 9896 11175 9952
rect 11231 9896 11299 9952
rect 11355 9896 11423 9952
rect 11479 9896 11547 9952
rect 11603 9896 11671 9952
rect 11727 9896 11795 9952
rect 11851 9896 11919 9952
rect 11975 9896 12043 9952
rect 12099 9896 12167 9952
rect 12223 9896 12291 9952
rect 12347 9896 12415 9952
rect 12471 9896 12481 9952
rect 10669 9828 12481 9896
rect 10669 9772 10679 9828
rect 10735 9772 10803 9828
rect 10859 9772 10927 9828
rect 10983 9772 11051 9828
rect 11107 9772 11175 9828
rect 11231 9772 11299 9828
rect 11355 9772 11423 9828
rect 11479 9772 11547 9828
rect 11603 9772 11671 9828
rect 11727 9772 11795 9828
rect 11851 9772 11919 9828
rect 11975 9772 12043 9828
rect 12099 9772 12167 9828
rect 12223 9772 12291 9828
rect 12347 9772 12415 9828
rect 12471 9772 12481 9828
rect 10669 9704 12481 9772
rect 10669 9648 10679 9704
rect 10735 9648 10803 9704
rect 10859 9648 10927 9704
rect 10983 9648 11051 9704
rect 11107 9648 11175 9704
rect 11231 9648 11299 9704
rect 11355 9648 11423 9704
rect 11479 9648 11547 9704
rect 11603 9648 11671 9704
rect 11727 9648 11795 9704
rect 11851 9648 11919 9704
rect 11975 9648 12043 9704
rect 12099 9648 12167 9704
rect 12223 9648 12291 9704
rect 12347 9648 12415 9704
rect 12471 9648 12481 9704
rect 10669 9638 12481 9648
rect 2497 9350 4309 9360
rect 2497 9294 2507 9350
rect 2563 9294 2631 9350
rect 2687 9294 2755 9350
rect 2811 9294 2879 9350
rect 2935 9294 3003 9350
rect 3059 9294 3127 9350
rect 3183 9294 3251 9350
rect 3307 9294 3375 9350
rect 3431 9294 3499 9350
rect 3555 9294 3623 9350
rect 3679 9294 3747 9350
rect 3803 9294 3871 9350
rect 3927 9294 3995 9350
rect 4051 9294 4119 9350
rect 4175 9294 4243 9350
rect 4299 9294 4309 9350
rect 2497 9226 4309 9294
rect 2497 9170 2507 9226
rect 2563 9170 2631 9226
rect 2687 9170 2755 9226
rect 2811 9170 2879 9226
rect 2935 9170 3003 9226
rect 3059 9170 3127 9226
rect 3183 9170 3251 9226
rect 3307 9170 3375 9226
rect 3431 9170 3499 9226
rect 3555 9170 3623 9226
rect 3679 9170 3747 9226
rect 3803 9170 3871 9226
rect 3927 9170 3995 9226
rect 4051 9170 4119 9226
rect 4175 9170 4243 9226
rect 4299 9170 4309 9226
rect 2497 9102 4309 9170
rect 2497 9046 2507 9102
rect 2563 9046 2631 9102
rect 2687 9046 2755 9102
rect 2811 9046 2879 9102
rect 2935 9046 3003 9102
rect 3059 9046 3127 9102
rect 3183 9046 3251 9102
rect 3307 9046 3375 9102
rect 3431 9046 3499 9102
rect 3555 9046 3623 9102
rect 3679 9046 3747 9102
rect 3803 9046 3871 9102
rect 3927 9046 3995 9102
rect 4051 9046 4119 9102
rect 4175 9046 4243 9102
rect 4299 9046 4309 9102
rect 2497 8978 4309 9046
rect 2497 8922 2507 8978
rect 2563 8922 2631 8978
rect 2687 8922 2755 8978
rect 2811 8922 2879 8978
rect 2935 8922 3003 8978
rect 3059 8922 3127 8978
rect 3183 8922 3251 8978
rect 3307 8922 3375 8978
rect 3431 8922 3499 8978
rect 3555 8922 3623 8978
rect 3679 8922 3747 8978
rect 3803 8922 3871 8978
rect 3927 8922 3995 8978
rect 4051 8922 4119 8978
rect 4175 8922 4243 8978
rect 4299 8922 4309 8978
rect 2497 8854 4309 8922
rect 2497 8798 2507 8854
rect 2563 8798 2631 8854
rect 2687 8798 2755 8854
rect 2811 8798 2879 8854
rect 2935 8798 3003 8854
rect 3059 8798 3127 8854
rect 3183 8798 3251 8854
rect 3307 8798 3375 8854
rect 3431 8798 3499 8854
rect 3555 8798 3623 8854
rect 3679 8798 3747 8854
rect 3803 8798 3871 8854
rect 3927 8798 3995 8854
rect 4051 8798 4119 8854
rect 4175 8798 4243 8854
rect 4299 8798 4309 8854
rect 2497 8730 4309 8798
rect 2497 8674 2507 8730
rect 2563 8674 2631 8730
rect 2687 8674 2755 8730
rect 2811 8674 2879 8730
rect 2935 8674 3003 8730
rect 3059 8674 3127 8730
rect 3183 8674 3251 8730
rect 3307 8674 3375 8730
rect 3431 8674 3499 8730
rect 3555 8674 3623 8730
rect 3679 8674 3747 8730
rect 3803 8674 3871 8730
rect 3927 8674 3995 8730
rect 4051 8674 4119 8730
rect 4175 8674 4243 8730
rect 4299 8674 4309 8730
rect 2497 8606 4309 8674
rect 2497 8550 2507 8606
rect 2563 8550 2631 8606
rect 2687 8550 2755 8606
rect 2811 8550 2879 8606
rect 2935 8550 3003 8606
rect 3059 8550 3127 8606
rect 3183 8550 3251 8606
rect 3307 8550 3375 8606
rect 3431 8550 3499 8606
rect 3555 8550 3623 8606
rect 3679 8550 3747 8606
rect 3803 8550 3871 8606
rect 3927 8550 3995 8606
rect 4051 8550 4119 8606
rect 4175 8550 4243 8606
rect 4299 8550 4309 8606
rect 2497 8482 4309 8550
rect 2497 8426 2507 8482
rect 2563 8426 2631 8482
rect 2687 8426 2755 8482
rect 2811 8426 2879 8482
rect 2935 8426 3003 8482
rect 3059 8426 3127 8482
rect 3183 8426 3251 8482
rect 3307 8426 3375 8482
rect 3431 8426 3499 8482
rect 3555 8426 3623 8482
rect 3679 8426 3747 8482
rect 3803 8426 3871 8482
rect 3927 8426 3995 8482
rect 4051 8426 4119 8482
rect 4175 8426 4243 8482
rect 4299 8426 4309 8482
rect 2497 8358 4309 8426
rect 2497 8302 2507 8358
rect 2563 8302 2631 8358
rect 2687 8302 2755 8358
rect 2811 8302 2879 8358
rect 2935 8302 3003 8358
rect 3059 8302 3127 8358
rect 3183 8302 3251 8358
rect 3307 8302 3375 8358
rect 3431 8302 3499 8358
rect 3555 8302 3623 8358
rect 3679 8302 3747 8358
rect 3803 8302 3871 8358
rect 3927 8302 3995 8358
rect 4051 8302 4119 8358
rect 4175 8302 4243 8358
rect 4299 8302 4309 8358
rect 2497 8234 4309 8302
rect 2497 8178 2507 8234
rect 2563 8178 2631 8234
rect 2687 8178 2755 8234
rect 2811 8178 2879 8234
rect 2935 8178 3003 8234
rect 3059 8178 3127 8234
rect 3183 8178 3251 8234
rect 3307 8178 3375 8234
rect 3431 8178 3499 8234
rect 3555 8178 3623 8234
rect 3679 8178 3747 8234
rect 3803 8178 3871 8234
rect 3927 8178 3995 8234
rect 4051 8178 4119 8234
rect 4175 8178 4243 8234
rect 4299 8178 4309 8234
rect 2497 8110 4309 8178
rect 2497 8054 2507 8110
rect 2563 8054 2631 8110
rect 2687 8054 2755 8110
rect 2811 8054 2879 8110
rect 2935 8054 3003 8110
rect 3059 8054 3127 8110
rect 3183 8054 3251 8110
rect 3307 8054 3375 8110
rect 3431 8054 3499 8110
rect 3555 8054 3623 8110
rect 3679 8054 3747 8110
rect 3803 8054 3871 8110
rect 3927 8054 3995 8110
rect 4051 8054 4119 8110
rect 4175 8054 4243 8110
rect 4299 8054 4309 8110
rect 2497 7986 4309 8054
rect 2497 7930 2507 7986
rect 2563 7930 2631 7986
rect 2687 7930 2755 7986
rect 2811 7930 2879 7986
rect 2935 7930 3003 7986
rect 3059 7930 3127 7986
rect 3183 7930 3251 7986
rect 3307 7930 3375 7986
rect 3431 7930 3499 7986
rect 3555 7930 3623 7986
rect 3679 7930 3747 7986
rect 3803 7930 3871 7986
rect 3927 7930 3995 7986
rect 4051 7930 4119 7986
rect 4175 7930 4243 7986
rect 4299 7930 4309 7986
rect 2497 7862 4309 7930
rect 2497 7806 2507 7862
rect 2563 7806 2631 7862
rect 2687 7806 2755 7862
rect 2811 7806 2879 7862
rect 2935 7806 3003 7862
rect 3059 7806 3127 7862
rect 3183 7806 3251 7862
rect 3307 7806 3375 7862
rect 3431 7806 3499 7862
rect 3555 7806 3623 7862
rect 3679 7806 3747 7862
rect 3803 7806 3871 7862
rect 3927 7806 3995 7862
rect 4051 7806 4119 7862
rect 4175 7806 4243 7862
rect 4299 7806 4309 7862
rect 2497 7738 4309 7806
rect 2497 7682 2507 7738
rect 2563 7682 2631 7738
rect 2687 7682 2755 7738
rect 2811 7682 2879 7738
rect 2935 7682 3003 7738
rect 3059 7682 3127 7738
rect 3183 7682 3251 7738
rect 3307 7682 3375 7738
rect 3431 7682 3499 7738
rect 3555 7682 3623 7738
rect 3679 7682 3747 7738
rect 3803 7682 3871 7738
rect 3927 7682 3995 7738
rect 4051 7682 4119 7738
rect 4175 7682 4243 7738
rect 4299 7682 4309 7738
rect 2497 7614 4309 7682
rect 2497 7558 2507 7614
rect 2563 7558 2631 7614
rect 2687 7558 2755 7614
rect 2811 7558 2879 7614
rect 2935 7558 3003 7614
rect 3059 7558 3127 7614
rect 3183 7558 3251 7614
rect 3307 7558 3375 7614
rect 3431 7558 3499 7614
rect 3555 7558 3623 7614
rect 3679 7558 3747 7614
rect 3803 7558 3871 7614
rect 3927 7558 3995 7614
rect 4051 7558 4119 7614
rect 4175 7558 4243 7614
rect 4299 7558 4309 7614
rect 2497 7490 4309 7558
rect 2497 7434 2507 7490
rect 2563 7434 2631 7490
rect 2687 7434 2755 7490
rect 2811 7434 2879 7490
rect 2935 7434 3003 7490
rect 3059 7434 3127 7490
rect 3183 7434 3251 7490
rect 3307 7434 3375 7490
rect 3431 7434 3499 7490
rect 3555 7434 3623 7490
rect 3679 7434 3747 7490
rect 3803 7434 3871 7490
rect 3927 7434 3995 7490
rect 4051 7434 4119 7490
rect 4175 7434 4243 7490
rect 4299 7434 4309 7490
rect 2497 7366 4309 7434
rect 2497 7310 2507 7366
rect 2563 7310 2631 7366
rect 2687 7310 2755 7366
rect 2811 7310 2879 7366
rect 2935 7310 3003 7366
rect 3059 7310 3127 7366
rect 3183 7310 3251 7366
rect 3307 7310 3375 7366
rect 3431 7310 3499 7366
rect 3555 7310 3623 7366
rect 3679 7310 3747 7366
rect 3803 7310 3871 7366
rect 3927 7310 3995 7366
rect 4051 7310 4119 7366
rect 4175 7310 4243 7366
rect 4299 7310 4309 7366
rect 2497 7242 4309 7310
rect 2497 7186 2507 7242
rect 2563 7186 2631 7242
rect 2687 7186 2755 7242
rect 2811 7186 2879 7242
rect 2935 7186 3003 7242
rect 3059 7186 3127 7242
rect 3183 7186 3251 7242
rect 3307 7186 3375 7242
rect 3431 7186 3499 7242
rect 3555 7186 3623 7242
rect 3679 7186 3747 7242
rect 3803 7186 3871 7242
rect 3927 7186 3995 7242
rect 4051 7186 4119 7242
rect 4175 7186 4243 7242
rect 4299 7186 4309 7242
rect 2497 7118 4309 7186
rect 2497 7062 2507 7118
rect 2563 7062 2631 7118
rect 2687 7062 2755 7118
rect 2811 7062 2879 7118
rect 2935 7062 3003 7118
rect 3059 7062 3127 7118
rect 3183 7062 3251 7118
rect 3307 7062 3375 7118
rect 3431 7062 3499 7118
rect 3555 7062 3623 7118
rect 3679 7062 3747 7118
rect 3803 7062 3871 7118
rect 3927 7062 3995 7118
rect 4051 7062 4119 7118
rect 4175 7062 4243 7118
rect 4299 7062 4309 7118
rect 2497 6994 4309 7062
rect 2497 6938 2507 6994
rect 2563 6938 2631 6994
rect 2687 6938 2755 6994
rect 2811 6938 2879 6994
rect 2935 6938 3003 6994
rect 3059 6938 3127 6994
rect 3183 6938 3251 6994
rect 3307 6938 3375 6994
rect 3431 6938 3499 6994
rect 3555 6938 3623 6994
rect 3679 6938 3747 6994
rect 3803 6938 3871 6994
rect 3927 6938 3995 6994
rect 4051 6938 4119 6994
rect 4175 6938 4243 6994
rect 4299 6938 4309 6994
rect 2497 6870 4309 6938
rect 2497 6814 2507 6870
rect 2563 6814 2631 6870
rect 2687 6814 2755 6870
rect 2811 6814 2879 6870
rect 2935 6814 3003 6870
rect 3059 6814 3127 6870
rect 3183 6814 3251 6870
rect 3307 6814 3375 6870
rect 3431 6814 3499 6870
rect 3555 6814 3623 6870
rect 3679 6814 3747 6870
rect 3803 6814 3871 6870
rect 3927 6814 3995 6870
rect 4051 6814 4119 6870
rect 4175 6814 4243 6870
rect 4299 6814 4309 6870
rect 2497 6746 4309 6814
rect 2497 6690 2507 6746
rect 2563 6690 2631 6746
rect 2687 6690 2755 6746
rect 2811 6690 2879 6746
rect 2935 6690 3003 6746
rect 3059 6690 3127 6746
rect 3183 6690 3251 6746
rect 3307 6690 3375 6746
rect 3431 6690 3499 6746
rect 3555 6690 3623 6746
rect 3679 6690 3747 6746
rect 3803 6690 3871 6746
rect 3927 6690 3995 6746
rect 4051 6690 4119 6746
rect 4175 6690 4243 6746
rect 4299 6690 4309 6746
rect 2497 6622 4309 6690
rect 2497 6566 2507 6622
rect 2563 6566 2631 6622
rect 2687 6566 2755 6622
rect 2811 6566 2879 6622
rect 2935 6566 3003 6622
rect 3059 6566 3127 6622
rect 3183 6566 3251 6622
rect 3307 6566 3375 6622
rect 3431 6566 3499 6622
rect 3555 6566 3623 6622
rect 3679 6566 3747 6622
rect 3803 6566 3871 6622
rect 3927 6566 3995 6622
rect 4051 6566 4119 6622
rect 4175 6566 4243 6622
rect 4299 6566 4309 6622
rect 2497 6498 4309 6566
rect 2497 6442 2507 6498
rect 2563 6442 2631 6498
rect 2687 6442 2755 6498
rect 2811 6442 2879 6498
rect 2935 6442 3003 6498
rect 3059 6442 3127 6498
rect 3183 6442 3251 6498
rect 3307 6442 3375 6498
rect 3431 6442 3499 6498
rect 3555 6442 3623 6498
rect 3679 6442 3747 6498
rect 3803 6442 3871 6498
rect 3927 6442 3995 6498
rect 4051 6442 4119 6498
rect 4175 6442 4243 6498
rect 4299 6442 4309 6498
rect 2497 6432 4309 6442
rect 6358 9350 7426 9360
rect 6358 9294 6368 9350
rect 6424 9294 6492 9350
rect 6548 9294 6616 9350
rect 6672 9294 6740 9350
rect 6796 9294 6864 9350
rect 6920 9294 6988 9350
rect 7044 9294 7112 9350
rect 7168 9294 7236 9350
rect 7292 9294 7360 9350
rect 7416 9294 7426 9350
rect 6358 9226 7426 9294
rect 6358 9170 6368 9226
rect 6424 9170 6492 9226
rect 6548 9170 6616 9226
rect 6672 9170 6740 9226
rect 6796 9170 6864 9226
rect 6920 9170 6988 9226
rect 7044 9170 7112 9226
rect 7168 9170 7236 9226
rect 7292 9170 7360 9226
rect 7416 9170 7426 9226
rect 6358 9102 7426 9170
rect 6358 9046 6368 9102
rect 6424 9046 6492 9102
rect 6548 9046 6616 9102
rect 6672 9046 6740 9102
rect 6796 9046 6864 9102
rect 6920 9046 6988 9102
rect 7044 9046 7112 9102
rect 7168 9046 7236 9102
rect 7292 9046 7360 9102
rect 7416 9046 7426 9102
rect 6358 8978 7426 9046
rect 6358 8922 6368 8978
rect 6424 8922 6492 8978
rect 6548 8922 6616 8978
rect 6672 8922 6740 8978
rect 6796 8922 6864 8978
rect 6920 8922 6988 8978
rect 7044 8922 7112 8978
rect 7168 8922 7236 8978
rect 7292 8922 7360 8978
rect 7416 8922 7426 8978
rect 6358 8854 7426 8922
rect 6358 8798 6368 8854
rect 6424 8798 6492 8854
rect 6548 8798 6616 8854
rect 6672 8798 6740 8854
rect 6796 8798 6864 8854
rect 6920 8798 6988 8854
rect 7044 8798 7112 8854
rect 7168 8798 7236 8854
rect 7292 8798 7360 8854
rect 7416 8798 7426 8854
rect 6358 8730 7426 8798
rect 6358 8674 6368 8730
rect 6424 8674 6492 8730
rect 6548 8674 6616 8730
rect 6672 8674 6740 8730
rect 6796 8674 6864 8730
rect 6920 8674 6988 8730
rect 7044 8674 7112 8730
rect 7168 8674 7236 8730
rect 7292 8674 7360 8730
rect 7416 8674 7426 8730
rect 6358 8606 7426 8674
rect 6358 8550 6368 8606
rect 6424 8550 6492 8606
rect 6548 8550 6616 8606
rect 6672 8550 6740 8606
rect 6796 8550 6864 8606
rect 6920 8550 6988 8606
rect 7044 8550 7112 8606
rect 7168 8550 7236 8606
rect 7292 8550 7360 8606
rect 7416 8550 7426 8606
rect 6358 8482 7426 8550
rect 6358 8426 6368 8482
rect 6424 8426 6492 8482
rect 6548 8426 6616 8482
rect 6672 8426 6740 8482
rect 6796 8426 6864 8482
rect 6920 8426 6988 8482
rect 7044 8426 7112 8482
rect 7168 8426 7236 8482
rect 7292 8426 7360 8482
rect 7416 8426 7426 8482
rect 6358 8358 7426 8426
rect 6358 8302 6368 8358
rect 6424 8302 6492 8358
rect 6548 8302 6616 8358
rect 6672 8302 6740 8358
rect 6796 8302 6864 8358
rect 6920 8302 6988 8358
rect 7044 8302 7112 8358
rect 7168 8302 7236 8358
rect 7292 8302 7360 8358
rect 7416 8302 7426 8358
rect 6358 8234 7426 8302
rect 6358 8178 6368 8234
rect 6424 8178 6492 8234
rect 6548 8178 6616 8234
rect 6672 8178 6740 8234
rect 6796 8178 6864 8234
rect 6920 8178 6988 8234
rect 7044 8178 7112 8234
rect 7168 8178 7236 8234
rect 7292 8178 7360 8234
rect 7416 8178 7426 8234
rect 6358 8110 7426 8178
rect 6358 8054 6368 8110
rect 6424 8054 6492 8110
rect 6548 8054 6616 8110
rect 6672 8054 6740 8110
rect 6796 8054 6864 8110
rect 6920 8054 6988 8110
rect 7044 8054 7112 8110
rect 7168 8054 7236 8110
rect 7292 8054 7360 8110
rect 7416 8054 7426 8110
rect 6358 7986 7426 8054
rect 6358 7930 6368 7986
rect 6424 7930 6492 7986
rect 6548 7930 6616 7986
rect 6672 7930 6740 7986
rect 6796 7930 6864 7986
rect 6920 7930 6988 7986
rect 7044 7930 7112 7986
rect 7168 7930 7236 7986
rect 7292 7930 7360 7986
rect 7416 7930 7426 7986
rect 6358 7862 7426 7930
rect 6358 7806 6368 7862
rect 6424 7806 6492 7862
rect 6548 7806 6616 7862
rect 6672 7806 6740 7862
rect 6796 7806 6864 7862
rect 6920 7806 6988 7862
rect 7044 7806 7112 7862
rect 7168 7806 7236 7862
rect 7292 7806 7360 7862
rect 7416 7806 7426 7862
rect 6358 7738 7426 7806
rect 6358 7682 6368 7738
rect 6424 7682 6492 7738
rect 6548 7682 6616 7738
rect 6672 7682 6740 7738
rect 6796 7682 6864 7738
rect 6920 7682 6988 7738
rect 7044 7682 7112 7738
rect 7168 7682 7236 7738
rect 7292 7682 7360 7738
rect 7416 7682 7426 7738
rect 6358 7614 7426 7682
rect 6358 7558 6368 7614
rect 6424 7558 6492 7614
rect 6548 7558 6616 7614
rect 6672 7558 6740 7614
rect 6796 7558 6864 7614
rect 6920 7558 6988 7614
rect 7044 7558 7112 7614
rect 7168 7558 7236 7614
rect 7292 7558 7360 7614
rect 7416 7558 7426 7614
rect 6358 7490 7426 7558
rect 6358 7434 6368 7490
rect 6424 7434 6492 7490
rect 6548 7434 6616 7490
rect 6672 7434 6740 7490
rect 6796 7434 6864 7490
rect 6920 7434 6988 7490
rect 7044 7434 7112 7490
rect 7168 7434 7236 7490
rect 7292 7434 7360 7490
rect 7416 7434 7426 7490
rect 6358 7366 7426 7434
rect 6358 7310 6368 7366
rect 6424 7310 6492 7366
rect 6548 7310 6616 7366
rect 6672 7310 6740 7366
rect 6796 7310 6864 7366
rect 6920 7310 6988 7366
rect 7044 7310 7112 7366
rect 7168 7310 7236 7366
rect 7292 7310 7360 7366
rect 7416 7310 7426 7366
rect 6358 7242 7426 7310
rect 6358 7186 6368 7242
rect 6424 7186 6492 7242
rect 6548 7186 6616 7242
rect 6672 7186 6740 7242
rect 6796 7186 6864 7242
rect 6920 7186 6988 7242
rect 7044 7186 7112 7242
rect 7168 7186 7236 7242
rect 7292 7186 7360 7242
rect 7416 7186 7426 7242
rect 6358 7118 7426 7186
rect 6358 7062 6368 7118
rect 6424 7062 6492 7118
rect 6548 7062 6616 7118
rect 6672 7062 6740 7118
rect 6796 7062 6864 7118
rect 6920 7062 6988 7118
rect 7044 7062 7112 7118
rect 7168 7062 7236 7118
rect 7292 7062 7360 7118
rect 7416 7062 7426 7118
rect 6358 6994 7426 7062
rect 6358 6938 6368 6994
rect 6424 6938 6492 6994
rect 6548 6938 6616 6994
rect 6672 6938 6740 6994
rect 6796 6938 6864 6994
rect 6920 6938 6988 6994
rect 7044 6938 7112 6994
rect 7168 6938 7236 6994
rect 7292 6938 7360 6994
rect 7416 6938 7426 6994
rect 6358 6870 7426 6938
rect 6358 6814 6368 6870
rect 6424 6814 6492 6870
rect 6548 6814 6616 6870
rect 6672 6814 6740 6870
rect 6796 6814 6864 6870
rect 6920 6814 6988 6870
rect 7044 6814 7112 6870
rect 7168 6814 7236 6870
rect 7292 6814 7360 6870
rect 7416 6814 7426 6870
rect 6358 6746 7426 6814
rect 6358 6690 6368 6746
rect 6424 6690 6492 6746
rect 6548 6690 6616 6746
rect 6672 6690 6740 6746
rect 6796 6690 6864 6746
rect 6920 6690 6988 6746
rect 7044 6690 7112 6746
rect 7168 6690 7236 6746
rect 7292 6690 7360 6746
rect 7416 6690 7426 6746
rect 6358 6622 7426 6690
rect 6358 6566 6368 6622
rect 6424 6566 6492 6622
rect 6548 6566 6616 6622
rect 6672 6566 6740 6622
rect 6796 6566 6864 6622
rect 6920 6566 6988 6622
rect 7044 6566 7112 6622
rect 7168 6566 7236 6622
rect 7292 6566 7360 6622
rect 7416 6566 7426 6622
rect 6358 6498 7426 6566
rect 6358 6442 6368 6498
rect 6424 6442 6492 6498
rect 6548 6442 6616 6498
rect 6672 6442 6740 6498
rect 6796 6442 6864 6498
rect 6920 6442 6988 6498
rect 7044 6442 7112 6498
rect 7168 6442 7236 6498
rect 7292 6442 7360 6498
rect 7416 6442 7426 6498
rect 6358 6432 7426 6442
rect 8741 9350 10553 9360
rect 8741 9294 8751 9350
rect 8807 9294 8875 9350
rect 8931 9294 8999 9350
rect 9055 9294 9123 9350
rect 9179 9294 9247 9350
rect 9303 9294 9371 9350
rect 9427 9294 9495 9350
rect 9551 9294 9619 9350
rect 9675 9294 9743 9350
rect 9799 9294 9867 9350
rect 9923 9294 9991 9350
rect 10047 9294 10115 9350
rect 10171 9294 10239 9350
rect 10295 9294 10363 9350
rect 10419 9294 10487 9350
rect 10543 9294 10553 9350
rect 8741 9226 10553 9294
rect 8741 9170 8751 9226
rect 8807 9170 8875 9226
rect 8931 9170 8999 9226
rect 9055 9170 9123 9226
rect 9179 9170 9247 9226
rect 9303 9170 9371 9226
rect 9427 9170 9495 9226
rect 9551 9170 9619 9226
rect 9675 9170 9743 9226
rect 9799 9170 9867 9226
rect 9923 9170 9991 9226
rect 10047 9170 10115 9226
rect 10171 9170 10239 9226
rect 10295 9170 10363 9226
rect 10419 9170 10487 9226
rect 10543 9170 10553 9226
rect 8741 9102 10553 9170
rect 8741 9046 8751 9102
rect 8807 9046 8875 9102
rect 8931 9046 8999 9102
rect 9055 9046 9123 9102
rect 9179 9046 9247 9102
rect 9303 9046 9371 9102
rect 9427 9046 9495 9102
rect 9551 9046 9619 9102
rect 9675 9046 9743 9102
rect 9799 9046 9867 9102
rect 9923 9046 9991 9102
rect 10047 9046 10115 9102
rect 10171 9046 10239 9102
rect 10295 9046 10363 9102
rect 10419 9046 10487 9102
rect 10543 9046 10553 9102
rect 8741 8978 10553 9046
rect 8741 8922 8751 8978
rect 8807 8922 8875 8978
rect 8931 8922 8999 8978
rect 9055 8922 9123 8978
rect 9179 8922 9247 8978
rect 9303 8922 9371 8978
rect 9427 8922 9495 8978
rect 9551 8922 9619 8978
rect 9675 8922 9743 8978
rect 9799 8922 9867 8978
rect 9923 8922 9991 8978
rect 10047 8922 10115 8978
rect 10171 8922 10239 8978
rect 10295 8922 10363 8978
rect 10419 8922 10487 8978
rect 10543 8922 10553 8978
rect 8741 8854 10553 8922
rect 8741 8798 8751 8854
rect 8807 8798 8875 8854
rect 8931 8798 8999 8854
rect 9055 8798 9123 8854
rect 9179 8798 9247 8854
rect 9303 8798 9371 8854
rect 9427 8798 9495 8854
rect 9551 8798 9619 8854
rect 9675 8798 9743 8854
rect 9799 8798 9867 8854
rect 9923 8798 9991 8854
rect 10047 8798 10115 8854
rect 10171 8798 10239 8854
rect 10295 8798 10363 8854
rect 10419 8798 10487 8854
rect 10543 8798 10553 8854
rect 8741 8730 10553 8798
rect 8741 8674 8751 8730
rect 8807 8674 8875 8730
rect 8931 8674 8999 8730
rect 9055 8674 9123 8730
rect 9179 8674 9247 8730
rect 9303 8674 9371 8730
rect 9427 8674 9495 8730
rect 9551 8674 9619 8730
rect 9675 8674 9743 8730
rect 9799 8674 9867 8730
rect 9923 8674 9991 8730
rect 10047 8674 10115 8730
rect 10171 8674 10239 8730
rect 10295 8674 10363 8730
rect 10419 8674 10487 8730
rect 10543 8674 10553 8730
rect 8741 8606 10553 8674
rect 8741 8550 8751 8606
rect 8807 8550 8875 8606
rect 8931 8550 8999 8606
rect 9055 8550 9123 8606
rect 9179 8550 9247 8606
rect 9303 8550 9371 8606
rect 9427 8550 9495 8606
rect 9551 8550 9619 8606
rect 9675 8550 9743 8606
rect 9799 8550 9867 8606
rect 9923 8550 9991 8606
rect 10047 8550 10115 8606
rect 10171 8550 10239 8606
rect 10295 8550 10363 8606
rect 10419 8550 10487 8606
rect 10543 8550 10553 8606
rect 8741 8482 10553 8550
rect 8741 8426 8751 8482
rect 8807 8426 8875 8482
rect 8931 8426 8999 8482
rect 9055 8426 9123 8482
rect 9179 8426 9247 8482
rect 9303 8426 9371 8482
rect 9427 8426 9495 8482
rect 9551 8426 9619 8482
rect 9675 8426 9743 8482
rect 9799 8426 9867 8482
rect 9923 8426 9991 8482
rect 10047 8426 10115 8482
rect 10171 8426 10239 8482
rect 10295 8426 10363 8482
rect 10419 8426 10487 8482
rect 10543 8426 10553 8482
rect 8741 8358 10553 8426
rect 8741 8302 8751 8358
rect 8807 8302 8875 8358
rect 8931 8302 8999 8358
rect 9055 8302 9123 8358
rect 9179 8302 9247 8358
rect 9303 8302 9371 8358
rect 9427 8302 9495 8358
rect 9551 8302 9619 8358
rect 9675 8302 9743 8358
rect 9799 8302 9867 8358
rect 9923 8302 9991 8358
rect 10047 8302 10115 8358
rect 10171 8302 10239 8358
rect 10295 8302 10363 8358
rect 10419 8302 10487 8358
rect 10543 8302 10553 8358
rect 8741 8234 10553 8302
rect 8741 8178 8751 8234
rect 8807 8178 8875 8234
rect 8931 8178 8999 8234
rect 9055 8178 9123 8234
rect 9179 8178 9247 8234
rect 9303 8178 9371 8234
rect 9427 8178 9495 8234
rect 9551 8178 9619 8234
rect 9675 8178 9743 8234
rect 9799 8178 9867 8234
rect 9923 8178 9991 8234
rect 10047 8178 10115 8234
rect 10171 8178 10239 8234
rect 10295 8178 10363 8234
rect 10419 8178 10487 8234
rect 10543 8178 10553 8234
rect 8741 8110 10553 8178
rect 8741 8054 8751 8110
rect 8807 8054 8875 8110
rect 8931 8054 8999 8110
rect 9055 8054 9123 8110
rect 9179 8054 9247 8110
rect 9303 8054 9371 8110
rect 9427 8054 9495 8110
rect 9551 8054 9619 8110
rect 9675 8054 9743 8110
rect 9799 8054 9867 8110
rect 9923 8054 9991 8110
rect 10047 8054 10115 8110
rect 10171 8054 10239 8110
rect 10295 8054 10363 8110
rect 10419 8054 10487 8110
rect 10543 8054 10553 8110
rect 8741 7986 10553 8054
rect 8741 7930 8751 7986
rect 8807 7930 8875 7986
rect 8931 7930 8999 7986
rect 9055 7930 9123 7986
rect 9179 7930 9247 7986
rect 9303 7930 9371 7986
rect 9427 7930 9495 7986
rect 9551 7930 9619 7986
rect 9675 7930 9743 7986
rect 9799 7930 9867 7986
rect 9923 7930 9991 7986
rect 10047 7930 10115 7986
rect 10171 7930 10239 7986
rect 10295 7930 10363 7986
rect 10419 7930 10487 7986
rect 10543 7930 10553 7986
rect 8741 7862 10553 7930
rect 8741 7806 8751 7862
rect 8807 7806 8875 7862
rect 8931 7806 8999 7862
rect 9055 7806 9123 7862
rect 9179 7806 9247 7862
rect 9303 7806 9371 7862
rect 9427 7806 9495 7862
rect 9551 7806 9619 7862
rect 9675 7806 9743 7862
rect 9799 7806 9867 7862
rect 9923 7806 9991 7862
rect 10047 7806 10115 7862
rect 10171 7806 10239 7862
rect 10295 7806 10363 7862
rect 10419 7806 10487 7862
rect 10543 7806 10553 7862
rect 8741 7738 10553 7806
rect 8741 7682 8751 7738
rect 8807 7682 8875 7738
rect 8931 7682 8999 7738
rect 9055 7682 9123 7738
rect 9179 7682 9247 7738
rect 9303 7682 9371 7738
rect 9427 7682 9495 7738
rect 9551 7682 9619 7738
rect 9675 7682 9743 7738
rect 9799 7682 9867 7738
rect 9923 7682 9991 7738
rect 10047 7682 10115 7738
rect 10171 7682 10239 7738
rect 10295 7682 10363 7738
rect 10419 7682 10487 7738
rect 10543 7682 10553 7738
rect 8741 7614 10553 7682
rect 8741 7558 8751 7614
rect 8807 7558 8875 7614
rect 8931 7558 8999 7614
rect 9055 7558 9123 7614
rect 9179 7558 9247 7614
rect 9303 7558 9371 7614
rect 9427 7558 9495 7614
rect 9551 7558 9619 7614
rect 9675 7558 9743 7614
rect 9799 7558 9867 7614
rect 9923 7558 9991 7614
rect 10047 7558 10115 7614
rect 10171 7558 10239 7614
rect 10295 7558 10363 7614
rect 10419 7558 10487 7614
rect 10543 7558 10553 7614
rect 8741 7490 10553 7558
rect 8741 7434 8751 7490
rect 8807 7434 8875 7490
rect 8931 7434 8999 7490
rect 9055 7434 9123 7490
rect 9179 7434 9247 7490
rect 9303 7434 9371 7490
rect 9427 7434 9495 7490
rect 9551 7434 9619 7490
rect 9675 7434 9743 7490
rect 9799 7434 9867 7490
rect 9923 7434 9991 7490
rect 10047 7434 10115 7490
rect 10171 7434 10239 7490
rect 10295 7434 10363 7490
rect 10419 7434 10487 7490
rect 10543 7434 10553 7490
rect 8741 7366 10553 7434
rect 8741 7310 8751 7366
rect 8807 7310 8875 7366
rect 8931 7310 8999 7366
rect 9055 7310 9123 7366
rect 9179 7310 9247 7366
rect 9303 7310 9371 7366
rect 9427 7310 9495 7366
rect 9551 7310 9619 7366
rect 9675 7310 9743 7366
rect 9799 7310 9867 7366
rect 9923 7310 9991 7366
rect 10047 7310 10115 7366
rect 10171 7310 10239 7366
rect 10295 7310 10363 7366
rect 10419 7310 10487 7366
rect 10543 7310 10553 7366
rect 8741 7242 10553 7310
rect 8741 7186 8751 7242
rect 8807 7186 8875 7242
rect 8931 7186 8999 7242
rect 9055 7186 9123 7242
rect 9179 7186 9247 7242
rect 9303 7186 9371 7242
rect 9427 7186 9495 7242
rect 9551 7186 9619 7242
rect 9675 7186 9743 7242
rect 9799 7186 9867 7242
rect 9923 7186 9991 7242
rect 10047 7186 10115 7242
rect 10171 7186 10239 7242
rect 10295 7186 10363 7242
rect 10419 7186 10487 7242
rect 10543 7186 10553 7242
rect 8741 7118 10553 7186
rect 8741 7062 8751 7118
rect 8807 7062 8875 7118
rect 8931 7062 8999 7118
rect 9055 7062 9123 7118
rect 9179 7062 9247 7118
rect 9303 7062 9371 7118
rect 9427 7062 9495 7118
rect 9551 7062 9619 7118
rect 9675 7062 9743 7118
rect 9799 7062 9867 7118
rect 9923 7062 9991 7118
rect 10047 7062 10115 7118
rect 10171 7062 10239 7118
rect 10295 7062 10363 7118
rect 10419 7062 10487 7118
rect 10543 7062 10553 7118
rect 8741 6994 10553 7062
rect 8741 6938 8751 6994
rect 8807 6938 8875 6994
rect 8931 6938 8999 6994
rect 9055 6938 9123 6994
rect 9179 6938 9247 6994
rect 9303 6938 9371 6994
rect 9427 6938 9495 6994
rect 9551 6938 9619 6994
rect 9675 6938 9743 6994
rect 9799 6938 9867 6994
rect 9923 6938 9991 6994
rect 10047 6938 10115 6994
rect 10171 6938 10239 6994
rect 10295 6938 10363 6994
rect 10419 6938 10487 6994
rect 10543 6938 10553 6994
rect 8741 6870 10553 6938
rect 8741 6814 8751 6870
rect 8807 6814 8875 6870
rect 8931 6814 8999 6870
rect 9055 6814 9123 6870
rect 9179 6814 9247 6870
rect 9303 6814 9371 6870
rect 9427 6814 9495 6870
rect 9551 6814 9619 6870
rect 9675 6814 9743 6870
rect 9799 6814 9867 6870
rect 9923 6814 9991 6870
rect 10047 6814 10115 6870
rect 10171 6814 10239 6870
rect 10295 6814 10363 6870
rect 10419 6814 10487 6870
rect 10543 6814 10553 6870
rect 8741 6746 10553 6814
rect 8741 6690 8751 6746
rect 8807 6690 8875 6746
rect 8931 6690 8999 6746
rect 9055 6690 9123 6746
rect 9179 6690 9247 6746
rect 9303 6690 9371 6746
rect 9427 6690 9495 6746
rect 9551 6690 9619 6746
rect 9675 6690 9743 6746
rect 9799 6690 9867 6746
rect 9923 6690 9991 6746
rect 10047 6690 10115 6746
rect 10171 6690 10239 6746
rect 10295 6690 10363 6746
rect 10419 6690 10487 6746
rect 10543 6690 10553 6746
rect 8741 6622 10553 6690
rect 8741 6566 8751 6622
rect 8807 6566 8875 6622
rect 8931 6566 8999 6622
rect 9055 6566 9123 6622
rect 9179 6566 9247 6622
rect 9303 6566 9371 6622
rect 9427 6566 9495 6622
rect 9551 6566 9619 6622
rect 9675 6566 9743 6622
rect 9799 6566 9867 6622
rect 9923 6566 9991 6622
rect 10047 6566 10115 6622
rect 10171 6566 10239 6622
rect 10295 6566 10363 6622
rect 10419 6566 10487 6622
rect 10543 6566 10553 6622
rect 8741 6498 10553 6566
rect 8741 6442 8751 6498
rect 8807 6442 8875 6498
rect 8931 6442 8999 6498
rect 9055 6442 9123 6498
rect 9179 6442 9247 6498
rect 9303 6442 9371 6498
rect 9427 6442 9495 6498
rect 9551 6442 9619 6498
rect 9675 6442 9743 6498
rect 9799 6442 9867 6498
rect 9923 6442 9991 6498
rect 10047 6442 10115 6498
rect 10171 6442 10239 6498
rect 10295 6442 10363 6498
rect 10419 6442 10487 6498
rect 10543 6442 10553 6498
rect 8741 6432 10553 6442
rect 12842 9350 13910 9360
rect 12842 9294 12852 9350
rect 12908 9294 12976 9350
rect 13032 9294 13100 9350
rect 13156 9294 13224 9350
rect 13280 9294 13348 9350
rect 13404 9294 13472 9350
rect 13528 9294 13596 9350
rect 13652 9294 13720 9350
rect 13776 9294 13844 9350
rect 13900 9294 13910 9350
rect 12842 9226 13910 9294
rect 12842 9170 12852 9226
rect 12908 9170 12976 9226
rect 13032 9170 13100 9226
rect 13156 9170 13224 9226
rect 13280 9170 13348 9226
rect 13404 9170 13472 9226
rect 13528 9170 13596 9226
rect 13652 9170 13720 9226
rect 13776 9170 13844 9226
rect 13900 9170 13910 9226
rect 12842 9102 13910 9170
rect 12842 9046 12852 9102
rect 12908 9046 12976 9102
rect 13032 9046 13100 9102
rect 13156 9046 13224 9102
rect 13280 9046 13348 9102
rect 13404 9046 13472 9102
rect 13528 9046 13596 9102
rect 13652 9046 13720 9102
rect 13776 9046 13844 9102
rect 13900 9046 13910 9102
rect 12842 8978 13910 9046
rect 12842 8922 12852 8978
rect 12908 8922 12976 8978
rect 13032 8922 13100 8978
rect 13156 8922 13224 8978
rect 13280 8922 13348 8978
rect 13404 8922 13472 8978
rect 13528 8922 13596 8978
rect 13652 8922 13720 8978
rect 13776 8922 13844 8978
rect 13900 8922 13910 8978
rect 12842 8854 13910 8922
rect 12842 8798 12852 8854
rect 12908 8798 12976 8854
rect 13032 8798 13100 8854
rect 13156 8798 13224 8854
rect 13280 8798 13348 8854
rect 13404 8798 13472 8854
rect 13528 8798 13596 8854
rect 13652 8798 13720 8854
rect 13776 8798 13844 8854
rect 13900 8798 13910 8854
rect 12842 8730 13910 8798
rect 12842 8674 12852 8730
rect 12908 8674 12976 8730
rect 13032 8674 13100 8730
rect 13156 8674 13224 8730
rect 13280 8674 13348 8730
rect 13404 8674 13472 8730
rect 13528 8674 13596 8730
rect 13652 8674 13720 8730
rect 13776 8674 13844 8730
rect 13900 8674 13910 8730
rect 12842 8606 13910 8674
rect 12842 8550 12852 8606
rect 12908 8550 12976 8606
rect 13032 8550 13100 8606
rect 13156 8550 13224 8606
rect 13280 8550 13348 8606
rect 13404 8550 13472 8606
rect 13528 8550 13596 8606
rect 13652 8550 13720 8606
rect 13776 8550 13844 8606
rect 13900 8550 13910 8606
rect 12842 8482 13910 8550
rect 12842 8426 12852 8482
rect 12908 8426 12976 8482
rect 13032 8426 13100 8482
rect 13156 8426 13224 8482
rect 13280 8426 13348 8482
rect 13404 8426 13472 8482
rect 13528 8426 13596 8482
rect 13652 8426 13720 8482
rect 13776 8426 13844 8482
rect 13900 8426 13910 8482
rect 12842 8358 13910 8426
rect 12842 8302 12852 8358
rect 12908 8302 12976 8358
rect 13032 8302 13100 8358
rect 13156 8302 13224 8358
rect 13280 8302 13348 8358
rect 13404 8302 13472 8358
rect 13528 8302 13596 8358
rect 13652 8302 13720 8358
rect 13776 8302 13844 8358
rect 13900 8302 13910 8358
rect 12842 8234 13910 8302
rect 12842 8178 12852 8234
rect 12908 8178 12976 8234
rect 13032 8178 13100 8234
rect 13156 8178 13224 8234
rect 13280 8178 13348 8234
rect 13404 8178 13472 8234
rect 13528 8178 13596 8234
rect 13652 8178 13720 8234
rect 13776 8178 13844 8234
rect 13900 8178 13910 8234
rect 12842 8110 13910 8178
rect 12842 8054 12852 8110
rect 12908 8054 12976 8110
rect 13032 8054 13100 8110
rect 13156 8054 13224 8110
rect 13280 8054 13348 8110
rect 13404 8054 13472 8110
rect 13528 8054 13596 8110
rect 13652 8054 13720 8110
rect 13776 8054 13844 8110
rect 13900 8054 13910 8110
rect 12842 7986 13910 8054
rect 12842 7930 12852 7986
rect 12908 7930 12976 7986
rect 13032 7930 13100 7986
rect 13156 7930 13224 7986
rect 13280 7930 13348 7986
rect 13404 7930 13472 7986
rect 13528 7930 13596 7986
rect 13652 7930 13720 7986
rect 13776 7930 13844 7986
rect 13900 7930 13910 7986
rect 12842 7862 13910 7930
rect 12842 7806 12852 7862
rect 12908 7806 12976 7862
rect 13032 7806 13100 7862
rect 13156 7806 13224 7862
rect 13280 7806 13348 7862
rect 13404 7806 13472 7862
rect 13528 7806 13596 7862
rect 13652 7806 13720 7862
rect 13776 7806 13844 7862
rect 13900 7806 13910 7862
rect 12842 7738 13910 7806
rect 12842 7682 12852 7738
rect 12908 7682 12976 7738
rect 13032 7682 13100 7738
rect 13156 7682 13224 7738
rect 13280 7682 13348 7738
rect 13404 7682 13472 7738
rect 13528 7682 13596 7738
rect 13652 7682 13720 7738
rect 13776 7682 13844 7738
rect 13900 7682 13910 7738
rect 12842 7614 13910 7682
rect 12842 7558 12852 7614
rect 12908 7558 12976 7614
rect 13032 7558 13100 7614
rect 13156 7558 13224 7614
rect 13280 7558 13348 7614
rect 13404 7558 13472 7614
rect 13528 7558 13596 7614
rect 13652 7558 13720 7614
rect 13776 7558 13844 7614
rect 13900 7558 13910 7614
rect 12842 7490 13910 7558
rect 12842 7434 12852 7490
rect 12908 7434 12976 7490
rect 13032 7434 13100 7490
rect 13156 7434 13224 7490
rect 13280 7434 13348 7490
rect 13404 7434 13472 7490
rect 13528 7434 13596 7490
rect 13652 7434 13720 7490
rect 13776 7434 13844 7490
rect 13900 7434 13910 7490
rect 12842 7366 13910 7434
rect 12842 7310 12852 7366
rect 12908 7310 12976 7366
rect 13032 7310 13100 7366
rect 13156 7310 13224 7366
rect 13280 7310 13348 7366
rect 13404 7310 13472 7366
rect 13528 7310 13596 7366
rect 13652 7310 13720 7366
rect 13776 7310 13844 7366
rect 13900 7310 13910 7366
rect 12842 7242 13910 7310
rect 12842 7186 12852 7242
rect 12908 7186 12976 7242
rect 13032 7186 13100 7242
rect 13156 7186 13224 7242
rect 13280 7186 13348 7242
rect 13404 7186 13472 7242
rect 13528 7186 13596 7242
rect 13652 7186 13720 7242
rect 13776 7186 13844 7242
rect 13900 7186 13910 7242
rect 12842 7118 13910 7186
rect 12842 7062 12852 7118
rect 12908 7062 12976 7118
rect 13032 7062 13100 7118
rect 13156 7062 13224 7118
rect 13280 7062 13348 7118
rect 13404 7062 13472 7118
rect 13528 7062 13596 7118
rect 13652 7062 13720 7118
rect 13776 7062 13844 7118
rect 13900 7062 13910 7118
rect 12842 6994 13910 7062
rect 12842 6938 12852 6994
rect 12908 6938 12976 6994
rect 13032 6938 13100 6994
rect 13156 6938 13224 6994
rect 13280 6938 13348 6994
rect 13404 6938 13472 6994
rect 13528 6938 13596 6994
rect 13652 6938 13720 6994
rect 13776 6938 13844 6994
rect 13900 6938 13910 6994
rect 12842 6870 13910 6938
rect 12842 6814 12852 6870
rect 12908 6814 12976 6870
rect 13032 6814 13100 6870
rect 13156 6814 13224 6870
rect 13280 6814 13348 6870
rect 13404 6814 13472 6870
rect 13528 6814 13596 6870
rect 13652 6814 13720 6870
rect 13776 6814 13844 6870
rect 13900 6814 13910 6870
rect 12842 6746 13910 6814
rect 12842 6690 12852 6746
rect 12908 6690 12976 6746
rect 13032 6690 13100 6746
rect 13156 6690 13224 6746
rect 13280 6690 13348 6746
rect 13404 6690 13472 6746
rect 13528 6690 13596 6746
rect 13652 6690 13720 6746
rect 13776 6690 13844 6746
rect 13900 6690 13910 6746
rect 12842 6622 13910 6690
rect 12842 6566 12852 6622
rect 12908 6566 12976 6622
rect 13032 6566 13100 6622
rect 13156 6566 13224 6622
rect 13280 6566 13348 6622
rect 13404 6566 13472 6622
rect 13528 6566 13596 6622
rect 13652 6566 13720 6622
rect 13776 6566 13844 6622
rect 13900 6566 13910 6622
rect 12842 6498 13910 6566
rect 12842 6442 12852 6498
rect 12908 6442 12976 6498
rect 13032 6442 13100 6498
rect 13156 6442 13224 6498
rect 13280 6442 13348 6498
rect 13404 6442 13472 6498
rect 13528 6442 13596 6498
rect 13652 6442 13720 6498
rect 13776 6442 13844 6498
rect 13900 6442 13910 6498
rect 12842 6432 13910 6442
rect 2497 6150 4309 6160
rect 2497 6094 2507 6150
rect 2563 6094 2631 6150
rect 2687 6094 2755 6150
rect 2811 6094 2879 6150
rect 2935 6094 3003 6150
rect 3059 6094 3127 6150
rect 3183 6094 3251 6150
rect 3307 6094 3375 6150
rect 3431 6094 3499 6150
rect 3555 6094 3623 6150
rect 3679 6094 3747 6150
rect 3803 6094 3871 6150
rect 3927 6094 3995 6150
rect 4051 6094 4119 6150
rect 4175 6094 4243 6150
rect 4299 6094 4309 6150
rect 2497 6026 4309 6094
rect 2497 5970 2507 6026
rect 2563 5970 2631 6026
rect 2687 5970 2755 6026
rect 2811 5970 2879 6026
rect 2935 5970 3003 6026
rect 3059 5970 3127 6026
rect 3183 5970 3251 6026
rect 3307 5970 3375 6026
rect 3431 5970 3499 6026
rect 3555 5970 3623 6026
rect 3679 5970 3747 6026
rect 3803 5970 3871 6026
rect 3927 5970 3995 6026
rect 4051 5970 4119 6026
rect 4175 5970 4243 6026
rect 4299 5970 4309 6026
rect 2497 5902 4309 5970
rect 2497 5846 2507 5902
rect 2563 5846 2631 5902
rect 2687 5846 2755 5902
rect 2811 5846 2879 5902
rect 2935 5846 3003 5902
rect 3059 5846 3127 5902
rect 3183 5846 3251 5902
rect 3307 5846 3375 5902
rect 3431 5846 3499 5902
rect 3555 5846 3623 5902
rect 3679 5846 3747 5902
rect 3803 5846 3871 5902
rect 3927 5846 3995 5902
rect 4051 5846 4119 5902
rect 4175 5846 4243 5902
rect 4299 5846 4309 5902
rect 2497 5778 4309 5846
rect 2497 5722 2507 5778
rect 2563 5722 2631 5778
rect 2687 5722 2755 5778
rect 2811 5722 2879 5778
rect 2935 5722 3003 5778
rect 3059 5722 3127 5778
rect 3183 5722 3251 5778
rect 3307 5722 3375 5778
rect 3431 5722 3499 5778
rect 3555 5722 3623 5778
rect 3679 5722 3747 5778
rect 3803 5722 3871 5778
rect 3927 5722 3995 5778
rect 4051 5722 4119 5778
rect 4175 5722 4243 5778
rect 4299 5722 4309 5778
rect 2497 5654 4309 5722
rect 2497 5598 2507 5654
rect 2563 5598 2631 5654
rect 2687 5598 2755 5654
rect 2811 5598 2879 5654
rect 2935 5598 3003 5654
rect 3059 5598 3127 5654
rect 3183 5598 3251 5654
rect 3307 5598 3375 5654
rect 3431 5598 3499 5654
rect 3555 5598 3623 5654
rect 3679 5598 3747 5654
rect 3803 5598 3871 5654
rect 3927 5598 3995 5654
rect 4051 5598 4119 5654
rect 4175 5598 4243 5654
rect 4299 5598 4309 5654
rect 2497 5530 4309 5598
rect 2497 5474 2507 5530
rect 2563 5474 2631 5530
rect 2687 5474 2755 5530
rect 2811 5474 2879 5530
rect 2935 5474 3003 5530
rect 3059 5474 3127 5530
rect 3183 5474 3251 5530
rect 3307 5474 3375 5530
rect 3431 5474 3499 5530
rect 3555 5474 3623 5530
rect 3679 5474 3747 5530
rect 3803 5474 3871 5530
rect 3927 5474 3995 5530
rect 4051 5474 4119 5530
rect 4175 5474 4243 5530
rect 4299 5474 4309 5530
rect 2497 5406 4309 5474
rect 2497 5350 2507 5406
rect 2563 5350 2631 5406
rect 2687 5350 2755 5406
rect 2811 5350 2879 5406
rect 2935 5350 3003 5406
rect 3059 5350 3127 5406
rect 3183 5350 3251 5406
rect 3307 5350 3375 5406
rect 3431 5350 3499 5406
rect 3555 5350 3623 5406
rect 3679 5350 3747 5406
rect 3803 5350 3871 5406
rect 3927 5350 3995 5406
rect 4051 5350 4119 5406
rect 4175 5350 4243 5406
rect 4299 5350 4309 5406
rect 2497 5282 4309 5350
rect 2497 5226 2507 5282
rect 2563 5226 2631 5282
rect 2687 5226 2755 5282
rect 2811 5226 2879 5282
rect 2935 5226 3003 5282
rect 3059 5226 3127 5282
rect 3183 5226 3251 5282
rect 3307 5226 3375 5282
rect 3431 5226 3499 5282
rect 3555 5226 3623 5282
rect 3679 5226 3747 5282
rect 3803 5226 3871 5282
rect 3927 5226 3995 5282
rect 4051 5226 4119 5282
rect 4175 5226 4243 5282
rect 4299 5226 4309 5282
rect 2497 5158 4309 5226
rect 2497 5102 2507 5158
rect 2563 5102 2631 5158
rect 2687 5102 2755 5158
rect 2811 5102 2879 5158
rect 2935 5102 3003 5158
rect 3059 5102 3127 5158
rect 3183 5102 3251 5158
rect 3307 5102 3375 5158
rect 3431 5102 3499 5158
rect 3555 5102 3623 5158
rect 3679 5102 3747 5158
rect 3803 5102 3871 5158
rect 3927 5102 3995 5158
rect 4051 5102 4119 5158
rect 4175 5102 4243 5158
rect 4299 5102 4309 5158
rect 2497 5034 4309 5102
rect 2497 4978 2507 5034
rect 2563 4978 2631 5034
rect 2687 4978 2755 5034
rect 2811 4978 2879 5034
rect 2935 4978 3003 5034
rect 3059 4978 3127 5034
rect 3183 4978 3251 5034
rect 3307 4978 3375 5034
rect 3431 4978 3499 5034
rect 3555 4978 3623 5034
rect 3679 4978 3747 5034
rect 3803 4978 3871 5034
rect 3927 4978 3995 5034
rect 4051 4978 4119 5034
rect 4175 4978 4243 5034
rect 4299 4978 4309 5034
rect 2497 4910 4309 4978
rect 2497 4854 2507 4910
rect 2563 4854 2631 4910
rect 2687 4854 2755 4910
rect 2811 4854 2879 4910
rect 2935 4854 3003 4910
rect 3059 4854 3127 4910
rect 3183 4854 3251 4910
rect 3307 4854 3375 4910
rect 3431 4854 3499 4910
rect 3555 4854 3623 4910
rect 3679 4854 3747 4910
rect 3803 4854 3871 4910
rect 3927 4854 3995 4910
rect 4051 4854 4119 4910
rect 4175 4854 4243 4910
rect 4299 4854 4309 4910
rect 2497 4786 4309 4854
rect 2497 4730 2507 4786
rect 2563 4730 2631 4786
rect 2687 4730 2755 4786
rect 2811 4730 2879 4786
rect 2935 4730 3003 4786
rect 3059 4730 3127 4786
rect 3183 4730 3251 4786
rect 3307 4730 3375 4786
rect 3431 4730 3499 4786
rect 3555 4730 3623 4786
rect 3679 4730 3747 4786
rect 3803 4730 3871 4786
rect 3927 4730 3995 4786
rect 4051 4730 4119 4786
rect 4175 4730 4243 4786
rect 4299 4730 4309 4786
rect 2497 4662 4309 4730
rect 2497 4606 2507 4662
rect 2563 4606 2631 4662
rect 2687 4606 2755 4662
rect 2811 4606 2879 4662
rect 2935 4606 3003 4662
rect 3059 4606 3127 4662
rect 3183 4606 3251 4662
rect 3307 4606 3375 4662
rect 3431 4606 3499 4662
rect 3555 4606 3623 4662
rect 3679 4606 3747 4662
rect 3803 4606 3871 4662
rect 3927 4606 3995 4662
rect 4051 4606 4119 4662
rect 4175 4606 4243 4662
rect 4299 4606 4309 4662
rect 2497 4538 4309 4606
rect 2497 4482 2507 4538
rect 2563 4482 2631 4538
rect 2687 4482 2755 4538
rect 2811 4482 2879 4538
rect 2935 4482 3003 4538
rect 3059 4482 3127 4538
rect 3183 4482 3251 4538
rect 3307 4482 3375 4538
rect 3431 4482 3499 4538
rect 3555 4482 3623 4538
rect 3679 4482 3747 4538
rect 3803 4482 3871 4538
rect 3927 4482 3995 4538
rect 4051 4482 4119 4538
rect 4175 4482 4243 4538
rect 4299 4482 4309 4538
rect 2497 4414 4309 4482
rect 2497 4358 2507 4414
rect 2563 4358 2631 4414
rect 2687 4358 2755 4414
rect 2811 4358 2879 4414
rect 2935 4358 3003 4414
rect 3059 4358 3127 4414
rect 3183 4358 3251 4414
rect 3307 4358 3375 4414
rect 3431 4358 3499 4414
rect 3555 4358 3623 4414
rect 3679 4358 3747 4414
rect 3803 4358 3871 4414
rect 3927 4358 3995 4414
rect 4051 4358 4119 4414
rect 4175 4358 4243 4414
rect 4299 4358 4309 4414
rect 2497 4290 4309 4358
rect 2497 4234 2507 4290
rect 2563 4234 2631 4290
rect 2687 4234 2755 4290
rect 2811 4234 2879 4290
rect 2935 4234 3003 4290
rect 3059 4234 3127 4290
rect 3183 4234 3251 4290
rect 3307 4234 3375 4290
rect 3431 4234 3499 4290
rect 3555 4234 3623 4290
rect 3679 4234 3747 4290
rect 3803 4234 3871 4290
rect 3927 4234 3995 4290
rect 4051 4234 4119 4290
rect 4175 4234 4243 4290
rect 4299 4234 4309 4290
rect 2497 4166 4309 4234
rect 2497 4110 2507 4166
rect 2563 4110 2631 4166
rect 2687 4110 2755 4166
rect 2811 4110 2879 4166
rect 2935 4110 3003 4166
rect 3059 4110 3127 4166
rect 3183 4110 3251 4166
rect 3307 4110 3375 4166
rect 3431 4110 3499 4166
rect 3555 4110 3623 4166
rect 3679 4110 3747 4166
rect 3803 4110 3871 4166
rect 3927 4110 3995 4166
rect 4051 4110 4119 4166
rect 4175 4110 4243 4166
rect 4299 4110 4309 4166
rect 2497 4042 4309 4110
rect 2497 3986 2507 4042
rect 2563 3986 2631 4042
rect 2687 3986 2755 4042
rect 2811 3986 2879 4042
rect 2935 3986 3003 4042
rect 3059 3986 3127 4042
rect 3183 3986 3251 4042
rect 3307 3986 3375 4042
rect 3431 3986 3499 4042
rect 3555 3986 3623 4042
rect 3679 3986 3747 4042
rect 3803 3986 3871 4042
rect 3927 3986 3995 4042
rect 4051 3986 4119 4042
rect 4175 3986 4243 4042
rect 4299 3986 4309 4042
rect 2497 3918 4309 3986
rect 2497 3862 2507 3918
rect 2563 3862 2631 3918
rect 2687 3862 2755 3918
rect 2811 3862 2879 3918
rect 2935 3862 3003 3918
rect 3059 3862 3127 3918
rect 3183 3862 3251 3918
rect 3307 3862 3375 3918
rect 3431 3862 3499 3918
rect 3555 3862 3623 3918
rect 3679 3862 3747 3918
rect 3803 3862 3871 3918
rect 3927 3862 3995 3918
rect 4051 3862 4119 3918
rect 4175 3862 4243 3918
rect 4299 3862 4309 3918
rect 2497 3794 4309 3862
rect 2497 3738 2507 3794
rect 2563 3738 2631 3794
rect 2687 3738 2755 3794
rect 2811 3738 2879 3794
rect 2935 3738 3003 3794
rect 3059 3738 3127 3794
rect 3183 3738 3251 3794
rect 3307 3738 3375 3794
rect 3431 3738 3499 3794
rect 3555 3738 3623 3794
rect 3679 3738 3747 3794
rect 3803 3738 3871 3794
rect 3927 3738 3995 3794
rect 4051 3738 4119 3794
rect 4175 3738 4243 3794
rect 4299 3738 4309 3794
rect 2497 3670 4309 3738
rect 2497 3614 2507 3670
rect 2563 3614 2631 3670
rect 2687 3614 2755 3670
rect 2811 3614 2879 3670
rect 2935 3614 3003 3670
rect 3059 3614 3127 3670
rect 3183 3614 3251 3670
rect 3307 3614 3375 3670
rect 3431 3614 3499 3670
rect 3555 3614 3623 3670
rect 3679 3614 3747 3670
rect 3803 3614 3871 3670
rect 3927 3614 3995 3670
rect 4051 3614 4119 3670
rect 4175 3614 4243 3670
rect 4299 3614 4309 3670
rect 2497 3546 4309 3614
rect 2497 3490 2507 3546
rect 2563 3490 2631 3546
rect 2687 3490 2755 3546
rect 2811 3490 2879 3546
rect 2935 3490 3003 3546
rect 3059 3490 3127 3546
rect 3183 3490 3251 3546
rect 3307 3490 3375 3546
rect 3431 3490 3499 3546
rect 3555 3490 3623 3546
rect 3679 3490 3747 3546
rect 3803 3490 3871 3546
rect 3927 3490 3995 3546
rect 4051 3490 4119 3546
rect 4175 3490 4243 3546
rect 4299 3490 4309 3546
rect 2497 3422 4309 3490
rect 2497 3366 2507 3422
rect 2563 3366 2631 3422
rect 2687 3366 2755 3422
rect 2811 3366 2879 3422
rect 2935 3366 3003 3422
rect 3059 3366 3127 3422
rect 3183 3366 3251 3422
rect 3307 3366 3375 3422
rect 3431 3366 3499 3422
rect 3555 3366 3623 3422
rect 3679 3366 3747 3422
rect 3803 3366 3871 3422
rect 3927 3366 3995 3422
rect 4051 3366 4119 3422
rect 4175 3366 4243 3422
rect 4299 3366 4309 3422
rect 2497 3298 4309 3366
rect 2497 3242 2507 3298
rect 2563 3242 2631 3298
rect 2687 3242 2755 3298
rect 2811 3242 2879 3298
rect 2935 3242 3003 3298
rect 3059 3242 3127 3298
rect 3183 3242 3251 3298
rect 3307 3242 3375 3298
rect 3431 3242 3499 3298
rect 3555 3242 3623 3298
rect 3679 3242 3747 3298
rect 3803 3242 3871 3298
rect 3927 3242 3995 3298
rect 4051 3242 4119 3298
rect 4175 3242 4243 3298
rect 4299 3242 4309 3298
rect 2497 3232 4309 3242
rect 6358 6150 7426 6160
rect 6358 6094 6368 6150
rect 6424 6094 6492 6150
rect 6548 6094 6616 6150
rect 6672 6094 6740 6150
rect 6796 6094 6864 6150
rect 6920 6094 6988 6150
rect 7044 6094 7112 6150
rect 7168 6094 7236 6150
rect 7292 6094 7360 6150
rect 7416 6094 7426 6150
rect 6358 6026 7426 6094
rect 6358 5970 6368 6026
rect 6424 5970 6492 6026
rect 6548 5970 6616 6026
rect 6672 5970 6740 6026
rect 6796 5970 6864 6026
rect 6920 5970 6988 6026
rect 7044 5970 7112 6026
rect 7168 5970 7236 6026
rect 7292 5970 7360 6026
rect 7416 5970 7426 6026
rect 6358 5902 7426 5970
rect 6358 5846 6368 5902
rect 6424 5846 6492 5902
rect 6548 5846 6616 5902
rect 6672 5846 6740 5902
rect 6796 5846 6864 5902
rect 6920 5846 6988 5902
rect 7044 5846 7112 5902
rect 7168 5846 7236 5902
rect 7292 5846 7360 5902
rect 7416 5846 7426 5902
rect 6358 5778 7426 5846
rect 6358 5722 6368 5778
rect 6424 5722 6492 5778
rect 6548 5722 6616 5778
rect 6672 5722 6740 5778
rect 6796 5722 6864 5778
rect 6920 5722 6988 5778
rect 7044 5722 7112 5778
rect 7168 5722 7236 5778
rect 7292 5722 7360 5778
rect 7416 5722 7426 5778
rect 6358 5654 7426 5722
rect 6358 5598 6368 5654
rect 6424 5598 6492 5654
rect 6548 5598 6616 5654
rect 6672 5598 6740 5654
rect 6796 5598 6864 5654
rect 6920 5598 6988 5654
rect 7044 5598 7112 5654
rect 7168 5598 7236 5654
rect 7292 5598 7360 5654
rect 7416 5598 7426 5654
rect 6358 5530 7426 5598
rect 6358 5474 6368 5530
rect 6424 5474 6492 5530
rect 6548 5474 6616 5530
rect 6672 5474 6740 5530
rect 6796 5474 6864 5530
rect 6920 5474 6988 5530
rect 7044 5474 7112 5530
rect 7168 5474 7236 5530
rect 7292 5474 7360 5530
rect 7416 5474 7426 5530
rect 6358 5406 7426 5474
rect 6358 5350 6368 5406
rect 6424 5350 6492 5406
rect 6548 5350 6616 5406
rect 6672 5350 6740 5406
rect 6796 5350 6864 5406
rect 6920 5350 6988 5406
rect 7044 5350 7112 5406
rect 7168 5350 7236 5406
rect 7292 5350 7360 5406
rect 7416 5350 7426 5406
rect 6358 5282 7426 5350
rect 6358 5226 6368 5282
rect 6424 5226 6492 5282
rect 6548 5226 6616 5282
rect 6672 5226 6740 5282
rect 6796 5226 6864 5282
rect 6920 5226 6988 5282
rect 7044 5226 7112 5282
rect 7168 5226 7236 5282
rect 7292 5226 7360 5282
rect 7416 5226 7426 5282
rect 6358 5158 7426 5226
rect 6358 5102 6368 5158
rect 6424 5102 6492 5158
rect 6548 5102 6616 5158
rect 6672 5102 6740 5158
rect 6796 5102 6864 5158
rect 6920 5102 6988 5158
rect 7044 5102 7112 5158
rect 7168 5102 7236 5158
rect 7292 5102 7360 5158
rect 7416 5102 7426 5158
rect 6358 5034 7426 5102
rect 6358 4978 6368 5034
rect 6424 4978 6492 5034
rect 6548 4978 6616 5034
rect 6672 4978 6740 5034
rect 6796 4978 6864 5034
rect 6920 4978 6988 5034
rect 7044 4978 7112 5034
rect 7168 4978 7236 5034
rect 7292 4978 7360 5034
rect 7416 4978 7426 5034
rect 6358 4910 7426 4978
rect 6358 4854 6368 4910
rect 6424 4854 6492 4910
rect 6548 4854 6616 4910
rect 6672 4854 6740 4910
rect 6796 4854 6864 4910
rect 6920 4854 6988 4910
rect 7044 4854 7112 4910
rect 7168 4854 7236 4910
rect 7292 4854 7360 4910
rect 7416 4854 7426 4910
rect 6358 4786 7426 4854
rect 6358 4730 6368 4786
rect 6424 4730 6492 4786
rect 6548 4730 6616 4786
rect 6672 4730 6740 4786
rect 6796 4730 6864 4786
rect 6920 4730 6988 4786
rect 7044 4730 7112 4786
rect 7168 4730 7236 4786
rect 7292 4730 7360 4786
rect 7416 4730 7426 4786
rect 6358 4662 7426 4730
rect 6358 4606 6368 4662
rect 6424 4606 6492 4662
rect 6548 4606 6616 4662
rect 6672 4606 6740 4662
rect 6796 4606 6864 4662
rect 6920 4606 6988 4662
rect 7044 4606 7112 4662
rect 7168 4606 7236 4662
rect 7292 4606 7360 4662
rect 7416 4606 7426 4662
rect 6358 4538 7426 4606
rect 6358 4482 6368 4538
rect 6424 4482 6492 4538
rect 6548 4482 6616 4538
rect 6672 4482 6740 4538
rect 6796 4482 6864 4538
rect 6920 4482 6988 4538
rect 7044 4482 7112 4538
rect 7168 4482 7236 4538
rect 7292 4482 7360 4538
rect 7416 4482 7426 4538
rect 6358 4414 7426 4482
rect 6358 4358 6368 4414
rect 6424 4358 6492 4414
rect 6548 4358 6616 4414
rect 6672 4358 6740 4414
rect 6796 4358 6864 4414
rect 6920 4358 6988 4414
rect 7044 4358 7112 4414
rect 7168 4358 7236 4414
rect 7292 4358 7360 4414
rect 7416 4358 7426 4414
rect 6358 4290 7426 4358
rect 6358 4234 6368 4290
rect 6424 4234 6492 4290
rect 6548 4234 6616 4290
rect 6672 4234 6740 4290
rect 6796 4234 6864 4290
rect 6920 4234 6988 4290
rect 7044 4234 7112 4290
rect 7168 4234 7236 4290
rect 7292 4234 7360 4290
rect 7416 4234 7426 4290
rect 6358 4166 7426 4234
rect 6358 4110 6368 4166
rect 6424 4110 6492 4166
rect 6548 4110 6616 4166
rect 6672 4110 6740 4166
rect 6796 4110 6864 4166
rect 6920 4110 6988 4166
rect 7044 4110 7112 4166
rect 7168 4110 7236 4166
rect 7292 4110 7360 4166
rect 7416 4110 7426 4166
rect 6358 4042 7426 4110
rect 6358 3986 6368 4042
rect 6424 3986 6492 4042
rect 6548 3986 6616 4042
rect 6672 3986 6740 4042
rect 6796 3986 6864 4042
rect 6920 3986 6988 4042
rect 7044 3986 7112 4042
rect 7168 3986 7236 4042
rect 7292 3986 7360 4042
rect 7416 3986 7426 4042
rect 6358 3918 7426 3986
rect 6358 3862 6368 3918
rect 6424 3862 6492 3918
rect 6548 3862 6616 3918
rect 6672 3862 6740 3918
rect 6796 3862 6864 3918
rect 6920 3862 6988 3918
rect 7044 3862 7112 3918
rect 7168 3862 7236 3918
rect 7292 3862 7360 3918
rect 7416 3862 7426 3918
rect 6358 3794 7426 3862
rect 6358 3738 6368 3794
rect 6424 3738 6492 3794
rect 6548 3738 6616 3794
rect 6672 3738 6740 3794
rect 6796 3738 6864 3794
rect 6920 3738 6988 3794
rect 7044 3738 7112 3794
rect 7168 3738 7236 3794
rect 7292 3738 7360 3794
rect 7416 3738 7426 3794
rect 6358 3670 7426 3738
rect 6358 3614 6368 3670
rect 6424 3614 6492 3670
rect 6548 3614 6616 3670
rect 6672 3614 6740 3670
rect 6796 3614 6864 3670
rect 6920 3614 6988 3670
rect 7044 3614 7112 3670
rect 7168 3614 7236 3670
rect 7292 3614 7360 3670
rect 7416 3614 7426 3670
rect 6358 3546 7426 3614
rect 6358 3490 6368 3546
rect 6424 3490 6492 3546
rect 6548 3490 6616 3546
rect 6672 3490 6740 3546
rect 6796 3490 6864 3546
rect 6920 3490 6988 3546
rect 7044 3490 7112 3546
rect 7168 3490 7236 3546
rect 7292 3490 7360 3546
rect 7416 3490 7426 3546
rect 6358 3422 7426 3490
rect 6358 3366 6368 3422
rect 6424 3366 6492 3422
rect 6548 3366 6616 3422
rect 6672 3366 6740 3422
rect 6796 3366 6864 3422
rect 6920 3366 6988 3422
rect 7044 3366 7112 3422
rect 7168 3366 7236 3422
rect 7292 3366 7360 3422
rect 7416 3366 7426 3422
rect 6358 3298 7426 3366
rect 6358 3242 6368 3298
rect 6424 3242 6492 3298
rect 6548 3242 6616 3298
rect 6672 3242 6740 3298
rect 6796 3242 6864 3298
rect 6920 3242 6988 3298
rect 7044 3242 7112 3298
rect 7168 3242 7236 3298
rect 7292 3242 7360 3298
rect 7416 3242 7426 3298
rect 6358 3232 7426 3242
rect 8741 6150 10553 6160
rect 8741 6094 8751 6150
rect 8807 6094 8875 6150
rect 8931 6094 8999 6150
rect 9055 6094 9123 6150
rect 9179 6094 9247 6150
rect 9303 6094 9371 6150
rect 9427 6094 9495 6150
rect 9551 6094 9619 6150
rect 9675 6094 9743 6150
rect 9799 6094 9867 6150
rect 9923 6094 9991 6150
rect 10047 6094 10115 6150
rect 10171 6094 10239 6150
rect 10295 6094 10363 6150
rect 10419 6094 10487 6150
rect 10543 6094 10553 6150
rect 8741 6026 10553 6094
rect 8741 5970 8751 6026
rect 8807 5970 8875 6026
rect 8931 5970 8999 6026
rect 9055 5970 9123 6026
rect 9179 5970 9247 6026
rect 9303 5970 9371 6026
rect 9427 5970 9495 6026
rect 9551 5970 9619 6026
rect 9675 5970 9743 6026
rect 9799 5970 9867 6026
rect 9923 5970 9991 6026
rect 10047 5970 10115 6026
rect 10171 5970 10239 6026
rect 10295 5970 10363 6026
rect 10419 5970 10487 6026
rect 10543 5970 10553 6026
rect 8741 5902 10553 5970
rect 8741 5846 8751 5902
rect 8807 5846 8875 5902
rect 8931 5846 8999 5902
rect 9055 5846 9123 5902
rect 9179 5846 9247 5902
rect 9303 5846 9371 5902
rect 9427 5846 9495 5902
rect 9551 5846 9619 5902
rect 9675 5846 9743 5902
rect 9799 5846 9867 5902
rect 9923 5846 9991 5902
rect 10047 5846 10115 5902
rect 10171 5846 10239 5902
rect 10295 5846 10363 5902
rect 10419 5846 10487 5902
rect 10543 5846 10553 5902
rect 8741 5778 10553 5846
rect 8741 5722 8751 5778
rect 8807 5722 8875 5778
rect 8931 5722 8999 5778
rect 9055 5722 9123 5778
rect 9179 5722 9247 5778
rect 9303 5722 9371 5778
rect 9427 5722 9495 5778
rect 9551 5722 9619 5778
rect 9675 5722 9743 5778
rect 9799 5722 9867 5778
rect 9923 5722 9991 5778
rect 10047 5722 10115 5778
rect 10171 5722 10239 5778
rect 10295 5722 10363 5778
rect 10419 5722 10487 5778
rect 10543 5722 10553 5778
rect 8741 5654 10553 5722
rect 8741 5598 8751 5654
rect 8807 5598 8875 5654
rect 8931 5598 8999 5654
rect 9055 5598 9123 5654
rect 9179 5598 9247 5654
rect 9303 5598 9371 5654
rect 9427 5598 9495 5654
rect 9551 5598 9619 5654
rect 9675 5598 9743 5654
rect 9799 5598 9867 5654
rect 9923 5598 9991 5654
rect 10047 5598 10115 5654
rect 10171 5598 10239 5654
rect 10295 5598 10363 5654
rect 10419 5598 10487 5654
rect 10543 5598 10553 5654
rect 8741 5530 10553 5598
rect 8741 5474 8751 5530
rect 8807 5474 8875 5530
rect 8931 5474 8999 5530
rect 9055 5474 9123 5530
rect 9179 5474 9247 5530
rect 9303 5474 9371 5530
rect 9427 5474 9495 5530
rect 9551 5474 9619 5530
rect 9675 5474 9743 5530
rect 9799 5474 9867 5530
rect 9923 5474 9991 5530
rect 10047 5474 10115 5530
rect 10171 5474 10239 5530
rect 10295 5474 10363 5530
rect 10419 5474 10487 5530
rect 10543 5474 10553 5530
rect 8741 5406 10553 5474
rect 8741 5350 8751 5406
rect 8807 5350 8875 5406
rect 8931 5350 8999 5406
rect 9055 5350 9123 5406
rect 9179 5350 9247 5406
rect 9303 5350 9371 5406
rect 9427 5350 9495 5406
rect 9551 5350 9619 5406
rect 9675 5350 9743 5406
rect 9799 5350 9867 5406
rect 9923 5350 9991 5406
rect 10047 5350 10115 5406
rect 10171 5350 10239 5406
rect 10295 5350 10363 5406
rect 10419 5350 10487 5406
rect 10543 5350 10553 5406
rect 8741 5282 10553 5350
rect 8741 5226 8751 5282
rect 8807 5226 8875 5282
rect 8931 5226 8999 5282
rect 9055 5226 9123 5282
rect 9179 5226 9247 5282
rect 9303 5226 9371 5282
rect 9427 5226 9495 5282
rect 9551 5226 9619 5282
rect 9675 5226 9743 5282
rect 9799 5226 9867 5282
rect 9923 5226 9991 5282
rect 10047 5226 10115 5282
rect 10171 5226 10239 5282
rect 10295 5226 10363 5282
rect 10419 5226 10487 5282
rect 10543 5226 10553 5282
rect 8741 5158 10553 5226
rect 8741 5102 8751 5158
rect 8807 5102 8875 5158
rect 8931 5102 8999 5158
rect 9055 5102 9123 5158
rect 9179 5102 9247 5158
rect 9303 5102 9371 5158
rect 9427 5102 9495 5158
rect 9551 5102 9619 5158
rect 9675 5102 9743 5158
rect 9799 5102 9867 5158
rect 9923 5102 9991 5158
rect 10047 5102 10115 5158
rect 10171 5102 10239 5158
rect 10295 5102 10363 5158
rect 10419 5102 10487 5158
rect 10543 5102 10553 5158
rect 8741 5034 10553 5102
rect 8741 4978 8751 5034
rect 8807 4978 8875 5034
rect 8931 4978 8999 5034
rect 9055 4978 9123 5034
rect 9179 4978 9247 5034
rect 9303 4978 9371 5034
rect 9427 4978 9495 5034
rect 9551 4978 9619 5034
rect 9675 4978 9743 5034
rect 9799 4978 9867 5034
rect 9923 4978 9991 5034
rect 10047 4978 10115 5034
rect 10171 4978 10239 5034
rect 10295 4978 10363 5034
rect 10419 4978 10487 5034
rect 10543 4978 10553 5034
rect 8741 4910 10553 4978
rect 8741 4854 8751 4910
rect 8807 4854 8875 4910
rect 8931 4854 8999 4910
rect 9055 4854 9123 4910
rect 9179 4854 9247 4910
rect 9303 4854 9371 4910
rect 9427 4854 9495 4910
rect 9551 4854 9619 4910
rect 9675 4854 9743 4910
rect 9799 4854 9867 4910
rect 9923 4854 9991 4910
rect 10047 4854 10115 4910
rect 10171 4854 10239 4910
rect 10295 4854 10363 4910
rect 10419 4854 10487 4910
rect 10543 4854 10553 4910
rect 8741 4786 10553 4854
rect 8741 4730 8751 4786
rect 8807 4730 8875 4786
rect 8931 4730 8999 4786
rect 9055 4730 9123 4786
rect 9179 4730 9247 4786
rect 9303 4730 9371 4786
rect 9427 4730 9495 4786
rect 9551 4730 9619 4786
rect 9675 4730 9743 4786
rect 9799 4730 9867 4786
rect 9923 4730 9991 4786
rect 10047 4730 10115 4786
rect 10171 4730 10239 4786
rect 10295 4730 10363 4786
rect 10419 4730 10487 4786
rect 10543 4730 10553 4786
rect 8741 4662 10553 4730
rect 8741 4606 8751 4662
rect 8807 4606 8875 4662
rect 8931 4606 8999 4662
rect 9055 4606 9123 4662
rect 9179 4606 9247 4662
rect 9303 4606 9371 4662
rect 9427 4606 9495 4662
rect 9551 4606 9619 4662
rect 9675 4606 9743 4662
rect 9799 4606 9867 4662
rect 9923 4606 9991 4662
rect 10047 4606 10115 4662
rect 10171 4606 10239 4662
rect 10295 4606 10363 4662
rect 10419 4606 10487 4662
rect 10543 4606 10553 4662
rect 8741 4538 10553 4606
rect 8741 4482 8751 4538
rect 8807 4482 8875 4538
rect 8931 4482 8999 4538
rect 9055 4482 9123 4538
rect 9179 4482 9247 4538
rect 9303 4482 9371 4538
rect 9427 4482 9495 4538
rect 9551 4482 9619 4538
rect 9675 4482 9743 4538
rect 9799 4482 9867 4538
rect 9923 4482 9991 4538
rect 10047 4482 10115 4538
rect 10171 4482 10239 4538
rect 10295 4482 10363 4538
rect 10419 4482 10487 4538
rect 10543 4482 10553 4538
rect 8741 4414 10553 4482
rect 8741 4358 8751 4414
rect 8807 4358 8875 4414
rect 8931 4358 8999 4414
rect 9055 4358 9123 4414
rect 9179 4358 9247 4414
rect 9303 4358 9371 4414
rect 9427 4358 9495 4414
rect 9551 4358 9619 4414
rect 9675 4358 9743 4414
rect 9799 4358 9867 4414
rect 9923 4358 9991 4414
rect 10047 4358 10115 4414
rect 10171 4358 10239 4414
rect 10295 4358 10363 4414
rect 10419 4358 10487 4414
rect 10543 4358 10553 4414
rect 8741 4290 10553 4358
rect 8741 4234 8751 4290
rect 8807 4234 8875 4290
rect 8931 4234 8999 4290
rect 9055 4234 9123 4290
rect 9179 4234 9247 4290
rect 9303 4234 9371 4290
rect 9427 4234 9495 4290
rect 9551 4234 9619 4290
rect 9675 4234 9743 4290
rect 9799 4234 9867 4290
rect 9923 4234 9991 4290
rect 10047 4234 10115 4290
rect 10171 4234 10239 4290
rect 10295 4234 10363 4290
rect 10419 4234 10487 4290
rect 10543 4234 10553 4290
rect 8741 4166 10553 4234
rect 8741 4110 8751 4166
rect 8807 4110 8875 4166
rect 8931 4110 8999 4166
rect 9055 4110 9123 4166
rect 9179 4110 9247 4166
rect 9303 4110 9371 4166
rect 9427 4110 9495 4166
rect 9551 4110 9619 4166
rect 9675 4110 9743 4166
rect 9799 4110 9867 4166
rect 9923 4110 9991 4166
rect 10047 4110 10115 4166
rect 10171 4110 10239 4166
rect 10295 4110 10363 4166
rect 10419 4110 10487 4166
rect 10543 4110 10553 4166
rect 8741 4042 10553 4110
rect 8741 3986 8751 4042
rect 8807 3986 8875 4042
rect 8931 3986 8999 4042
rect 9055 3986 9123 4042
rect 9179 3986 9247 4042
rect 9303 3986 9371 4042
rect 9427 3986 9495 4042
rect 9551 3986 9619 4042
rect 9675 3986 9743 4042
rect 9799 3986 9867 4042
rect 9923 3986 9991 4042
rect 10047 3986 10115 4042
rect 10171 3986 10239 4042
rect 10295 3986 10363 4042
rect 10419 3986 10487 4042
rect 10543 3986 10553 4042
rect 8741 3918 10553 3986
rect 8741 3862 8751 3918
rect 8807 3862 8875 3918
rect 8931 3862 8999 3918
rect 9055 3862 9123 3918
rect 9179 3862 9247 3918
rect 9303 3862 9371 3918
rect 9427 3862 9495 3918
rect 9551 3862 9619 3918
rect 9675 3862 9743 3918
rect 9799 3862 9867 3918
rect 9923 3862 9991 3918
rect 10047 3862 10115 3918
rect 10171 3862 10239 3918
rect 10295 3862 10363 3918
rect 10419 3862 10487 3918
rect 10543 3862 10553 3918
rect 8741 3794 10553 3862
rect 8741 3738 8751 3794
rect 8807 3738 8875 3794
rect 8931 3738 8999 3794
rect 9055 3738 9123 3794
rect 9179 3738 9247 3794
rect 9303 3738 9371 3794
rect 9427 3738 9495 3794
rect 9551 3738 9619 3794
rect 9675 3738 9743 3794
rect 9799 3738 9867 3794
rect 9923 3738 9991 3794
rect 10047 3738 10115 3794
rect 10171 3738 10239 3794
rect 10295 3738 10363 3794
rect 10419 3738 10487 3794
rect 10543 3738 10553 3794
rect 8741 3670 10553 3738
rect 8741 3614 8751 3670
rect 8807 3614 8875 3670
rect 8931 3614 8999 3670
rect 9055 3614 9123 3670
rect 9179 3614 9247 3670
rect 9303 3614 9371 3670
rect 9427 3614 9495 3670
rect 9551 3614 9619 3670
rect 9675 3614 9743 3670
rect 9799 3614 9867 3670
rect 9923 3614 9991 3670
rect 10047 3614 10115 3670
rect 10171 3614 10239 3670
rect 10295 3614 10363 3670
rect 10419 3614 10487 3670
rect 10543 3614 10553 3670
rect 8741 3546 10553 3614
rect 8741 3490 8751 3546
rect 8807 3490 8875 3546
rect 8931 3490 8999 3546
rect 9055 3490 9123 3546
rect 9179 3490 9247 3546
rect 9303 3490 9371 3546
rect 9427 3490 9495 3546
rect 9551 3490 9619 3546
rect 9675 3490 9743 3546
rect 9799 3490 9867 3546
rect 9923 3490 9991 3546
rect 10047 3490 10115 3546
rect 10171 3490 10239 3546
rect 10295 3490 10363 3546
rect 10419 3490 10487 3546
rect 10543 3490 10553 3546
rect 8741 3422 10553 3490
rect 8741 3366 8751 3422
rect 8807 3366 8875 3422
rect 8931 3366 8999 3422
rect 9055 3366 9123 3422
rect 9179 3366 9247 3422
rect 9303 3366 9371 3422
rect 9427 3366 9495 3422
rect 9551 3366 9619 3422
rect 9675 3366 9743 3422
rect 9799 3366 9867 3422
rect 9923 3366 9991 3422
rect 10047 3366 10115 3422
rect 10171 3366 10239 3422
rect 10295 3366 10363 3422
rect 10419 3366 10487 3422
rect 10543 3366 10553 3422
rect 8741 3298 10553 3366
rect 8741 3242 8751 3298
rect 8807 3242 8875 3298
rect 8931 3242 8999 3298
rect 9055 3242 9123 3298
rect 9179 3242 9247 3298
rect 9303 3242 9371 3298
rect 9427 3242 9495 3298
rect 9551 3242 9619 3298
rect 9675 3242 9743 3298
rect 9799 3242 9867 3298
rect 9923 3242 9991 3298
rect 10047 3242 10115 3298
rect 10171 3242 10239 3298
rect 10295 3242 10363 3298
rect 10419 3242 10487 3298
rect 10543 3242 10553 3298
rect 8741 3232 10553 3242
rect 12842 6150 13910 6160
rect 12842 6094 12852 6150
rect 12908 6094 12976 6150
rect 13032 6094 13100 6150
rect 13156 6094 13224 6150
rect 13280 6094 13348 6150
rect 13404 6094 13472 6150
rect 13528 6094 13596 6150
rect 13652 6094 13720 6150
rect 13776 6094 13844 6150
rect 13900 6094 13910 6150
rect 12842 6026 13910 6094
rect 12842 5970 12852 6026
rect 12908 5970 12976 6026
rect 13032 5970 13100 6026
rect 13156 5970 13224 6026
rect 13280 5970 13348 6026
rect 13404 5970 13472 6026
rect 13528 5970 13596 6026
rect 13652 5970 13720 6026
rect 13776 5970 13844 6026
rect 13900 5970 13910 6026
rect 12842 5902 13910 5970
rect 12842 5846 12852 5902
rect 12908 5846 12976 5902
rect 13032 5846 13100 5902
rect 13156 5846 13224 5902
rect 13280 5846 13348 5902
rect 13404 5846 13472 5902
rect 13528 5846 13596 5902
rect 13652 5846 13720 5902
rect 13776 5846 13844 5902
rect 13900 5846 13910 5902
rect 12842 5778 13910 5846
rect 12842 5722 12852 5778
rect 12908 5722 12976 5778
rect 13032 5722 13100 5778
rect 13156 5722 13224 5778
rect 13280 5722 13348 5778
rect 13404 5722 13472 5778
rect 13528 5722 13596 5778
rect 13652 5722 13720 5778
rect 13776 5722 13844 5778
rect 13900 5722 13910 5778
rect 12842 5654 13910 5722
rect 12842 5598 12852 5654
rect 12908 5598 12976 5654
rect 13032 5598 13100 5654
rect 13156 5598 13224 5654
rect 13280 5598 13348 5654
rect 13404 5598 13472 5654
rect 13528 5598 13596 5654
rect 13652 5598 13720 5654
rect 13776 5598 13844 5654
rect 13900 5598 13910 5654
rect 12842 5530 13910 5598
rect 12842 5474 12852 5530
rect 12908 5474 12976 5530
rect 13032 5474 13100 5530
rect 13156 5474 13224 5530
rect 13280 5474 13348 5530
rect 13404 5474 13472 5530
rect 13528 5474 13596 5530
rect 13652 5474 13720 5530
rect 13776 5474 13844 5530
rect 13900 5474 13910 5530
rect 12842 5406 13910 5474
rect 12842 5350 12852 5406
rect 12908 5350 12976 5406
rect 13032 5350 13100 5406
rect 13156 5350 13224 5406
rect 13280 5350 13348 5406
rect 13404 5350 13472 5406
rect 13528 5350 13596 5406
rect 13652 5350 13720 5406
rect 13776 5350 13844 5406
rect 13900 5350 13910 5406
rect 12842 5282 13910 5350
rect 12842 5226 12852 5282
rect 12908 5226 12976 5282
rect 13032 5226 13100 5282
rect 13156 5226 13224 5282
rect 13280 5226 13348 5282
rect 13404 5226 13472 5282
rect 13528 5226 13596 5282
rect 13652 5226 13720 5282
rect 13776 5226 13844 5282
rect 13900 5226 13910 5282
rect 12842 5158 13910 5226
rect 12842 5102 12852 5158
rect 12908 5102 12976 5158
rect 13032 5102 13100 5158
rect 13156 5102 13224 5158
rect 13280 5102 13348 5158
rect 13404 5102 13472 5158
rect 13528 5102 13596 5158
rect 13652 5102 13720 5158
rect 13776 5102 13844 5158
rect 13900 5102 13910 5158
rect 12842 5034 13910 5102
rect 12842 4978 12852 5034
rect 12908 4978 12976 5034
rect 13032 4978 13100 5034
rect 13156 4978 13224 5034
rect 13280 4978 13348 5034
rect 13404 4978 13472 5034
rect 13528 4978 13596 5034
rect 13652 4978 13720 5034
rect 13776 4978 13844 5034
rect 13900 4978 13910 5034
rect 12842 4910 13910 4978
rect 12842 4854 12852 4910
rect 12908 4854 12976 4910
rect 13032 4854 13100 4910
rect 13156 4854 13224 4910
rect 13280 4854 13348 4910
rect 13404 4854 13472 4910
rect 13528 4854 13596 4910
rect 13652 4854 13720 4910
rect 13776 4854 13844 4910
rect 13900 4854 13910 4910
rect 12842 4786 13910 4854
rect 12842 4730 12852 4786
rect 12908 4730 12976 4786
rect 13032 4730 13100 4786
rect 13156 4730 13224 4786
rect 13280 4730 13348 4786
rect 13404 4730 13472 4786
rect 13528 4730 13596 4786
rect 13652 4730 13720 4786
rect 13776 4730 13844 4786
rect 13900 4730 13910 4786
rect 12842 4662 13910 4730
rect 12842 4606 12852 4662
rect 12908 4606 12976 4662
rect 13032 4606 13100 4662
rect 13156 4606 13224 4662
rect 13280 4606 13348 4662
rect 13404 4606 13472 4662
rect 13528 4606 13596 4662
rect 13652 4606 13720 4662
rect 13776 4606 13844 4662
rect 13900 4606 13910 4662
rect 12842 4538 13910 4606
rect 12842 4482 12852 4538
rect 12908 4482 12976 4538
rect 13032 4482 13100 4538
rect 13156 4482 13224 4538
rect 13280 4482 13348 4538
rect 13404 4482 13472 4538
rect 13528 4482 13596 4538
rect 13652 4482 13720 4538
rect 13776 4482 13844 4538
rect 13900 4482 13910 4538
rect 12842 4414 13910 4482
rect 12842 4358 12852 4414
rect 12908 4358 12976 4414
rect 13032 4358 13100 4414
rect 13156 4358 13224 4414
rect 13280 4358 13348 4414
rect 13404 4358 13472 4414
rect 13528 4358 13596 4414
rect 13652 4358 13720 4414
rect 13776 4358 13844 4414
rect 13900 4358 13910 4414
rect 12842 4290 13910 4358
rect 12842 4234 12852 4290
rect 12908 4234 12976 4290
rect 13032 4234 13100 4290
rect 13156 4234 13224 4290
rect 13280 4234 13348 4290
rect 13404 4234 13472 4290
rect 13528 4234 13596 4290
rect 13652 4234 13720 4290
rect 13776 4234 13844 4290
rect 13900 4234 13910 4290
rect 12842 4166 13910 4234
rect 12842 4110 12852 4166
rect 12908 4110 12976 4166
rect 13032 4110 13100 4166
rect 13156 4110 13224 4166
rect 13280 4110 13348 4166
rect 13404 4110 13472 4166
rect 13528 4110 13596 4166
rect 13652 4110 13720 4166
rect 13776 4110 13844 4166
rect 13900 4110 13910 4166
rect 12842 4042 13910 4110
rect 12842 3986 12852 4042
rect 12908 3986 12976 4042
rect 13032 3986 13100 4042
rect 13156 3986 13224 4042
rect 13280 3986 13348 4042
rect 13404 3986 13472 4042
rect 13528 3986 13596 4042
rect 13652 3986 13720 4042
rect 13776 3986 13844 4042
rect 13900 3986 13910 4042
rect 12842 3918 13910 3986
rect 12842 3862 12852 3918
rect 12908 3862 12976 3918
rect 13032 3862 13100 3918
rect 13156 3862 13224 3918
rect 13280 3862 13348 3918
rect 13404 3862 13472 3918
rect 13528 3862 13596 3918
rect 13652 3862 13720 3918
rect 13776 3862 13844 3918
rect 13900 3862 13910 3918
rect 12842 3794 13910 3862
rect 12842 3738 12852 3794
rect 12908 3738 12976 3794
rect 13032 3738 13100 3794
rect 13156 3738 13224 3794
rect 13280 3738 13348 3794
rect 13404 3738 13472 3794
rect 13528 3738 13596 3794
rect 13652 3738 13720 3794
rect 13776 3738 13844 3794
rect 13900 3738 13910 3794
rect 12842 3670 13910 3738
rect 12842 3614 12852 3670
rect 12908 3614 12976 3670
rect 13032 3614 13100 3670
rect 13156 3614 13224 3670
rect 13280 3614 13348 3670
rect 13404 3614 13472 3670
rect 13528 3614 13596 3670
rect 13652 3614 13720 3670
rect 13776 3614 13844 3670
rect 13900 3614 13910 3670
rect 12842 3546 13910 3614
rect 12842 3490 12852 3546
rect 12908 3490 12976 3546
rect 13032 3490 13100 3546
rect 13156 3490 13224 3546
rect 13280 3490 13348 3546
rect 13404 3490 13472 3546
rect 13528 3490 13596 3546
rect 13652 3490 13720 3546
rect 13776 3490 13844 3546
rect 13900 3490 13910 3546
rect 12842 3422 13910 3490
rect 12842 3366 12852 3422
rect 12908 3366 12976 3422
rect 13032 3366 13100 3422
rect 13156 3366 13224 3422
rect 13280 3366 13348 3422
rect 13404 3366 13472 3422
rect 13528 3366 13596 3422
rect 13652 3366 13720 3422
rect 13776 3366 13844 3422
rect 13900 3366 13910 3422
rect 12842 3298 13910 3366
rect 12842 3242 12852 3298
rect 12908 3242 12976 3298
rect 13032 3242 13100 3298
rect 13156 3242 13224 3298
rect 13280 3242 13348 3298
rect 13404 3242 13472 3298
rect 13528 3242 13596 3298
rect 13652 3242 13720 3298
rect 13776 3242 13844 3298
rect 13900 3242 13910 3298
rect 12842 3232 13910 3242
rect 2497 2950 4309 2960
rect 2497 2894 2507 2950
rect 2563 2894 2631 2950
rect 2687 2894 2755 2950
rect 2811 2894 2879 2950
rect 2935 2894 3003 2950
rect 3059 2894 3127 2950
rect 3183 2894 3251 2950
rect 3307 2894 3375 2950
rect 3431 2894 3499 2950
rect 3555 2894 3623 2950
rect 3679 2894 3747 2950
rect 3803 2894 3871 2950
rect 3927 2894 3995 2950
rect 4051 2894 4119 2950
rect 4175 2894 4243 2950
rect 4299 2894 4309 2950
rect 2497 2826 4309 2894
rect 2497 2770 2507 2826
rect 2563 2770 2631 2826
rect 2687 2770 2755 2826
rect 2811 2770 2879 2826
rect 2935 2770 3003 2826
rect 3059 2770 3127 2826
rect 3183 2770 3251 2826
rect 3307 2770 3375 2826
rect 3431 2770 3499 2826
rect 3555 2770 3623 2826
rect 3679 2770 3747 2826
rect 3803 2770 3871 2826
rect 3927 2770 3995 2826
rect 4051 2770 4119 2826
rect 4175 2770 4243 2826
rect 4299 2770 4309 2826
rect 2497 2702 4309 2770
rect 2497 2646 2507 2702
rect 2563 2646 2631 2702
rect 2687 2646 2755 2702
rect 2811 2646 2879 2702
rect 2935 2646 3003 2702
rect 3059 2646 3127 2702
rect 3183 2646 3251 2702
rect 3307 2646 3375 2702
rect 3431 2646 3499 2702
rect 3555 2646 3623 2702
rect 3679 2646 3747 2702
rect 3803 2646 3871 2702
rect 3927 2646 3995 2702
rect 4051 2646 4119 2702
rect 4175 2646 4243 2702
rect 4299 2646 4309 2702
rect 2497 2578 4309 2646
rect 2497 2522 2507 2578
rect 2563 2522 2631 2578
rect 2687 2522 2755 2578
rect 2811 2522 2879 2578
rect 2935 2522 3003 2578
rect 3059 2522 3127 2578
rect 3183 2522 3251 2578
rect 3307 2522 3375 2578
rect 3431 2522 3499 2578
rect 3555 2522 3623 2578
rect 3679 2522 3747 2578
rect 3803 2522 3871 2578
rect 3927 2522 3995 2578
rect 4051 2522 4119 2578
rect 4175 2522 4243 2578
rect 4299 2522 4309 2578
rect 2497 2454 4309 2522
rect 2497 2398 2507 2454
rect 2563 2398 2631 2454
rect 2687 2398 2755 2454
rect 2811 2398 2879 2454
rect 2935 2398 3003 2454
rect 3059 2398 3127 2454
rect 3183 2398 3251 2454
rect 3307 2398 3375 2454
rect 3431 2398 3499 2454
rect 3555 2398 3623 2454
rect 3679 2398 3747 2454
rect 3803 2398 3871 2454
rect 3927 2398 3995 2454
rect 4051 2398 4119 2454
rect 4175 2398 4243 2454
rect 4299 2398 4309 2454
rect 2497 2330 4309 2398
rect 2497 2274 2507 2330
rect 2563 2274 2631 2330
rect 2687 2274 2755 2330
rect 2811 2274 2879 2330
rect 2935 2274 3003 2330
rect 3059 2274 3127 2330
rect 3183 2274 3251 2330
rect 3307 2274 3375 2330
rect 3431 2274 3499 2330
rect 3555 2274 3623 2330
rect 3679 2274 3747 2330
rect 3803 2274 3871 2330
rect 3927 2274 3995 2330
rect 4051 2274 4119 2330
rect 4175 2274 4243 2330
rect 4299 2274 4309 2330
rect 2497 2206 4309 2274
rect 2497 2150 2507 2206
rect 2563 2150 2631 2206
rect 2687 2150 2755 2206
rect 2811 2150 2879 2206
rect 2935 2150 3003 2206
rect 3059 2150 3127 2206
rect 3183 2150 3251 2206
rect 3307 2150 3375 2206
rect 3431 2150 3499 2206
rect 3555 2150 3623 2206
rect 3679 2150 3747 2206
rect 3803 2150 3871 2206
rect 3927 2150 3995 2206
rect 4051 2150 4119 2206
rect 4175 2150 4243 2206
rect 4299 2150 4309 2206
rect 2497 2082 4309 2150
rect 2497 2026 2507 2082
rect 2563 2026 2631 2082
rect 2687 2026 2755 2082
rect 2811 2026 2879 2082
rect 2935 2026 3003 2082
rect 3059 2026 3127 2082
rect 3183 2026 3251 2082
rect 3307 2026 3375 2082
rect 3431 2026 3499 2082
rect 3555 2026 3623 2082
rect 3679 2026 3747 2082
rect 3803 2026 3871 2082
rect 3927 2026 3995 2082
rect 4051 2026 4119 2082
rect 4175 2026 4243 2082
rect 4299 2026 4309 2082
rect 2497 1958 4309 2026
rect 2497 1902 2507 1958
rect 2563 1902 2631 1958
rect 2687 1902 2755 1958
rect 2811 1902 2879 1958
rect 2935 1902 3003 1958
rect 3059 1902 3127 1958
rect 3183 1902 3251 1958
rect 3307 1902 3375 1958
rect 3431 1902 3499 1958
rect 3555 1902 3623 1958
rect 3679 1902 3747 1958
rect 3803 1902 3871 1958
rect 3927 1902 3995 1958
rect 4051 1902 4119 1958
rect 4175 1902 4243 1958
rect 4299 1902 4309 1958
rect 2497 1834 4309 1902
rect 2497 1778 2507 1834
rect 2563 1778 2631 1834
rect 2687 1778 2755 1834
rect 2811 1778 2879 1834
rect 2935 1778 3003 1834
rect 3059 1778 3127 1834
rect 3183 1778 3251 1834
rect 3307 1778 3375 1834
rect 3431 1778 3499 1834
rect 3555 1778 3623 1834
rect 3679 1778 3747 1834
rect 3803 1778 3871 1834
rect 3927 1778 3995 1834
rect 4051 1778 4119 1834
rect 4175 1778 4243 1834
rect 4299 1778 4309 1834
rect 2497 1710 4309 1778
rect 2497 1654 2507 1710
rect 2563 1654 2631 1710
rect 2687 1654 2755 1710
rect 2811 1654 2879 1710
rect 2935 1654 3003 1710
rect 3059 1654 3127 1710
rect 3183 1654 3251 1710
rect 3307 1654 3375 1710
rect 3431 1654 3499 1710
rect 3555 1654 3623 1710
rect 3679 1654 3747 1710
rect 3803 1654 3871 1710
rect 3927 1654 3995 1710
rect 4051 1654 4119 1710
rect 4175 1654 4243 1710
rect 4299 1654 4309 1710
rect 2497 1586 4309 1654
rect 2497 1530 2507 1586
rect 2563 1530 2631 1586
rect 2687 1530 2755 1586
rect 2811 1530 2879 1586
rect 2935 1530 3003 1586
rect 3059 1530 3127 1586
rect 3183 1530 3251 1586
rect 3307 1530 3375 1586
rect 3431 1530 3499 1586
rect 3555 1530 3623 1586
rect 3679 1530 3747 1586
rect 3803 1530 3871 1586
rect 3927 1530 3995 1586
rect 4051 1530 4119 1586
rect 4175 1530 4243 1586
rect 4299 1530 4309 1586
rect 2497 1462 4309 1530
rect 2497 1406 2507 1462
rect 2563 1406 2631 1462
rect 2687 1406 2755 1462
rect 2811 1406 2879 1462
rect 2935 1406 3003 1462
rect 3059 1406 3127 1462
rect 3183 1406 3251 1462
rect 3307 1406 3375 1462
rect 3431 1406 3499 1462
rect 3555 1406 3623 1462
rect 3679 1406 3747 1462
rect 3803 1406 3871 1462
rect 3927 1406 3995 1462
rect 4051 1406 4119 1462
rect 4175 1406 4243 1462
rect 4299 1406 4309 1462
rect 2497 1338 4309 1406
rect 2497 1282 2507 1338
rect 2563 1282 2631 1338
rect 2687 1282 2755 1338
rect 2811 1282 2879 1338
rect 2935 1282 3003 1338
rect 3059 1282 3127 1338
rect 3183 1282 3251 1338
rect 3307 1282 3375 1338
rect 3431 1282 3499 1338
rect 3555 1282 3623 1338
rect 3679 1282 3747 1338
rect 3803 1282 3871 1338
rect 3927 1282 3995 1338
rect 4051 1282 4119 1338
rect 4175 1282 4243 1338
rect 4299 1282 4309 1338
rect 2497 1214 4309 1282
rect 2497 1158 2507 1214
rect 2563 1158 2631 1214
rect 2687 1158 2755 1214
rect 2811 1158 2879 1214
rect 2935 1158 3003 1214
rect 3059 1158 3127 1214
rect 3183 1158 3251 1214
rect 3307 1158 3375 1214
rect 3431 1158 3499 1214
rect 3555 1158 3623 1214
rect 3679 1158 3747 1214
rect 3803 1158 3871 1214
rect 3927 1158 3995 1214
rect 4051 1158 4119 1214
rect 4175 1158 4243 1214
rect 4299 1158 4309 1214
rect 2497 1090 4309 1158
rect 2497 1034 2507 1090
rect 2563 1034 2631 1090
rect 2687 1034 2755 1090
rect 2811 1034 2879 1090
rect 2935 1034 3003 1090
rect 3059 1034 3127 1090
rect 3183 1034 3251 1090
rect 3307 1034 3375 1090
rect 3431 1034 3499 1090
rect 3555 1034 3623 1090
rect 3679 1034 3747 1090
rect 3803 1034 3871 1090
rect 3927 1034 3995 1090
rect 4051 1034 4119 1090
rect 4175 1034 4243 1090
rect 4299 1034 4309 1090
rect 2497 966 4309 1034
rect 2497 910 2507 966
rect 2563 910 2631 966
rect 2687 910 2755 966
rect 2811 910 2879 966
rect 2935 910 3003 966
rect 3059 910 3127 966
rect 3183 910 3251 966
rect 3307 910 3375 966
rect 3431 910 3499 966
rect 3555 910 3623 966
rect 3679 910 3747 966
rect 3803 910 3871 966
rect 3927 910 3995 966
rect 4051 910 4119 966
rect 4175 910 4243 966
rect 4299 910 4309 966
rect 2497 842 4309 910
rect 2497 786 2507 842
rect 2563 786 2631 842
rect 2687 786 2755 842
rect 2811 786 2879 842
rect 2935 786 3003 842
rect 3059 786 3127 842
rect 3183 786 3251 842
rect 3307 786 3375 842
rect 3431 786 3499 842
rect 3555 786 3623 842
rect 3679 786 3747 842
rect 3803 786 3871 842
rect 3927 786 3995 842
rect 4051 786 4119 842
rect 4175 786 4243 842
rect 4299 786 4309 842
rect 2497 718 4309 786
rect 2497 662 2507 718
rect 2563 662 2631 718
rect 2687 662 2755 718
rect 2811 662 2879 718
rect 2935 662 3003 718
rect 3059 662 3127 718
rect 3183 662 3251 718
rect 3307 662 3375 718
rect 3431 662 3499 718
rect 3555 662 3623 718
rect 3679 662 3747 718
rect 3803 662 3871 718
rect 3927 662 3995 718
rect 4051 662 4119 718
rect 4175 662 4243 718
rect 4299 662 4309 718
rect 2497 594 4309 662
rect 2497 538 2507 594
rect 2563 538 2631 594
rect 2687 538 2755 594
rect 2811 538 2879 594
rect 2935 538 3003 594
rect 3059 538 3127 594
rect 3183 538 3251 594
rect 3307 538 3375 594
rect 3431 538 3499 594
rect 3555 538 3623 594
rect 3679 538 3747 594
rect 3803 538 3871 594
rect 3927 538 3995 594
rect 4051 538 4119 594
rect 4175 538 4243 594
rect 4299 538 4309 594
rect 2497 470 4309 538
rect 2497 414 2507 470
rect 2563 414 2631 470
rect 2687 414 2755 470
rect 2811 414 2879 470
rect 2935 414 3003 470
rect 3059 414 3127 470
rect 3183 414 3251 470
rect 3307 414 3375 470
rect 3431 414 3499 470
rect 3555 414 3623 470
rect 3679 414 3747 470
rect 3803 414 3871 470
rect 3927 414 3995 470
rect 4051 414 4119 470
rect 4175 414 4243 470
rect 4299 414 4309 470
rect 2497 346 4309 414
rect 2497 290 2507 346
rect 2563 290 2631 346
rect 2687 290 2755 346
rect 2811 290 2879 346
rect 2935 290 3003 346
rect 3059 290 3127 346
rect 3183 290 3251 346
rect 3307 290 3375 346
rect 3431 290 3499 346
rect 3555 290 3623 346
rect 3679 290 3747 346
rect 3803 290 3871 346
rect 3927 290 3995 346
rect 4051 290 4119 346
rect 4175 290 4243 346
rect 4299 290 4309 346
rect 2497 222 4309 290
rect 2497 166 2507 222
rect 2563 166 2631 222
rect 2687 166 2755 222
rect 2811 166 2879 222
rect 2935 166 3003 222
rect 3059 166 3127 222
rect 3183 166 3251 222
rect 3307 166 3375 222
rect 3431 166 3499 222
rect 3555 166 3623 222
rect 3679 166 3747 222
rect 3803 166 3871 222
rect 3927 166 3995 222
rect 4051 166 4119 222
rect 4175 166 4243 222
rect 4299 166 4309 222
rect 2497 98 4309 166
rect 2497 42 2507 98
rect 2563 42 2631 98
rect 2687 42 2755 98
rect 2811 42 2879 98
rect 2935 42 3003 98
rect 3059 42 3127 98
rect 3183 42 3251 98
rect 3307 42 3375 98
rect 3431 42 3499 98
rect 3555 42 3623 98
rect 3679 42 3747 98
rect 3803 42 3871 98
rect 3927 42 3995 98
rect 4051 42 4119 98
rect 4175 42 4243 98
rect 4299 42 4309 98
rect 2497 32 4309 42
rect 6358 2950 7426 2960
rect 6358 2894 6368 2950
rect 6424 2894 6492 2950
rect 6548 2894 6616 2950
rect 6672 2894 6740 2950
rect 6796 2894 6864 2950
rect 6920 2894 6988 2950
rect 7044 2894 7112 2950
rect 7168 2894 7236 2950
rect 7292 2894 7360 2950
rect 7416 2894 7426 2950
rect 6358 2826 7426 2894
rect 6358 2770 6368 2826
rect 6424 2770 6492 2826
rect 6548 2770 6616 2826
rect 6672 2770 6740 2826
rect 6796 2770 6864 2826
rect 6920 2770 6988 2826
rect 7044 2770 7112 2826
rect 7168 2770 7236 2826
rect 7292 2770 7360 2826
rect 7416 2770 7426 2826
rect 6358 2702 7426 2770
rect 6358 2646 6368 2702
rect 6424 2646 6492 2702
rect 6548 2646 6616 2702
rect 6672 2646 6740 2702
rect 6796 2646 6864 2702
rect 6920 2646 6988 2702
rect 7044 2646 7112 2702
rect 7168 2646 7236 2702
rect 7292 2646 7360 2702
rect 7416 2646 7426 2702
rect 6358 2578 7426 2646
rect 6358 2522 6368 2578
rect 6424 2522 6492 2578
rect 6548 2522 6616 2578
rect 6672 2522 6740 2578
rect 6796 2522 6864 2578
rect 6920 2522 6988 2578
rect 7044 2522 7112 2578
rect 7168 2522 7236 2578
rect 7292 2522 7360 2578
rect 7416 2522 7426 2578
rect 6358 2454 7426 2522
rect 6358 2398 6368 2454
rect 6424 2398 6492 2454
rect 6548 2398 6616 2454
rect 6672 2398 6740 2454
rect 6796 2398 6864 2454
rect 6920 2398 6988 2454
rect 7044 2398 7112 2454
rect 7168 2398 7236 2454
rect 7292 2398 7360 2454
rect 7416 2398 7426 2454
rect 6358 2330 7426 2398
rect 6358 2274 6368 2330
rect 6424 2274 6492 2330
rect 6548 2274 6616 2330
rect 6672 2274 6740 2330
rect 6796 2274 6864 2330
rect 6920 2274 6988 2330
rect 7044 2274 7112 2330
rect 7168 2274 7236 2330
rect 7292 2274 7360 2330
rect 7416 2274 7426 2330
rect 6358 2206 7426 2274
rect 6358 2150 6368 2206
rect 6424 2150 6492 2206
rect 6548 2150 6616 2206
rect 6672 2150 6740 2206
rect 6796 2150 6864 2206
rect 6920 2150 6988 2206
rect 7044 2150 7112 2206
rect 7168 2150 7236 2206
rect 7292 2150 7360 2206
rect 7416 2150 7426 2206
rect 6358 2082 7426 2150
rect 6358 2026 6368 2082
rect 6424 2026 6492 2082
rect 6548 2026 6616 2082
rect 6672 2026 6740 2082
rect 6796 2026 6864 2082
rect 6920 2026 6988 2082
rect 7044 2026 7112 2082
rect 7168 2026 7236 2082
rect 7292 2026 7360 2082
rect 7416 2026 7426 2082
rect 6358 1958 7426 2026
rect 6358 1902 6368 1958
rect 6424 1902 6492 1958
rect 6548 1902 6616 1958
rect 6672 1902 6740 1958
rect 6796 1902 6864 1958
rect 6920 1902 6988 1958
rect 7044 1902 7112 1958
rect 7168 1902 7236 1958
rect 7292 1902 7360 1958
rect 7416 1902 7426 1958
rect 6358 1834 7426 1902
rect 6358 1778 6368 1834
rect 6424 1778 6492 1834
rect 6548 1778 6616 1834
rect 6672 1778 6740 1834
rect 6796 1778 6864 1834
rect 6920 1778 6988 1834
rect 7044 1778 7112 1834
rect 7168 1778 7236 1834
rect 7292 1778 7360 1834
rect 7416 1778 7426 1834
rect 6358 1710 7426 1778
rect 6358 1654 6368 1710
rect 6424 1654 6492 1710
rect 6548 1654 6616 1710
rect 6672 1654 6740 1710
rect 6796 1654 6864 1710
rect 6920 1654 6988 1710
rect 7044 1654 7112 1710
rect 7168 1654 7236 1710
rect 7292 1654 7360 1710
rect 7416 1654 7426 1710
rect 6358 1586 7426 1654
rect 6358 1530 6368 1586
rect 6424 1530 6492 1586
rect 6548 1530 6616 1586
rect 6672 1530 6740 1586
rect 6796 1530 6864 1586
rect 6920 1530 6988 1586
rect 7044 1530 7112 1586
rect 7168 1530 7236 1586
rect 7292 1530 7360 1586
rect 7416 1530 7426 1586
rect 6358 1462 7426 1530
rect 6358 1406 6368 1462
rect 6424 1406 6492 1462
rect 6548 1406 6616 1462
rect 6672 1406 6740 1462
rect 6796 1406 6864 1462
rect 6920 1406 6988 1462
rect 7044 1406 7112 1462
rect 7168 1406 7236 1462
rect 7292 1406 7360 1462
rect 7416 1406 7426 1462
rect 6358 1338 7426 1406
rect 6358 1282 6368 1338
rect 6424 1282 6492 1338
rect 6548 1282 6616 1338
rect 6672 1282 6740 1338
rect 6796 1282 6864 1338
rect 6920 1282 6988 1338
rect 7044 1282 7112 1338
rect 7168 1282 7236 1338
rect 7292 1282 7360 1338
rect 7416 1282 7426 1338
rect 6358 1214 7426 1282
rect 6358 1158 6368 1214
rect 6424 1158 6492 1214
rect 6548 1158 6616 1214
rect 6672 1158 6740 1214
rect 6796 1158 6864 1214
rect 6920 1158 6988 1214
rect 7044 1158 7112 1214
rect 7168 1158 7236 1214
rect 7292 1158 7360 1214
rect 7416 1158 7426 1214
rect 6358 1090 7426 1158
rect 6358 1034 6368 1090
rect 6424 1034 6492 1090
rect 6548 1034 6616 1090
rect 6672 1034 6740 1090
rect 6796 1034 6864 1090
rect 6920 1034 6988 1090
rect 7044 1034 7112 1090
rect 7168 1034 7236 1090
rect 7292 1034 7360 1090
rect 7416 1034 7426 1090
rect 6358 966 7426 1034
rect 6358 910 6368 966
rect 6424 910 6492 966
rect 6548 910 6616 966
rect 6672 910 6740 966
rect 6796 910 6864 966
rect 6920 910 6988 966
rect 7044 910 7112 966
rect 7168 910 7236 966
rect 7292 910 7360 966
rect 7416 910 7426 966
rect 6358 842 7426 910
rect 6358 786 6368 842
rect 6424 786 6492 842
rect 6548 786 6616 842
rect 6672 786 6740 842
rect 6796 786 6864 842
rect 6920 786 6988 842
rect 7044 786 7112 842
rect 7168 786 7236 842
rect 7292 786 7360 842
rect 7416 786 7426 842
rect 6358 718 7426 786
rect 6358 662 6368 718
rect 6424 662 6492 718
rect 6548 662 6616 718
rect 6672 662 6740 718
rect 6796 662 6864 718
rect 6920 662 6988 718
rect 7044 662 7112 718
rect 7168 662 7236 718
rect 7292 662 7360 718
rect 7416 662 7426 718
rect 6358 594 7426 662
rect 6358 538 6368 594
rect 6424 538 6492 594
rect 6548 538 6616 594
rect 6672 538 6740 594
rect 6796 538 6864 594
rect 6920 538 6988 594
rect 7044 538 7112 594
rect 7168 538 7236 594
rect 7292 538 7360 594
rect 7416 538 7426 594
rect 6358 470 7426 538
rect 6358 414 6368 470
rect 6424 414 6492 470
rect 6548 414 6616 470
rect 6672 414 6740 470
rect 6796 414 6864 470
rect 6920 414 6988 470
rect 7044 414 7112 470
rect 7168 414 7236 470
rect 7292 414 7360 470
rect 7416 414 7426 470
rect 6358 346 7426 414
rect 6358 290 6368 346
rect 6424 290 6492 346
rect 6548 290 6616 346
rect 6672 290 6740 346
rect 6796 290 6864 346
rect 6920 290 6988 346
rect 7044 290 7112 346
rect 7168 290 7236 346
rect 7292 290 7360 346
rect 7416 290 7426 346
rect 6358 222 7426 290
rect 6358 166 6368 222
rect 6424 166 6492 222
rect 6548 166 6616 222
rect 6672 166 6740 222
rect 6796 166 6864 222
rect 6920 166 6988 222
rect 7044 166 7112 222
rect 7168 166 7236 222
rect 7292 166 7360 222
rect 7416 166 7426 222
rect 6358 98 7426 166
rect 6358 42 6368 98
rect 6424 42 6492 98
rect 6548 42 6616 98
rect 6672 42 6740 98
rect 6796 42 6864 98
rect 6920 42 6988 98
rect 7044 42 7112 98
rect 7168 42 7236 98
rect 7292 42 7360 98
rect 7416 42 7426 98
rect 6358 32 7426 42
rect 8741 2950 10553 2960
rect 8741 2894 8751 2950
rect 8807 2894 8875 2950
rect 8931 2894 8999 2950
rect 9055 2894 9123 2950
rect 9179 2894 9247 2950
rect 9303 2894 9371 2950
rect 9427 2894 9495 2950
rect 9551 2894 9619 2950
rect 9675 2894 9743 2950
rect 9799 2894 9867 2950
rect 9923 2894 9991 2950
rect 10047 2894 10115 2950
rect 10171 2894 10239 2950
rect 10295 2894 10363 2950
rect 10419 2894 10487 2950
rect 10543 2894 10553 2950
rect 8741 2826 10553 2894
rect 8741 2770 8751 2826
rect 8807 2770 8875 2826
rect 8931 2770 8999 2826
rect 9055 2770 9123 2826
rect 9179 2770 9247 2826
rect 9303 2770 9371 2826
rect 9427 2770 9495 2826
rect 9551 2770 9619 2826
rect 9675 2770 9743 2826
rect 9799 2770 9867 2826
rect 9923 2770 9991 2826
rect 10047 2770 10115 2826
rect 10171 2770 10239 2826
rect 10295 2770 10363 2826
rect 10419 2770 10487 2826
rect 10543 2770 10553 2826
rect 8741 2702 10553 2770
rect 8741 2646 8751 2702
rect 8807 2646 8875 2702
rect 8931 2646 8999 2702
rect 9055 2646 9123 2702
rect 9179 2646 9247 2702
rect 9303 2646 9371 2702
rect 9427 2646 9495 2702
rect 9551 2646 9619 2702
rect 9675 2646 9743 2702
rect 9799 2646 9867 2702
rect 9923 2646 9991 2702
rect 10047 2646 10115 2702
rect 10171 2646 10239 2702
rect 10295 2646 10363 2702
rect 10419 2646 10487 2702
rect 10543 2646 10553 2702
rect 8741 2578 10553 2646
rect 8741 2522 8751 2578
rect 8807 2522 8875 2578
rect 8931 2522 8999 2578
rect 9055 2522 9123 2578
rect 9179 2522 9247 2578
rect 9303 2522 9371 2578
rect 9427 2522 9495 2578
rect 9551 2522 9619 2578
rect 9675 2522 9743 2578
rect 9799 2522 9867 2578
rect 9923 2522 9991 2578
rect 10047 2522 10115 2578
rect 10171 2522 10239 2578
rect 10295 2522 10363 2578
rect 10419 2522 10487 2578
rect 10543 2522 10553 2578
rect 8741 2454 10553 2522
rect 8741 2398 8751 2454
rect 8807 2398 8875 2454
rect 8931 2398 8999 2454
rect 9055 2398 9123 2454
rect 9179 2398 9247 2454
rect 9303 2398 9371 2454
rect 9427 2398 9495 2454
rect 9551 2398 9619 2454
rect 9675 2398 9743 2454
rect 9799 2398 9867 2454
rect 9923 2398 9991 2454
rect 10047 2398 10115 2454
rect 10171 2398 10239 2454
rect 10295 2398 10363 2454
rect 10419 2398 10487 2454
rect 10543 2398 10553 2454
rect 8741 2330 10553 2398
rect 8741 2274 8751 2330
rect 8807 2274 8875 2330
rect 8931 2274 8999 2330
rect 9055 2274 9123 2330
rect 9179 2274 9247 2330
rect 9303 2274 9371 2330
rect 9427 2274 9495 2330
rect 9551 2274 9619 2330
rect 9675 2274 9743 2330
rect 9799 2274 9867 2330
rect 9923 2274 9991 2330
rect 10047 2274 10115 2330
rect 10171 2274 10239 2330
rect 10295 2274 10363 2330
rect 10419 2274 10487 2330
rect 10543 2274 10553 2330
rect 8741 2206 10553 2274
rect 8741 2150 8751 2206
rect 8807 2150 8875 2206
rect 8931 2150 8999 2206
rect 9055 2150 9123 2206
rect 9179 2150 9247 2206
rect 9303 2150 9371 2206
rect 9427 2150 9495 2206
rect 9551 2150 9619 2206
rect 9675 2150 9743 2206
rect 9799 2150 9867 2206
rect 9923 2150 9991 2206
rect 10047 2150 10115 2206
rect 10171 2150 10239 2206
rect 10295 2150 10363 2206
rect 10419 2150 10487 2206
rect 10543 2150 10553 2206
rect 8741 2082 10553 2150
rect 8741 2026 8751 2082
rect 8807 2026 8875 2082
rect 8931 2026 8999 2082
rect 9055 2026 9123 2082
rect 9179 2026 9247 2082
rect 9303 2026 9371 2082
rect 9427 2026 9495 2082
rect 9551 2026 9619 2082
rect 9675 2026 9743 2082
rect 9799 2026 9867 2082
rect 9923 2026 9991 2082
rect 10047 2026 10115 2082
rect 10171 2026 10239 2082
rect 10295 2026 10363 2082
rect 10419 2026 10487 2082
rect 10543 2026 10553 2082
rect 8741 1958 10553 2026
rect 8741 1902 8751 1958
rect 8807 1902 8875 1958
rect 8931 1902 8999 1958
rect 9055 1902 9123 1958
rect 9179 1902 9247 1958
rect 9303 1902 9371 1958
rect 9427 1902 9495 1958
rect 9551 1902 9619 1958
rect 9675 1902 9743 1958
rect 9799 1902 9867 1958
rect 9923 1902 9991 1958
rect 10047 1902 10115 1958
rect 10171 1902 10239 1958
rect 10295 1902 10363 1958
rect 10419 1902 10487 1958
rect 10543 1902 10553 1958
rect 8741 1834 10553 1902
rect 8741 1778 8751 1834
rect 8807 1778 8875 1834
rect 8931 1778 8999 1834
rect 9055 1778 9123 1834
rect 9179 1778 9247 1834
rect 9303 1778 9371 1834
rect 9427 1778 9495 1834
rect 9551 1778 9619 1834
rect 9675 1778 9743 1834
rect 9799 1778 9867 1834
rect 9923 1778 9991 1834
rect 10047 1778 10115 1834
rect 10171 1778 10239 1834
rect 10295 1778 10363 1834
rect 10419 1778 10487 1834
rect 10543 1778 10553 1834
rect 8741 1710 10553 1778
rect 8741 1654 8751 1710
rect 8807 1654 8875 1710
rect 8931 1654 8999 1710
rect 9055 1654 9123 1710
rect 9179 1654 9247 1710
rect 9303 1654 9371 1710
rect 9427 1654 9495 1710
rect 9551 1654 9619 1710
rect 9675 1654 9743 1710
rect 9799 1654 9867 1710
rect 9923 1654 9991 1710
rect 10047 1654 10115 1710
rect 10171 1654 10239 1710
rect 10295 1654 10363 1710
rect 10419 1654 10487 1710
rect 10543 1654 10553 1710
rect 8741 1586 10553 1654
rect 8741 1530 8751 1586
rect 8807 1530 8875 1586
rect 8931 1530 8999 1586
rect 9055 1530 9123 1586
rect 9179 1530 9247 1586
rect 9303 1530 9371 1586
rect 9427 1530 9495 1586
rect 9551 1530 9619 1586
rect 9675 1530 9743 1586
rect 9799 1530 9867 1586
rect 9923 1530 9991 1586
rect 10047 1530 10115 1586
rect 10171 1530 10239 1586
rect 10295 1530 10363 1586
rect 10419 1530 10487 1586
rect 10543 1530 10553 1586
rect 8741 1462 10553 1530
rect 8741 1406 8751 1462
rect 8807 1406 8875 1462
rect 8931 1406 8999 1462
rect 9055 1406 9123 1462
rect 9179 1406 9247 1462
rect 9303 1406 9371 1462
rect 9427 1406 9495 1462
rect 9551 1406 9619 1462
rect 9675 1406 9743 1462
rect 9799 1406 9867 1462
rect 9923 1406 9991 1462
rect 10047 1406 10115 1462
rect 10171 1406 10239 1462
rect 10295 1406 10363 1462
rect 10419 1406 10487 1462
rect 10543 1406 10553 1462
rect 8741 1338 10553 1406
rect 8741 1282 8751 1338
rect 8807 1282 8875 1338
rect 8931 1282 8999 1338
rect 9055 1282 9123 1338
rect 9179 1282 9247 1338
rect 9303 1282 9371 1338
rect 9427 1282 9495 1338
rect 9551 1282 9619 1338
rect 9675 1282 9743 1338
rect 9799 1282 9867 1338
rect 9923 1282 9991 1338
rect 10047 1282 10115 1338
rect 10171 1282 10239 1338
rect 10295 1282 10363 1338
rect 10419 1282 10487 1338
rect 10543 1282 10553 1338
rect 8741 1214 10553 1282
rect 8741 1158 8751 1214
rect 8807 1158 8875 1214
rect 8931 1158 8999 1214
rect 9055 1158 9123 1214
rect 9179 1158 9247 1214
rect 9303 1158 9371 1214
rect 9427 1158 9495 1214
rect 9551 1158 9619 1214
rect 9675 1158 9743 1214
rect 9799 1158 9867 1214
rect 9923 1158 9991 1214
rect 10047 1158 10115 1214
rect 10171 1158 10239 1214
rect 10295 1158 10363 1214
rect 10419 1158 10487 1214
rect 10543 1158 10553 1214
rect 8741 1090 10553 1158
rect 8741 1034 8751 1090
rect 8807 1034 8875 1090
rect 8931 1034 8999 1090
rect 9055 1034 9123 1090
rect 9179 1034 9247 1090
rect 9303 1034 9371 1090
rect 9427 1034 9495 1090
rect 9551 1034 9619 1090
rect 9675 1034 9743 1090
rect 9799 1034 9867 1090
rect 9923 1034 9991 1090
rect 10047 1034 10115 1090
rect 10171 1034 10239 1090
rect 10295 1034 10363 1090
rect 10419 1034 10487 1090
rect 10543 1034 10553 1090
rect 8741 966 10553 1034
rect 8741 910 8751 966
rect 8807 910 8875 966
rect 8931 910 8999 966
rect 9055 910 9123 966
rect 9179 910 9247 966
rect 9303 910 9371 966
rect 9427 910 9495 966
rect 9551 910 9619 966
rect 9675 910 9743 966
rect 9799 910 9867 966
rect 9923 910 9991 966
rect 10047 910 10115 966
rect 10171 910 10239 966
rect 10295 910 10363 966
rect 10419 910 10487 966
rect 10543 910 10553 966
rect 8741 842 10553 910
rect 8741 786 8751 842
rect 8807 786 8875 842
rect 8931 786 8999 842
rect 9055 786 9123 842
rect 9179 786 9247 842
rect 9303 786 9371 842
rect 9427 786 9495 842
rect 9551 786 9619 842
rect 9675 786 9743 842
rect 9799 786 9867 842
rect 9923 786 9991 842
rect 10047 786 10115 842
rect 10171 786 10239 842
rect 10295 786 10363 842
rect 10419 786 10487 842
rect 10543 786 10553 842
rect 8741 718 10553 786
rect 8741 662 8751 718
rect 8807 662 8875 718
rect 8931 662 8999 718
rect 9055 662 9123 718
rect 9179 662 9247 718
rect 9303 662 9371 718
rect 9427 662 9495 718
rect 9551 662 9619 718
rect 9675 662 9743 718
rect 9799 662 9867 718
rect 9923 662 9991 718
rect 10047 662 10115 718
rect 10171 662 10239 718
rect 10295 662 10363 718
rect 10419 662 10487 718
rect 10543 662 10553 718
rect 8741 594 10553 662
rect 8741 538 8751 594
rect 8807 538 8875 594
rect 8931 538 8999 594
rect 9055 538 9123 594
rect 9179 538 9247 594
rect 9303 538 9371 594
rect 9427 538 9495 594
rect 9551 538 9619 594
rect 9675 538 9743 594
rect 9799 538 9867 594
rect 9923 538 9991 594
rect 10047 538 10115 594
rect 10171 538 10239 594
rect 10295 538 10363 594
rect 10419 538 10487 594
rect 10543 538 10553 594
rect 8741 470 10553 538
rect 8741 414 8751 470
rect 8807 414 8875 470
rect 8931 414 8999 470
rect 9055 414 9123 470
rect 9179 414 9247 470
rect 9303 414 9371 470
rect 9427 414 9495 470
rect 9551 414 9619 470
rect 9675 414 9743 470
rect 9799 414 9867 470
rect 9923 414 9991 470
rect 10047 414 10115 470
rect 10171 414 10239 470
rect 10295 414 10363 470
rect 10419 414 10487 470
rect 10543 414 10553 470
rect 8741 346 10553 414
rect 8741 290 8751 346
rect 8807 290 8875 346
rect 8931 290 8999 346
rect 9055 290 9123 346
rect 9179 290 9247 346
rect 9303 290 9371 346
rect 9427 290 9495 346
rect 9551 290 9619 346
rect 9675 290 9743 346
rect 9799 290 9867 346
rect 9923 290 9991 346
rect 10047 290 10115 346
rect 10171 290 10239 346
rect 10295 290 10363 346
rect 10419 290 10487 346
rect 10543 290 10553 346
rect 8741 222 10553 290
rect 8741 166 8751 222
rect 8807 166 8875 222
rect 8931 166 8999 222
rect 9055 166 9123 222
rect 9179 166 9247 222
rect 9303 166 9371 222
rect 9427 166 9495 222
rect 9551 166 9619 222
rect 9675 166 9743 222
rect 9799 166 9867 222
rect 9923 166 9991 222
rect 10047 166 10115 222
rect 10171 166 10239 222
rect 10295 166 10363 222
rect 10419 166 10487 222
rect 10543 166 10553 222
rect 8741 98 10553 166
rect 8741 42 8751 98
rect 8807 42 8875 98
rect 8931 42 8999 98
rect 9055 42 9123 98
rect 9179 42 9247 98
rect 9303 42 9371 98
rect 9427 42 9495 98
rect 9551 42 9619 98
rect 9675 42 9743 98
rect 9799 42 9867 98
rect 9923 42 9991 98
rect 10047 42 10115 98
rect 10171 42 10239 98
rect 10295 42 10363 98
rect 10419 42 10487 98
rect 10543 42 10553 98
rect 8741 32 10553 42
rect 12842 2950 13910 2960
rect 12842 2894 12852 2950
rect 12908 2894 12976 2950
rect 13032 2894 13100 2950
rect 13156 2894 13224 2950
rect 13280 2894 13348 2950
rect 13404 2894 13472 2950
rect 13528 2894 13596 2950
rect 13652 2894 13720 2950
rect 13776 2894 13844 2950
rect 13900 2894 13910 2950
rect 12842 2826 13910 2894
rect 12842 2770 12852 2826
rect 12908 2770 12976 2826
rect 13032 2770 13100 2826
rect 13156 2770 13224 2826
rect 13280 2770 13348 2826
rect 13404 2770 13472 2826
rect 13528 2770 13596 2826
rect 13652 2770 13720 2826
rect 13776 2770 13844 2826
rect 13900 2770 13910 2826
rect 12842 2702 13910 2770
rect 12842 2646 12852 2702
rect 12908 2646 12976 2702
rect 13032 2646 13100 2702
rect 13156 2646 13224 2702
rect 13280 2646 13348 2702
rect 13404 2646 13472 2702
rect 13528 2646 13596 2702
rect 13652 2646 13720 2702
rect 13776 2646 13844 2702
rect 13900 2646 13910 2702
rect 12842 2578 13910 2646
rect 12842 2522 12852 2578
rect 12908 2522 12976 2578
rect 13032 2522 13100 2578
rect 13156 2522 13224 2578
rect 13280 2522 13348 2578
rect 13404 2522 13472 2578
rect 13528 2522 13596 2578
rect 13652 2522 13720 2578
rect 13776 2522 13844 2578
rect 13900 2522 13910 2578
rect 12842 2454 13910 2522
rect 12842 2398 12852 2454
rect 12908 2398 12976 2454
rect 13032 2398 13100 2454
rect 13156 2398 13224 2454
rect 13280 2398 13348 2454
rect 13404 2398 13472 2454
rect 13528 2398 13596 2454
rect 13652 2398 13720 2454
rect 13776 2398 13844 2454
rect 13900 2398 13910 2454
rect 12842 2330 13910 2398
rect 12842 2274 12852 2330
rect 12908 2274 12976 2330
rect 13032 2274 13100 2330
rect 13156 2274 13224 2330
rect 13280 2274 13348 2330
rect 13404 2274 13472 2330
rect 13528 2274 13596 2330
rect 13652 2274 13720 2330
rect 13776 2274 13844 2330
rect 13900 2274 13910 2330
rect 12842 2206 13910 2274
rect 12842 2150 12852 2206
rect 12908 2150 12976 2206
rect 13032 2150 13100 2206
rect 13156 2150 13224 2206
rect 13280 2150 13348 2206
rect 13404 2150 13472 2206
rect 13528 2150 13596 2206
rect 13652 2150 13720 2206
rect 13776 2150 13844 2206
rect 13900 2150 13910 2206
rect 12842 2082 13910 2150
rect 12842 2026 12852 2082
rect 12908 2026 12976 2082
rect 13032 2026 13100 2082
rect 13156 2026 13224 2082
rect 13280 2026 13348 2082
rect 13404 2026 13472 2082
rect 13528 2026 13596 2082
rect 13652 2026 13720 2082
rect 13776 2026 13844 2082
rect 13900 2026 13910 2082
rect 12842 1958 13910 2026
rect 12842 1902 12852 1958
rect 12908 1902 12976 1958
rect 13032 1902 13100 1958
rect 13156 1902 13224 1958
rect 13280 1902 13348 1958
rect 13404 1902 13472 1958
rect 13528 1902 13596 1958
rect 13652 1902 13720 1958
rect 13776 1902 13844 1958
rect 13900 1902 13910 1958
rect 12842 1834 13910 1902
rect 12842 1778 12852 1834
rect 12908 1778 12976 1834
rect 13032 1778 13100 1834
rect 13156 1778 13224 1834
rect 13280 1778 13348 1834
rect 13404 1778 13472 1834
rect 13528 1778 13596 1834
rect 13652 1778 13720 1834
rect 13776 1778 13844 1834
rect 13900 1778 13910 1834
rect 12842 1710 13910 1778
rect 12842 1654 12852 1710
rect 12908 1654 12976 1710
rect 13032 1654 13100 1710
rect 13156 1654 13224 1710
rect 13280 1654 13348 1710
rect 13404 1654 13472 1710
rect 13528 1654 13596 1710
rect 13652 1654 13720 1710
rect 13776 1654 13844 1710
rect 13900 1654 13910 1710
rect 12842 1586 13910 1654
rect 12842 1530 12852 1586
rect 12908 1530 12976 1586
rect 13032 1530 13100 1586
rect 13156 1530 13224 1586
rect 13280 1530 13348 1586
rect 13404 1530 13472 1586
rect 13528 1530 13596 1586
rect 13652 1530 13720 1586
rect 13776 1530 13844 1586
rect 13900 1530 13910 1586
rect 12842 1462 13910 1530
rect 12842 1406 12852 1462
rect 12908 1406 12976 1462
rect 13032 1406 13100 1462
rect 13156 1406 13224 1462
rect 13280 1406 13348 1462
rect 13404 1406 13472 1462
rect 13528 1406 13596 1462
rect 13652 1406 13720 1462
rect 13776 1406 13844 1462
rect 13900 1406 13910 1462
rect 12842 1338 13910 1406
rect 12842 1282 12852 1338
rect 12908 1282 12976 1338
rect 13032 1282 13100 1338
rect 13156 1282 13224 1338
rect 13280 1282 13348 1338
rect 13404 1282 13472 1338
rect 13528 1282 13596 1338
rect 13652 1282 13720 1338
rect 13776 1282 13844 1338
rect 13900 1282 13910 1338
rect 12842 1214 13910 1282
rect 12842 1158 12852 1214
rect 12908 1158 12976 1214
rect 13032 1158 13100 1214
rect 13156 1158 13224 1214
rect 13280 1158 13348 1214
rect 13404 1158 13472 1214
rect 13528 1158 13596 1214
rect 13652 1158 13720 1214
rect 13776 1158 13844 1214
rect 13900 1158 13910 1214
rect 12842 1090 13910 1158
rect 12842 1034 12852 1090
rect 12908 1034 12976 1090
rect 13032 1034 13100 1090
rect 13156 1034 13224 1090
rect 13280 1034 13348 1090
rect 13404 1034 13472 1090
rect 13528 1034 13596 1090
rect 13652 1034 13720 1090
rect 13776 1034 13844 1090
rect 13900 1034 13910 1090
rect 12842 966 13910 1034
rect 12842 910 12852 966
rect 12908 910 12976 966
rect 13032 910 13100 966
rect 13156 910 13224 966
rect 13280 910 13348 966
rect 13404 910 13472 966
rect 13528 910 13596 966
rect 13652 910 13720 966
rect 13776 910 13844 966
rect 13900 910 13910 966
rect 12842 842 13910 910
rect 12842 786 12852 842
rect 12908 786 12976 842
rect 13032 786 13100 842
rect 13156 786 13224 842
rect 13280 786 13348 842
rect 13404 786 13472 842
rect 13528 786 13596 842
rect 13652 786 13720 842
rect 13776 786 13844 842
rect 13900 786 13910 842
rect 12842 718 13910 786
rect 12842 662 12852 718
rect 12908 662 12976 718
rect 13032 662 13100 718
rect 13156 662 13224 718
rect 13280 662 13348 718
rect 13404 662 13472 718
rect 13528 662 13596 718
rect 13652 662 13720 718
rect 13776 662 13844 718
rect 13900 662 13910 718
rect 12842 594 13910 662
rect 12842 538 12852 594
rect 12908 538 12976 594
rect 13032 538 13100 594
rect 13156 538 13224 594
rect 13280 538 13348 594
rect 13404 538 13472 594
rect 13528 538 13596 594
rect 13652 538 13720 594
rect 13776 538 13844 594
rect 13900 538 13910 594
rect 12842 470 13910 538
rect 12842 414 12852 470
rect 12908 414 12976 470
rect 13032 414 13100 470
rect 13156 414 13224 470
rect 13280 414 13348 470
rect 13404 414 13472 470
rect 13528 414 13596 470
rect 13652 414 13720 470
rect 13776 414 13844 470
rect 13900 414 13910 470
rect 12842 346 13910 414
rect 12842 290 12852 346
rect 12908 290 12976 346
rect 13032 290 13100 346
rect 13156 290 13224 346
rect 13280 290 13348 346
rect 13404 290 13472 346
rect 13528 290 13596 346
rect 13652 290 13720 346
rect 13776 290 13844 346
rect 13900 290 13910 346
rect 12842 222 13910 290
rect 12842 166 12852 222
rect 12908 166 12976 222
rect 13032 166 13100 222
rect 13156 166 13224 222
rect 13280 166 13348 222
rect 13404 166 13472 222
rect 13528 166 13596 222
rect 13652 166 13720 222
rect 13776 166 13844 222
rect 13900 166 13910 222
rect 12842 98 13910 166
rect 12842 42 12852 98
rect 12908 42 12976 98
rect 13032 42 13100 98
rect 13156 42 13224 98
rect 13280 42 13348 98
rect 13404 42 13472 98
rect 13528 42 13596 98
rect 13652 42 13720 98
rect 13776 42 13844 98
rect 13900 42 13910 98
rect 12842 32 13910 42
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_0
timestamp 1755005639
transform 1 0 14795 0 1 35896
box 0 0 1 1
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_1
timestamp 1755005639
transform 1 0 14795 0 1 50296
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_0
timestamp 1755005639
transform 1 0 9647 0 1 4696
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_1
timestamp 1755005639
transform 1 0 9647 0 1 7896
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_2
timestamp 1755005639
transform 1 0 11575 0 1 14296
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_3
timestamp 1755005639
transform 1 0 11575 0 1 17496
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_4
timestamp 1755005639
transform 1 0 11575 0 1 20696
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_5
timestamp 1755005639
transform 1 0 11575 0 1 23896
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_6
timestamp 1755005639
transform 1 0 9647 0 1 1496
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_7
timestamp 1755005639
transform 1 0 5331 0 1 17496
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_8
timestamp 1755005639
transform 1 0 5331 0 1 20696
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_9
timestamp 1755005639
transform 1 0 5331 0 1 23896
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_10
timestamp 1755005639
transform 1 0 3403 0 1 1496
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_11
timestamp 1755005639
transform 1 0 3403 0 1 4696
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_12
timestamp 1755005639
transform 1 0 3403 0 1 7896
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_13
timestamp 1755005639
transform 1 0 5331 0 1 14296
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_14
timestamp 1755005639
transform 1 0 5331 0 1 30296
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_15
timestamp 1755005639
transform 1 0 9647 0 1 33496
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_16
timestamp 1755005639
transform 1 0 11575 0 1 30296
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_0
timestamp 1755005639
transform 1 0 14795 0 1 35896
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_1
timestamp 1755005639
transform 1 0 14795 0 1 50296
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_0
timestamp 1755005639
transform 1 0 9647 0 1 11896
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_1
timestamp 1755005639
transform 1 0 11575 0 1 10296
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_2
timestamp 1755005639
transform 1 0 5331 0 1 10296
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_3
timestamp 1755005639
transform 1 0 3403 0 1 11896
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_4
timestamp 1755005639
transform 1 0 5331 0 1 27896
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_5
timestamp 1755005639
transform 1 0 3403 0 1 26296
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_6
timestamp 1755005639
transform 1 0 11575 0 1 27896
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_7
timestamp 1755005639
transform 1 0 11575 0 1 39096
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_8
timestamp 1755005639
transform 1 0 11575 0 1 40696
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_9
timestamp 1755005639
transform 1 0 11575 0 1 42296
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_10
timestamp 1755005639
transform 1 0 9647 0 1 26296
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_11
timestamp 1755005639
transform 1 0 9647 0 1 43896
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_0
timestamp 1755005639
transform 1 0 13376 0 1 11896
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_1
timestamp 1755005639
transform 1 0 6892 0 1 11896
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_2
timestamp 1755005639
transform 1 0 1602 0 1 10296
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_3
timestamp 1755005639
transform 1 0 6892 0 1 26296
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_4
timestamp 1755005639
transform 1 0 13376 0 1 43896
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_5
timestamp 1755005639
transform 1 0 13376 0 1 26296
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_6
timestamp 1755005639
transform 1 0 8086 0 1 39096
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_7
timestamp 1755005639
transform 1 0 8086 0 1 40696
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_8
timestamp 1755005639
transform 1 0 8086 0 1 27896
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_9
timestamp 1755005639
transform 1 0 8086 0 1 10296
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_10
timestamp 1755005639
transform 1 0 8086 0 1 42296
box 0 0 1 1
use M3_M2_CDNS_40661953145782  M3_M2_CDNS_40661953145782_0
timestamp 1755005639
transform 1 0 4498 0 1 45489
box 0 0 1 1
use M3_M2_CDNS_40661953145782  M3_M2_CDNS_40661953145782_1
timestamp 1755005639
transform 1 0 4498 0 1 40955
box 0 0 1 1
use M3_M2_CDNS_40661953145782  M3_M2_CDNS_40661953145782_2
timestamp 1755005639
transform 1 0 4498 0 1 43190
box 0 0 1 1
use M3_M2_CDNS_40661953145783  M3_M2_CDNS_40661953145783_0
timestamp 1755005639
transform 1 0 2023 0 1 27889
box 0 0 1 1
use M3_M2_CDNS_40661953145783  M3_M2_CDNS_40661953145783_1
timestamp 1755005639
transform 1 0 1899 0 1 27891
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_0
timestamp 1755005639
transform 1 0 6110 0 1 39343
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_1
timestamp 1755005639
transform 1 0 5490 0 1 44497
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_2
timestamp 1755005639
transform 1 0 6422 0 1 45836
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_3
timestamp 1755005639
transform 1 0 4622 0 1 45365
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_4
timestamp 1755005639
transform 1 0 4746 0 1 45241
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_5
timestamp 1755005639
transform 1 0 7166 0 1 45092
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_6
timestamp 1755005639
transform 1 0 7042 0 1 45216
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_7
timestamp 1755005639
transform 1 0 4870 0 1 45117
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_8
timestamp 1755005639
transform 1 0 5738 0 1 39715
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_9
timestamp 1755005639
transform 1 0 5862 0 1 39591
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_10
timestamp 1755005639
transform 1 0 5986 0 1 39467
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_11
timestamp 1755005639
transform 1 0 4622 0 1 40831
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_12
timestamp 1755005639
transform 1 0 4746 0 1 40707
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_13
timestamp 1755005639
transform 1 0 4870 0 1 40583
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_14
timestamp 1755005639
transform 1 0 4994 0 1 40459
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_15
timestamp 1755005639
transform 1 0 5118 0 1 40335
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_16
timestamp 1755005639
transform 1 0 5242 0 1 40211
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_17
timestamp 1755005639
transform 1 0 5366 0 1 40087
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_18
timestamp 1755005639
transform 1 0 5490 0 1 39963
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_19
timestamp 1755005639
transform 1 0 5614 0 1 39839
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_20
timestamp 1755005639
transform 1 0 5614 0 1 42074
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_21
timestamp 1755005639
transform 1 0 1527 0 1 28088
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_22
timestamp 1755005639
transform 1 0 4994 0 1 44993
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_23
timestamp 1755005639
transform 1 0 5366 0 1 44621
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_24
timestamp 1755005639
transform 1 0 6670 0 1 45588
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_25
timestamp 1755005639
transform 1 0 5490 0 1 42198
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_26
timestamp 1755005639
transform 1 0 7290 0 1 44968
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_27
timestamp 1755005639
transform 1 0 5366 0 1 42322
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_28
timestamp 1755005639
transform 1 0 6110 0 1 41578
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_29
timestamp 1755005639
transform 1 0 5986 0 1 41702
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_30
timestamp 1755005639
transform 1 0 5862 0 1 41826
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_31
timestamp 1755005639
transform 1 0 5738 0 1 41950
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_32
timestamp 1755005639
transform 1 0 5242 0 1 42446
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_33
timestamp 1755005639
transform 1 0 4622 0 1 43066
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_34
timestamp 1755005639
transform 1 0 5614 0 1 44373
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_35
timestamp 1755005639
transform 1 0 4746 0 1 42942
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_36
timestamp 1755005639
transform 1 0 4994 0 1 42694
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_37
timestamp 1755005639
transform 1 0 6546 0 1 45712
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_38
timestamp 1755005639
transform 1 0 6794 0 1 45464
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_39
timestamp 1755005639
transform 1 0 6918 0 1 45340
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_40
timestamp 1755005639
transform 1 0 4870 0 1 42818
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_41
timestamp 1755005639
transform 1 0 5118 0 1 42570
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_42
timestamp 1755005639
transform 1 0 5242 0 1 44745
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_43
timestamp 1755005639
transform 1 0 5118 0 1 44869
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_44
timestamp 1755005639
transform 1 0 6110 0 1 43877
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_45
timestamp 1755005639
transform 1 0 5986 0 1 44001
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_46
timestamp 1755005639
transform 1 0 5862 0 1 44125
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_47
timestamp 1755005639
transform 1 0 5738 0 1 44249
box 0 0 1 1
use M3_M2_CDNS_40661953145785  M3_M2_CDNS_40661953145785_0
timestamp 1755005639
transform 1 0 1651 0 1 28036
box 0 0 1 1
use M3_M2_CDNS_40661953145786  M3_M2_CDNS_40661953145786_0
timestamp 1755005639
transform 1 0 1775 0 1 27943
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_0
timestamp 1755005639
transform 1 0 13376 0 1 1496
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_1
timestamp 1755005639
transform 1 0 13376 0 1 4696
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_2
timestamp 1755005639
transform 1 0 13376 0 1 7896
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_3
timestamp 1755005639
transform 1 0 1602 0 1 20696
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_4
timestamp 1755005639
transform 1 0 1602 0 1 14296
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_5
timestamp 1755005639
transform 1 0 1602 0 1 17496
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_6
timestamp 1755005639
transform 1 0 1602 0 1 23896
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_7
timestamp 1755005639
transform 1 0 6892 0 1 1496
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_8
timestamp 1755005639
transform 1 0 6892 0 1 4696
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_9
timestamp 1755005639
transform 1 0 6892 0 1 7896
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_10
timestamp 1755005639
transform 1 0 6892 0 1 33496
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_11
timestamp 1755005639
transform 1 0 13376 0 1 33496
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_12
timestamp 1755005639
transform 1 0 8086 0 1 30296
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_13
timestamp 1755005639
transform 1 0 8086 0 1 14296
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_14
timestamp 1755005639
transform 1 0 8086 0 1 17496
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_15
timestamp 1755005639
transform 1 0 8086 0 1 20696
box 0 0 1 1
use M3_M2_CDNS_40661953145795  M3_M2_CDNS_40661953145795_16
timestamp 1755005639
transform 1 0 8086 0 1 23896
box 0 0 1 1
use M3_M2_CDNS_40661953145796  M3_M2_CDNS_40661953145796_0
timestamp 1755005639
transform 1 0 2555 0 1 34988
box 0 0 1 1
use M3_M2_CDNS_40661953145796  M3_M2_CDNS_40661953145796_1
timestamp 1755005639
transform 1 0 1183 0 1 31754
box 0 0 1 1
use M3_M2_CDNS_40661953145797  M3_M2_CDNS_40661953145797_0
timestamp 1755005639
transform 1 0 4167 0 1 33715
box 0 0 1 1
use M3_M2_CDNS_40661953145798  M3_M2_CDNS_40661953145798_0
timestamp 1755005639
transform 1 0 3919 0 1 33842
box 0 0 1 1
use M3_M2_CDNS_40661953145798  M3_M2_CDNS_40661953145798_1
timestamp 1755005639
transform 1 0 4043 0 1 33771
box 0 0 1 1
use M3_M2_CDNS_40661953145799  M3_M2_CDNS_40661953145799_0
timestamp 1755005639
transform 1 0 3795 0 1 33884
box 0 0 1 1
use M3_M2_CDNS_40661953145800  M3_M2_CDNS_40661953145800_0
timestamp 1755005639
transform 1 0 3671 0 1 33925
box 0 0 1 1
use M3_M2_CDNS_40661953145801  M3_M2_CDNS_40661953145801_0
timestamp 1755005639
transform 1 0 3547 0 1 33996
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_0
timestamp 1755005639
transform 1 0 3175 0 1 34368
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_1
timestamp 1755005639
transform 1 0 1927 0 1 31010
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_2
timestamp 1755005639
transform 1 0 2051 0 1 30886
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_3
timestamp 1755005639
transform 1 0 1307 0 1 31630
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_4
timestamp 1755005639
transform 1 0 2927 0 1 34616
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_5
timestamp 1755005639
transform 1 0 2679 0 1 34864
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_6
timestamp 1755005639
transform 1 0 3051 0 1 34492
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_7
timestamp 1755005639
transform 1 0 3423 0 1 34120
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_8
timestamp 1755005639
transform 1 0 1431 0 1 31506
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_9
timestamp 1755005639
transform 1 0 1679 0 1 31258
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_10
timestamp 1755005639
transform 1 0 1803 0 1 31134
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_11
timestamp 1755005639
transform 1 0 1555 0 1 31382
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_12
timestamp 1755005639
transform 1 0 2803 0 1 34740
box 0 0 1 1
use M3_M2_CDNS_40661953145802  M3_M2_CDNS_40661953145802_13
timestamp 1755005639
transform 1 0 3299 0 1 34244
box 0 0 1 1
use M3_M2_CDNS_40661953145803  M3_M2_CDNS_40661953145803_0
timestamp 1755005639
transform 1 0 1132 0 1 44359
box 0 0 1 1
use M3_M2_CDNS_40661953145803  M3_M2_CDNS_40661953145803_1
timestamp 1755005639
transform 1 0 1155 0 1 28411
box 0 0 1 1
use M3_M2_CDNS_40661953145804  M3_M2_CDNS_40661953145804_0
timestamp 1755005639
transform 1 0 1403 0 1 28163
box 0 0 1 1
use M3_M2_CDNS_40661953145804  M3_M2_CDNS_40661953145804_1
timestamp 1755005639
transform 1 0 1279 0 1 28287
box 0 0 1 1
use M3_M2_CDNS_40661953145804  M3_M2_CDNS_40661953145804_2
timestamp 1755005639
transform 1 0 1380 0 1 44111
box 0 0 1 1
use M3_M2_CDNS_40661953145804  M3_M2_CDNS_40661953145804_3
timestamp 1755005639
transform 1 0 1256 0 1 44235
box 0 0 1 1
use M3_M2_CDNS_40661953145804  M3_M2_CDNS_40661953145804_4
timestamp 1755005639
transform 1 0 1876 0 1 43615
box 0 0 1 1
use M3_M2_CDNS_40661953145804  M3_M2_CDNS_40661953145804_5
timestamp 1755005639
transform 1 0 1752 0 1 43739
box 0 0 1 1
use M3_M2_CDNS_40661953145804  M3_M2_CDNS_40661953145804_6
timestamp 1755005639
transform 1 0 1628 0 1 43863
box 0 0 1 1
use M3_M2_CDNS_40661953145804  M3_M2_CDNS_40661953145804_7
timestamp 1755005639
transform 1 0 1504 0 1 43987
box 0 0 1 1
use M3_M2_CDNS_40661953145804  M3_M2_CDNS_40661953145804_8
timestamp 1755005639
transform 1 0 2000 0 1 43491
box 0 0 1 1
<< properties >>
string GDS_END 7041524
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 7034136
<< end >>
