magic
tech gf180mcuD
timestamp 1755005639
<< properties >>
string GDS_END 816232
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 814756
<< end >>
