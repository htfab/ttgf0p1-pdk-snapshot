magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect 314 14615 1690 68707
<< obsm1 >>
rect -32 13108 2032 69957
<< obsm2 >>
rect 0 13611 2000 69620
<< metal3 >>
rect 0 68400 200 69678
rect 1800 68400 2000 69678
rect 0 66800 200 68200
rect 1800 66800 2000 68200
rect 0 65200 200 66600
rect 1800 65200 2000 66600
rect 0 63600 200 65000
rect 1800 63600 2000 65000
rect 0 62000 200 63400
rect 1800 62000 2000 63400
rect 0 60400 200 61800
rect 1800 60400 2000 61800
rect 0 58800 200 60200
rect 1800 58800 2000 60200
rect 0 57200 200 58600
rect 1800 57200 2000 58600
rect 0 55600 200 57000
rect 1800 55600 2000 57000
rect 0 54000 200 55400
rect 1800 54000 2000 55400
rect 0 52400 200 53800
rect 1800 52400 2000 53800
rect 0 50800 200 52200
rect 1800 50800 2000 52200
rect 0 49200 200 50600
rect 1800 49200 2000 50600
rect 0 46000 200 49000
rect 1800 46000 2000 49000
rect 0 42800 200 45800
rect 1800 42800 2000 45800
rect 0 41200 200 42600
rect 1800 41200 2000 42600
rect 0 39600 200 41000
rect 1800 39600 2000 41000
rect 0 36400 200 39400
rect 1800 36400 2000 39400
rect 0 33200 200 36200
rect 1800 33200 2000 36200
rect 0 30000 200 33000
rect 1800 30000 2000 33000
rect 0 26800 200 29800
rect 1800 26800 2000 29800
rect 0 25200 200 26600
rect 1800 25200 2000 26600
rect 0 23600 200 25000
rect 1800 23600 2000 25000
rect 0 20400 200 23400
rect 1800 20400 2000 23400
rect 0 17200 200 20200
rect 1800 17200 2000 20200
rect 0 14000 200 17000
rect 1800 14000 2000 17000
<< obsm3 >>
rect 260 68340 1740 69678
rect 200 68260 1800 68340
rect 260 66740 1740 68260
rect 200 66660 1800 66740
rect 260 65140 1740 66660
rect 200 65060 1800 65140
rect 260 63540 1740 65060
rect 200 63460 1800 63540
rect 260 61940 1740 63460
rect 200 61860 1800 61940
rect 260 60340 1740 61860
rect 200 60260 1800 60340
rect 260 58740 1740 60260
rect 200 58660 1800 58740
rect 260 57140 1740 58660
rect 200 57060 1800 57140
rect 260 55540 1740 57060
rect 200 55460 1800 55540
rect 260 53940 1740 55460
rect 200 53860 1800 53940
rect 260 52340 1740 53860
rect 200 52260 1800 52340
rect 260 50740 1740 52260
rect 200 50660 1800 50740
rect 260 49140 1740 50660
rect 200 49060 1800 49140
rect 260 45940 1740 49060
rect 200 45860 1800 45940
rect 260 42740 1740 45860
rect 200 42660 1800 42740
rect 260 41140 1740 42660
rect 200 41060 1800 41140
rect 260 39540 1740 41060
rect 200 39460 1800 39540
rect 260 36340 1740 39460
rect 200 36260 1800 36340
rect 260 33140 1740 36260
rect 200 33060 1800 33140
rect 260 29940 1740 33060
rect 200 29860 1800 29940
rect 260 26740 1740 29860
rect 200 26660 1800 26740
rect 260 25140 1740 26660
rect 200 25060 1800 25140
rect 260 23540 1740 25060
rect 200 23460 1800 23540
rect 260 20340 1740 23460
rect 200 20260 1800 20340
rect 260 17140 1740 20260
rect 200 17060 1800 17140
rect 260 14000 1740 17060
<< metal4 >>
rect 0 68400 200 69678
rect 1800 68400 2000 69678
rect 0 66800 200 68200
rect 1800 66800 2000 68200
rect 0 65200 200 66600
rect 1800 65200 2000 66600
rect 0 63600 200 65000
rect 1800 63600 2000 65000
rect 0 62000 200 63400
rect 1800 62000 2000 63400
rect 0 60400 200 61800
rect 1800 60400 2000 61800
rect 0 58800 200 60200
rect 1800 58800 2000 60200
rect 0 57200 200 58600
rect 1800 57200 2000 58600
rect 0 55600 200 57000
rect 1800 55600 2000 57000
rect 0 54000 200 55400
rect 1800 54000 2000 55400
rect 0 52400 200 53800
rect 1800 52400 2000 53800
rect 0 50800 200 52200
rect 1800 50800 2000 52200
rect 0 49200 200 50600
rect 1800 49200 2000 50600
rect 0 46000 200 49000
rect 1800 46000 2000 49000
rect 0 42800 200 45800
rect 1800 42800 2000 45800
rect 0 41200 200 42600
rect 1800 41200 2000 42600
rect 0 39600 200 41000
rect 1800 39600 2000 41000
rect 0 36400 200 39400
rect 1800 36400 2000 39400
rect 0 33200 200 36200
rect 1800 33200 2000 36200
rect 0 30000 200 33000
rect 1800 30000 2000 33000
rect 0 26800 200 29800
rect 1800 26800 2000 29800
rect 0 25200 200 26600
rect 1800 25200 2000 26600
rect 0 23600 200 25000
rect 1800 23600 2000 25000
rect 0 20400 200 23400
rect 1800 20400 2000 23400
rect 0 17200 200 20200
rect 1800 17200 2000 20200
rect 0 14000 200 17000
rect 1800 14000 2000 17000
<< obsm4 >>
rect 260 68340 1740 69678
rect 200 68260 1800 68340
rect 260 66740 1740 68260
rect 200 66660 1800 66740
rect 260 65140 1740 66660
rect 200 65060 1800 65140
rect 260 63540 1740 65060
rect 200 63460 1800 63540
rect 260 61940 1740 63460
rect 200 61860 1800 61940
rect 260 60340 1740 61860
rect 200 60260 1800 60340
rect 260 58740 1740 60260
rect 200 58660 1800 58740
rect 260 57140 1740 58660
rect 200 57060 1800 57140
rect 260 55540 1740 57060
rect 200 55460 1800 55540
rect 260 53940 1740 55460
rect 200 53860 1800 53940
rect 260 52340 1740 53860
rect 200 52260 1800 52340
rect 260 50740 1740 52260
rect 200 50660 1800 50740
rect 260 49140 1740 50660
rect 200 49060 1800 49140
rect 260 45940 1740 49060
rect 200 45860 1800 45940
rect 260 42740 1740 45860
rect 200 42660 1800 42740
rect 260 41140 1740 42660
rect 200 41060 1800 41140
rect 260 39540 1740 41060
rect 200 39460 1800 39540
rect 260 36340 1740 39460
rect 200 36260 1800 36340
rect 260 33140 1740 36260
rect 200 33060 1800 33140
rect 260 29940 1740 33060
rect 200 29860 1800 29940
rect 260 26740 1740 29860
rect 200 26660 1800 26740
rect 260 25140 1740 26660
rect 200 25060 1800 25140
rect 260 23540 1740 25060
rect 200 23460 1800 23540
rect 260 20340 1740 23460
rect 200 20260 1800 20340
rect 260 17140 1740 20260
rect 200 17060 1800 17140
rect 260 14000 1740 17060
<< metal5 >>
rect 0 68400 200 69678
rect 0 66800 200 68200
rect 0 65200 200 66600
rect 0 63600 200 65000
rect 0 62000 200 63400
rect 0 60400 200 61800
rect 0 58800 200 60200
rect 0 57200 200 58600
rect 0 55600 200 57000
rect 0 54000 200 55400
rect 0 52400 200 53800
rect 0 50800 200 52200
rect 0 49200 200 50600
rect 0 46000 200 49000
rect 0 42800 200 45800
rect 0 41200 200 42600
rect 0 39600 200 41000
rect 0 36400 200 39400
rect 0 33200 200 36200
rect 0 30000 200 33000
rect 0 26800 200 29800
rect 0 25200 200 26600
rect 0 23600 200 25000
rect 0 20400 200 23400
rect 0 17200 200 20200
rect 0 14000 200 17000
rect 1800 68400 2000 69678
rect 1800 66800 2000 68200
rect 1800 65200 2000 66600
rect 1800 63600 2000 65000
rect 1800 62000 2000 63400
rect 1800 60400 2000 61800
rect 1800 58800 2000 60200
rect 1800 57200 2000 58600
rect 1800 55600 2000 57000
rect 1800 54000 2000 55400
rect 1800 52400 2000 53800
rect 1800 50800 2000 52200
rect 1800 49200 2000 50600
rect 1800 46000 2000 49000
rect 1800 42800 2000 45800
rect 1800 41200 2000 42600
rect 1800 39600 2000 41000
rect 1800 36400 2000 39400
rect 1800 33200 2000 36200
rect 1800 30000 2000 33000
rect 1800 26800 2000 29800
rect 1800 25200 2000 26600
rect 1800 23600 2000 25000
rect 1800 20400 2000 23400
rect 1800 17200 2000 20200
rect 1800 14000 2000 17000
<< obsm5 >>
rect 300 14000 1700 69678
<< labels >>
rlabel metal5 s 1800 26800 2000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 30000 2000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 33200 2000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 36400 2000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 42800 2000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 23600 2000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 41200 2000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 52400 2000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 54000 2000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 55600 2000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 58800 2000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 66800 2000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 26800 2000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 30000 2000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 33200 2000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 36400 2000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 42800 2000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 23600 2000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 41200 2000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 52400 2000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 54000 2000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 55600 2000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 58800 2000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 1800 66800 2000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 26800 2000 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 30000 2000 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 33200 2000 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 36400 2000 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 42800 2000 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 23600 2000 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 41200 2000 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 52400 2000 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 54000 2000 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 55600 2000 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 58800 2000 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 1800 66800 2000 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 66800 200 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 58800 200 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 55600 200 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 54000 200 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 52400 200 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 42800 200 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 41200 200 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 36400 200 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 33200 200 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 30000 200 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 26800 200 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 66800 200 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 58800 200 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 55600 200 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 54000 200 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 52400 200 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 42800 200 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 41200 200 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 36400 200 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 33200 200 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 30000 200 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 26800 200 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 66800 200 68200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 58800 200 60200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 55600 200 57000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 54000 200 55400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 52400 200 53800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 42800 200 45800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 41200 200 42600 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 36400 200 39400 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 33200 200 36200 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 30000 200 33000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 26800 200 29800 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 0 23600 200 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 23600 200 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 23600 200 25000 6 DVDD
port 1 nsew power bidirectional
rlabel metal5 s 1800 14000 2000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 1800 17200 2000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 1800 20400 2000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 1800 46000 2000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 1800 25200 2000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 1800 39600 2000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 1800 57200 2000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 1800 60400 2000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 1800 65200 2000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 1800 68400 2000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 1800 14000 2000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 1800 17200 2000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 1800 20400 2000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 1800 46000 2000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 1800 25200 2000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 1800 39600 2000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 1800 57200 2000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 1800 60400 2000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 1800 65200 2000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 1800 68400 2000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 1800 14000 2000 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 1800 17200 2000 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 1800 20400 2000 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 1800 46000 2000 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 1800 25200 2000 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 1800 39600 2000 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 1800 57200 2000 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 1800 60400 2000 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 1800 65200 2000 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 1800 68400 2000 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 68400 200 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 65200 200 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 60400 200 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 57200 200 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 46000 200 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 39600 200 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 25200 200 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 20400 200 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 17200 200 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 68400 200 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 65200 200 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 60400 200 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 57200 200 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 46000 200 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 39600 200 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 25200 200 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 20400 200 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 17200 200 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 68400 200 69678 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 65200 200 66600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 60400 200 61800 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 57200 200 58600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 46000 200 49000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 39600 200 41000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 25200 200 26600 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 20400 200 23400 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 17200 200 20200 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 0 14000 200 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 14000 200 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 14000 200 17000 6 DVSS
port 2 nsew ground bidirectional
rlabel metal5 s 1800 50800 2000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 1800 62000 2000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 1800 50800 2000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 1800 62000 2000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 1800 50800 2000 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 1800 62000 2000 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 62000 200 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 62000 200 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 0 62000 200 63400 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 0 50800 200 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 50800 200 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 50800 200 52200 6 VDD
port 3 nsew power bidirectional
rlabel metal5 s 1800 49200 2000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 1800 63600 2000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 1800 49200 2000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 1800 63600 2000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 1800 49200 2000 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 1800 63600 2000 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 63600 200 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 0 63600 200 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 63600 200 65000 6 VSS
port 4 nsew ground bidirectional
rlabel metal5 s 0 49200 200 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 0 49200 200 50600 6 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 49200 200 50600 6 VSS
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 2000 70000
string LEFclass PAD SPACER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 17619454
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17612986
<< end >>
