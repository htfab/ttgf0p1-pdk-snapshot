magic
tech gf180mcuD
magscale 1 5
timestamp 1755005639
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_0
timestamp 1755005639
transform -1 0 10200 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_1
timestamp 1755005639
transform -1 0 9900 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_2
timestamp 1755005639
transform -1 0 9600 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_3
timestamp 1755005639
transform -1 0 9300 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_4
timestamp 1755005639
transform -1 0 9000 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_5
timestamp 1755005639
transform -1 0 8700 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_6
timestamp 1755005639
transform -1 0 10800 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_7
timestamp 1755005639
transform -1 0 10500 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_8
timestamp 1755005639
transform -1 0 10200 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_9
timestamp 1755005639
transform -1 0 9900 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_10
timestamp 1755005639
transform -1 0 9600 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_11
timestamp 1755005639
transform -1 0 9300 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_12
timestamp 1755005639
transform -1 0 9000 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_13
timestamp 1755005639
transform -1 0 10800 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_14
timestamp 1755005639
transform -1 0 8700 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_15
timestamp 1755005639
transform -1 0 10800 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_16
timestamp 1755005639
transform -1 0 10500 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_17
timestamp 1755005639
transform -1 0 10200 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_18
timestamp 1755005639
transform -1 0 9900 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_19
timestamp 1755005639
transform -1 0 9600 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_20
timestamp 1755005639
transform -1 0 9300 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_21
timestamp 1755005639
transform -1 0 9000 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_22
timestamp 1755005639
transform -1 0 8700 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_23
timestamp 1755005639
transform -1 0 10500 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_24
timestamp 1755005639
transform 1 0 6600 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_25
timestamp 1755005639
transform 1 0 6900 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_26
timestamp 1755005639
transform 1 0 7200 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_27
timestamp 1755005639
transform 1 0 7500 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_28
timestamp 1755005639
transform 1 0 7800 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_29
timestamp 1755005639
transform 1 0 5700 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_30
timestamp 1755005639
transform 1 0 6300 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_31
timestamp 1755005639
transform 1 0 6600 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_32
timestamp 1755005639
transform 1 0 6900 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_33
timestamp 1755005639
transform 1 0 7200 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_34
timestamp 1755005639
transform 1 0 7500 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_35
timestamp 1755005639
transform 1 0 7800 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_36
timestamp 1755005639
transform 1 0 6000 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_37
timestamp 1755005639
transform 1 0 5700 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_38
timestamp 1755005639
transform 1 0 6000 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_39
timestamp 1755005639
transform 1 0 6300 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_40
timestamp 1755005639
transform 1 0 6600 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_41
timestamp 1755005639
transform 1 0 6900 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_42
timestamp 1755005639
transform 1 0 7200 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_43
timestamp 1755005639
transform 1 0 7500 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_44
timestamp 1755005639
transform 1 0 7800 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_45
timestamp 1755005639
transform 1 0 5700 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_46
timestamp 1755005639
transform 1 0 6000 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_47
timestamp 1755005639
transform 1 0 6300 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_48
timestamp 1755005639
transform 1 0 5700 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_49
timestamp 1755005639
transform 1 0 6000 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_50
timestamp 1755005639
transform 1 0 6300 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_51
timestamp 1755005639
transform 1 0 6600 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_52
timestamp 1755005639
transform 1 0 6300 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_53
timestamp 1755005639
transform 1 0 6600 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_54
timestamp 1755005639
transform 1 0 6900 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_55
timestamp 1755005639
transform 1 0 7200 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_56
timestamp 1755005639
transform 1 0 7500 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_57
timestamp 1755005639
transform 1 0 7800 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_58
timestamp 1755005639
transform 1 0 6900 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_59
timestamp 1755005639
transform 1 0 7200 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_60
timestamp 1755005639
transform 1 0 7500 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_61
timestamp 1755005639
transform 1 0 7800 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_62
timestamp 1755005639
transform 1 0 5700 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_63
timestamp 1755005639
transform 1 0 6000 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_64
timestamp 1755005639
transform -1 0 9300 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_65
timestamp 1755005639
transform -1 0 9900 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_66
timestamp 1755005639
transform -1 0 9000 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_67
timestamp 1755005639
transform -1 0 8700 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_68
timestamp 1755005639
transform -1 0 9600 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_69
timestamp 1755005639
transform -1 0 10800 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_70
timestamp 1755005639
transform -1 0 10500 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_71
timestamp 1755005639
transform -1 0 10200 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_72
timestamp 1755005639
transform -1 0 9900 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_73
timestamp 1755005639
transform -1 0 9600 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_74
timestamp 1755005639
transform -1 0 9300 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_75
timestamp 1755005639
transform -1 0 9000 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_76
timestamp 1755005639
transform -1 0 8700 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_77
timestamp 1755005639
transform -1 0 10800 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_78
timestamp 1755005639
transform -1 0 10500 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_79
timestamp 1755005639
transform -1 0 10200 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_80
timestamp 1755005639
transform 1 0 5700 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_81
timestamp 1755005639
transform 1 0 6000 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_82
timestamp 1755005639
transform 1 0 6300 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_83
timestamp 1755005639
transform 1 0 6600 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_84
timestamp 1755005639
transform 1 0 6900 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_85
timestamp 1755005639
transform 1 0 7200 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_86
timestamp 1755005639
transform 1 0 7500 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_87
timestamp 1755005639
transform 1 0 7800 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_88
timestamp 1755005639
transform 1 0 5700 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_89
timestamp 1755005639
transform 1 0 6000 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_90
timestamp 1755005639
transform 1 0 6300 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_91
timestamp 1755005639
transform 1 0 6600 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_92
timestamp 1755005639
transform 1 0 6900 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_93
timestamp 1755005639
transform 1 0 7200 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_94
timestamp 1755005639
transform 1 0 7500 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_95
timestamp 1755005639
transform 1 0 7800 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_96
timestamp 1755005639
transform -1 0 10800 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_97
timestamp 1755005639
transform -1 0 10500 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_98
timestamp 1755005639
transform -1 0 10200 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_99
timestamp 1755005639
transform -1 0 9900 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_100
timestamp 1755005639
transform -1 0 9600 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_101
timestamp 1755005639
transform -1 0 9300 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_102
timestamp 1755005639
transform -1 0 9000 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_103
timestamp 1755005639
transform -1 0 8700 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_104
timestamp 1755005639
transform -1 0 10800 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_105
timestamp 1755005639
transform -1 0 10500 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_106
timestamp 1755005639
transform -1 0 10200 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_107
timestamp 1755005639
transform -1 0 9900 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_108
timestamp 1755005639
transform -1 0 9600 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_109
timestamp 1755005639
transform -1 0 9300 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_110
timestamp 1755005639
transform -1 0 9000 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_111
timestamp 1755005639
transform -1 0 8700 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_112
timestamp 1755005639
transform -1 0 3600 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_113
timestamp 1755005639
transform -1 0 3300 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_114
timestamp 1755005639
transform -1 0 5400 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_115
timestamp 1755005639
transform -1 0 5100 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_116
timestamp 1755005639
transform -1 0 4800 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_117
timestamp 1755005639
transform -1 0 4500 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_118
timestamp 1755005639
transform -1 0 4200 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_119
timestamp 1755005639
transform -1 0 3900 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_120
timestamp 1755005639
transform -1 0 3600 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_121
timestamp 1755005639
transform -1 0 3300 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_122
timestamp 1755005639
transform -1 0 5100 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_123
timestamp 1755005639
transform -1 0 4800 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_124
timestamp 1755005639
transform -1 0 4500 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_125
timestamp 1755005639
transform -1 0 4200 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_126
timestamp 1755005639
transform -1 0 3900 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_127
timestamp 1755005639
transform -1 0 3600 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_128
timestamp 1755005639
transform -1 0 3300 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_129
timestamp 1755005639
transform -1 0 5400 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_130
timestamp 1755005639
transform -1 0 5100 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_131
timestamp 1755005639
transform -1 0 4800 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_132
timestamp 1755005639
transform -1 0 4500 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_133
timestamp 1755005639
transform -1 0 4200 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_134
timestamp 1755005639
transform -1 0 3900 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_135
timestamp 1755005639
transform -1 0 5400 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_136
timestamp 1755005639
transform 1 0 1200 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_137
timestamp 1755005639
transform 1 0 900 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_138
timestamp 1755005639
transform 1 0 600 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_139
timestamp 1755005639
transform 1 0 1500 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_140
timestamp 1755005639
transform 1 0 300 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_141
timestamp 1755005639
transform 1 0 1200 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_142
timestamp 1755005639
transform 1 0 900 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_143
timestamp 1755005639
transform 1 0 600 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_144
timestamp 1755005639
transform 1 0 2400 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_145
timestamp 1755005639
transform 1 0 2100 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_146
timestamp 1755005639
transform 1 0 1800 0 1 900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_147
timestamp 1755005639
transform 1 0 1500 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_148
timestamp 1755005639
transform 1 0 300 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_149
timestamp 1755005639
transform 1 0 2100 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_150
timestamp 1755005639
transform 1 0 600 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_151
timestamp 1755005639
transform 1 0 2400 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_152
timestamp 1755005639
transform 1 0 2100 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_153
timestamp 1755005639
transform 1 0 1800 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_154
timestamp 1755005639
transform 1 0 1200 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_155
timestamp 1755005639
transform 1 0 900 0 1 0
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_156
timestamp 1755005639
transform 1 0 2400 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_157
timestamp 1755005639
transform 1 0 1800 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_158
timestamp 1755005639
transform 1 0 1500 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_159
timestamp 1755005639
transform 1 0 300 0 1 1800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_160
timestamp 1755005639
transform 1 0 600 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_161
timestamp 1755005639
transform 1 0 900 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_162
timestamp 1755005639
transform 1 0 1200 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_163
timestamp 1755005639
transform 1 0 1500 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_164
timestamp 1755005639
transform 1 0 1800 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_165
timestamp 1755005639
transform 1 0 2100 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_166
timestamp 1755005639
transform 1 0 2400 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_167
timestamp 1755005639
transform 1 0 300 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_168
timestamp 1755005639
transform 1 0 600 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_169
timestamp 1755005639
transform 1 0 900 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_170
timestamp 1755005639
transform 1 0 1200 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_171
timestamp 1755005639
transform 1 0 1500 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_172
timestamp 1755005639
transform 1 0 1800 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_173
timestamp 1755005639
transform 1 0 2100 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_174
timestamp 1755005639
transform 1 0 2400 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_175
timestamp 1755005639
transform 1 0 300 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_176
timestamp 1755005639
transform -1 0 4200 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_177
timestamp 1755005639
transform -1 0 3900 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_178
timestamp 1755005639
transform -1 0 3600 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_179
timestamp 1755005639
transform -1 0 3300 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_180
timestamp 1755005639
transform -1 0 5400 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_181
timestamp 1755005639
transform -1 0 5100 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_182
timestamp 1755005639
transform -1 0 4800 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_183
timestamp 1755005639
transform -1 0 4500 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_184
timestamp 1755005639
transform -1 0 4200 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_185
timestamp 1755005639
transform -1 0 3900 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_186
timestamp 1755005639
transform -1 0 3600 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_187
timestamp 1755005639
transform -1 0 3300 0 1 5400
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_188
timestamp 1755005639
transform -1 0 5400 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_189
timestamp 1755005639
transform -1 0 5100 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_190
timestamp 1755005639
transform -1 0 4800 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_191
timestamp 1755005639
transform -1 0 4500 0 1 4500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_192
timestamp 1755005639
transform 1 0 300 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_193
timestamp 1755005639
transform 1 0 600 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_194
timestamp 1755005639
transform 1 0 900 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_195
timestamp 1755005639
transform -1 0 5400 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_196
timestamp 1755005639
transform -1 0 5100 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_197
timestamp 1755005639
transform -1 0 4800 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_198
timestamp 1755005639
transform -1 0 4500 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_199
timestamp 1755005639
transform -1 0 4200 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_200
timestamp 1755005639
transform -1 0 3900 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_201
timestamp 1755005639
transform -1 0 3600 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_202
timestamp 1755005639
transform -1 0 3300 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_203
timestamp 1755005639
transform -1 0 5400 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_204
timestamp 1755005639
transform -1 0 5100 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_205
timestamp 1755005639
transform -1 0 4800 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_206
timestamp 1755005639
transform -1 0 4500 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_207
timestamp 1755005639
transform -1 0 4200 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_208
timestamp 1755005639
transform -1 0 3900 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_209
timestamp 1755005639
transform -1 0 3600 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_210
timestamp 1755005639
transform -1 0 3300 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_211
timestamp 1755005639
transform 1 0 1200 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_212
timestamp 1755005639
transform 1 0 1500 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_213
timestamp 1755005639
transform 1 0 1800 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_214
timestamp 1755005639
transform 1 0 2100 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_215
timestamp 1755005639
transform 1 0 2400 0 1 2700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_216
timestamp 1755005639
transform 1 0 300 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_217
timestamp 1755005639
transform 1 0 600 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_218
timestamp 1755005639
transform 1 0 900 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_219
timestamp 1755005639
transform 1 0 1200 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_220
timestamp 1755005639
transform 1 0 1500 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_221
timestamp 1755005639
transform 1 0 1800 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_222
timestamp 1755005639
transform 1 0 2100 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_223
timestamp 1755005639
transform 1 0 2400 0 1 3600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_224
timestamp 1755005639
transform -1 0 3900 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_225
timestamp 1755005639
transform -1 0 3600 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_226
timestamp 1755005639
transform -1 0 3300 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_227
timestamp 1755005639
transform -1 0 5400 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_228
timestamp 1755005639
transform -1 0 5100 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_229
timestamp 1755005639
transform -1 0 4800 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_230
timestamp 1755005639
transform -1 0 4500 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_231
timestamp 1755005639
transform -1 0 4200 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_232
timestamp 1755005639
transform -1 0 3900 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_233
timestamp 1755005639
transform -1 0 3600 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_234
timestamp 1755005639
transform -1 0 3300 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_235
timestamp 1755005639
transform -1 0 5400 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_236
timestamp 1755005639
transform -1 0 5100 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_237
timestamp 1755005639
transform -1 0 4800 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_238
timestamp 1755005639
transform -1 0 4500 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_239
timestamp 1755005639
transform -1 0 4200 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_240
timestamp 1755005639
transform 1 0 1200 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_241
timestamp 1755005639
transform 1 0 1500 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_242
timestamp 1755005639
transform 1 0 1800 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_243
timestamp 1755005639
transform 1 0 2100 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_244
timestamp 1755005639
transform 1 0 2400 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_245
timestamp 1755005639
transform 1 0 300 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_246
timestamp 1755005639
transform 1 0 600 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_247
timestamp 1755005639
transform 1 0 900 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_248
timestamp 1755005639
transform 1 0 300 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_249
timestamp 1755005639
transform 1 0 600 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_250
timestamp 1755005639
transform 1 0 900 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_251
timestamp 1755005639
transform 1 0 1200 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_252
timestamp 1755005639
transform 1 0 1500 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_253
timestamp 1755005639
transform 1 0 1800 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_254
timestamp 1755005639
transform 1 0 2100 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_255
timestamp 1755005639
transform 1 0 2400 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_256
timestamp 1755005639
transform 1 0 1200 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_257
timestamp 1755005639
transform 1 0 1500 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_258
timestamp 1755005639
transform 1 0 1800 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_259
timestamp 1755005639
transform 1 0 2100 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_260
timestamp 1755005639
transform 1 0 2400 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_261
timestamp 1755005639
transform 1 0 300 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_262
timestamp 1755005639
transform 1 0 600 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_263
timestamp 1755005639
transform 1 0 900 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_264
timestamp 1755005639
transform 1 0 1200 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_265
timestamp 1755005639
transform 1 0 1500 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_266
timestamp 1755005639
transform 1 0 1800 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_267
timestamp 1755005639
transform 1 0 2100 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_268
timestamp 1755005639
transform 1 0 2400 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_269
timestamp 1755005639
transform 1 0 300 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_270
timestamp 1755005639
transform 1 0 600 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_271
timestamp 1755005639
transform 1 0 900 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_272
timestamp 1755005639
transform 1 0 1200 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_273
timestamp 1755005639
transform 1 0 1500 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_274
timestamp 1755005639
transform 1 0 2400 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_275
timestamp 1755005639
transform 1 0 900 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_276
timestamp 1755005639
transform 1 0 300 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_277
timestamp 1755005639
transform 1 0 600 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_278
timestamp 1755005639
transform 1 0 1800 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_279
timestamp 1755005639
transform 1 0 2100 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_280
timestamp 1755005639
transform -1 0 3300 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_281
timestamp 1755005639
transform -1 0 5400 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_282
timestamp 1755005639
transform -1 0 5100 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_283
timestamp 1755005639
transform -1 0 4800 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_284
timestamp 1755005639
transform -1 0 4500 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_285
timestamp 1755005639
transform -1 0 4200 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_286
timestamp 1755005639
transform -1 0 3900 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_287
timestamp 1755005639
transform -1 0 3600 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_288
timestamp 1755005639
transform -1 0 3300 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_289
timestamp 1755005639
transform -1 0 5400 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_290
timestamp 1755005639
transform -1 0 5100 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_291
timestamp 1755005639
transform -1 0 4800 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_292
timestamp 1755005639
transform -1 0 4500 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_293
timestamp 1755005639
transform -1 0 4200 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_294
timestamp 1755005639
transform -1 0 3900 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_295
timestamp 1755005639
transform -1 0 3600 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_296
timestamp 1755005639
transform -1 0 3300 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_297
timestamp 1755005639
transform -1 0 5400 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_298
timestamp 1755005639
transform -1 0 5100 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_299
timestamp 1755005639
transform -1 0 4800 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_300
timestamp 1755005639
transform -1 0 4500 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_301
timestamp 1755005639
transform -1 0 4200 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_302
timestamp 1755005639
transform -1 0 3900 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_303
timestamp 1755005639
transform -1 0 3600 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_304
timestamp 1755005639
transform 1 0 300 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_305
timestamp 1755005639
transform 1 0 600 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_306
timestamp 1755005639
transform 1 0 900 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_307
timestamp 1755005639
transform 1 0 1200 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_308
timestamp 1755005639
transform 1 0 1500 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_309
timestamp 1755005639
transform 1 0 1800 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_310
timestamp 1755005639
transform 1 0 2100 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_311
timestamp 1755005639
transform 1 0 2400 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_312
timestamp 1755005639
transform -1 0 5400 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_313
timestamp 1755005639
transform -1 0 5100 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_314
timestamp 1755005639
transform -1 0 4800 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_315
timestamp 1755005639
transform -1 0 4500 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_316
timestamp 1755005639
transform -1 0 4200 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_317
timestamp 1755005639
transform -1 0 3900 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_318
timestamp 1755005639
transform -1 0 3600 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_319
timestamp 1755005639
transform -1 0 3300 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_320
timestamp 1755005639
transform -1 0 5400 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_321
timestamp 1755005639
transform -1 0 5100 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_322
timestamp 1755005639
transform -1 0 4800 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_323
timestamp 1755005639
transform -1 0 4500 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_324
timestamp 1755005639
transform -1 0 4200 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_325
timestamp 1755005639
transform -1 0 3900 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_326
timestamp 1755005639
transform -1 0 3600 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_327
timestamp 1755005639
transform -1 0 3300 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_328
timestamp 1755005639
transform 1 0 300 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_329
timestamp 1755005639
transform 1 0 600 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_330
timestamp 1755005639
transform 1 0 900 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_331
timestamp 1755005639
transform 1 0 1200 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_332
timestamp 1755005639
transform 1 0 1500 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_333
timestamp 1755005639
transform 1 0 1800 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_334
timestamp 1755005639
transform 1 0 2100 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_335
timestamp 1755005639
transform 1 0 2400 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_336
timestamp 1755005639
transform -1 0 8700 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_337
timestamp 1755005639
transform -1 0 10800 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_338
timestamp 1755005639
transform -1 0 10500 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_339
timestamp 1755005639
transform -1 0 10200 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_340
timestamp 1755005639
transform -1 0 9900 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_341
timestamp 1755005639
transform -1 0 9600 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_342
timestamp 1755005639
transform -1 0 9300 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_343
timestamp 1755005639
transform -1 0 9000 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_344
timestamp 1755005639
transform -1 0 8700 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_345
timestamp 1755005639
transform -1 0 10800 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_346
timestamp 1755005639
transform -1 0 10500 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_347
timestamp 1755005639
transform -1 0 10200 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_348
timestamp 1755005639
transform -1 0 9900 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_349
timestamp 1755005639
transform -1 0 9600 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_350
timestamp 1755005639
transform -1 0 9300 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_351
timestamp 1755005639
transform -1 0 9000 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_352
timestamp 1755005639
transform 1 0 6900 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_353
timestamp 1755005639
transform 1 0 7200 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_354
timestamp 1755005639
transform 1 0 7500 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_355
timestamp 1755005639
transform 1 0 7800 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_356
timestamp 1755005639
transform 1 0 5700 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_357
timestamp 1755005639
transform 1 0 6000 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_358
timestamp 1755005639
transform 1 0 6300 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_359
timestamp 1755005639
transform 1 0 6600 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_360
timestamp 1755005639
transform 1 0 6900 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_361
timestamp 1755005639
transform 1 0 7200 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_362
timestamp 1755005639
transform 1 0 7500 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_363
timestamp 1755005639
transform 1 0 7800 0 1 9000
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_364
timestamp 1755005639
transform 1 0 5700 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_365
timestamp 1755005639
transform 1 0 6000 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_366
timestamp 1755005639
transform 1 0 6300 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_367
timestamp 1755005639
transform 1 0 6600 0 1 8100
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_368
timestamp 1755005639
transform 1 0 5700 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_369
timestamp 1755005639
transform 1 0 6000 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_370
timestamp 1755005639
transform 1 0 6300 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_371
timestamp 1755005639
transform 1 0 6600 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_372
timestamp 1755005639
transform 1 0 6900 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_373
timestamp 1755005639
transform 1 0 7200 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_374
timestamp 1755005639
transform 1 0 7500 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_375
timestamp 1755005639
transform 1 0 7800 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_376
timestamp 1755005639
transform 1 0 5700 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_377
timestamp 1755005639
transform 1 0 6000 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_378
timestamp 1755005639
transform 1 0 6300 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_379
timestamp 1755005639
transform 1 0 6600 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_380
timestamp 1755005639
transform 1 0 6900 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_381
timestamp 1755005639
transform 1 0 7200 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_382
timestamp 1755005639
transform 1 0 7500 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_383
timestamp 1755005639
transform 1 0 7800 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_384
timestamp 1755005639
transform 1 0 6900 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_385
timestamp 1755005639
transform 1 0 7200 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_386
timestamp 1755005639
transform 1 0 7500 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_387
timestamp 1755005639
transform 1 0 7800 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_388
timestamp 1755005639
transform 1 0 5700 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_389
timestamp 1755005639
transform 1 0 6000 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_390
timestamp 1755005639
transform 1 0 6300 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_391
timestamp 1755005639
transform 1 0 6600 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_392
timestamp 1755005639
transform -1 0 10800 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_393
timestamp 1755005639
transform -1 0 10500 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_394
timestamp 1755005639
transform -1 0 10200 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_395
timestamp 1755005639
transform -1 0 9900 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_396
timestamp 1755005639
transform -1 0 9600 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_397
timestamp 1755005639
transform -1 0 9300 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_398
timestamp 1755005639
transform -1 0 9000 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_399
timestamp 1755005639
transform -1 0 8700 0 1 12600
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_400
timestamp 1755005639
transform -1 0 10800 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_401
timestamp 1755005639
transform -1 0 10500 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_402
timestamp 1755005639
transform -1 0 10200 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_403
timestamp 1755005639
transform -1 0 9900 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_404
timestamp 1755005639
transform -1 0 9600 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_405
timestamp 1755005639
transform -1 0 9300 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_406
timestamp 1755005639
transform -1 0 9000 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_407
timestamp 1755005639
transform -1 0 8700 0 1 13500
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_408
timestamp 1755005639
transform -1 0 10800 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_409
timestamp 1755005639
transform -1 0 10500 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_410
timestamp 1755005639
transform -1 0 10200 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_411
timestamp 1755005639
transform -1 0 9900 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_412
timestamp 1755005639
transform -1 0 9600 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_413
timestamp 1755005639
transform -1 0 9300 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_414
timestamp 1755005639
transform -1 0 9000 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_415
timestamp 1755005639
transform -1 0 8700 0 1 11700
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_416
timestamp 1755005639
transform 1 0 5700 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_417
timestamp 1755005639
transform 1 0 6000 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_418
timestamp 1755005639
transform 1 0 6300 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_419
timestamp 1755005639
transform 1 0 6600 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_420
timestamp 1755005639
transform 1 0 6900 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_421
timestamp 1755005639
transform 1 0 7200 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_422
timestamp 1755005639
transform 1 0 7500 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_423
timestamp 1755005639
transform 1 0 7800 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_424
timestamp 1755005639
transform 1 0 5700 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_425
timestamp 1755005639
transform 1 0 6000 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_426
timestamp 1755005639
transform 1 0 6300 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_427
timestamp 1755005639
transform 1 0 6600 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_428
timestamp 1755005639
transform 1 0 6900 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_429
timestamp 1755005639
transform 1 0 7200 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_430
timestamp 1755005639
transform 1 0 7500 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_431
timestamp 1755005639
transform -1 0 10800 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_432
timestamp 1755005639
transform -1 0 10500 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_433
timestamp 1755005639
transform -1 0 10200 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_434
timestamp 1755005639
transform -1 0 9900 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_435
timestamp 1755005639
transform -1 0 9600 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_436
timestamp 1755005639
transform -1 0 9300 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_437
timestamp 1755005639
transform -1 0 9000 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_438
timestamp 1755005639
transform -1 0 8700 0 1 9900
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_439
timestamp 1755005639
transform -1 0 10800 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_440
timestamp 1755005639
transform -1 0 10500 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_441
timestamp 1755005639
transform -1 0 10200 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_442
timestamp 1755005639
transform -1 0 9900 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_443
timestamp 1755005639
transform -1 0 9600 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_444
timestamp 1755005639
transform -1 0 9300 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_445
timestamp 1755005639
transform -1 0 9000 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_446
timestamp 1755005639
transform -1 0 8700 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_447
timestamp 1755005639
transform 1 0 7800 0 1 10800
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_448
timestamp 1755005639
transform -1 0 5400 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_449
timestamp 1755005639
transform -1 0 5100 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_450
timestamp 1755005639
transform -1 0 4800 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_451
timestamp 1755005639
transform -1 0 4500 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_452
timestamp 1755005639
transform -1 0 4200 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_453
timestamp 1755005639
transform -1 0 3900 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_454
timestamp 1755005639
transform -1 0 3600 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_455
timestamp 1755005639
transform -1 0 3300 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_456
timestamp 1755005639
transform -1 0 5400 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_457
timestamp 1755005639
transform -1 0 5100 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_458
timestamp 1755005639
transform -1 0 4800 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_459
timestamp 1755005639
transform -1 0 4500 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_460
timestamp 1755005639
transform -1 0 4200 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_461
timestamp 1755005639
transform -1 0 3900 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_462
timestamp 1755005639
transform -1 0 3600 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_463
timestamp 1755005639
transform -1 0 3300 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_464
timestamp 1755005639
transform -1 0 10800 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_465
timestamp 1755005639
transform -1 0 10500 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_466
timestamp 1755005639
transform -1 0 10200 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_467
timestamp 1755005639
transform -1 0 9900 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_468
timestamp 1755005639
transform -1 0 9600 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_469
timestamp 1755005639
transform -1 0 9300 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_470
timestamp 1755005639
transform -1 0 9000 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_471
timestamp 1755005639
transform -1 0 8700 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_472
timestamp 1755005639
transform -1 0 10800 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_473
timestamp 1755005639
transform -1 0 10500 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_474
timestamp 1755005639
transform -1 0 10200 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_475
timestamp 1755005639
transform -1 0 9900 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_476
timestamp 1755005639
transform -1 0 9600 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_477
timestamp 1755005639
transform -1 0 9300 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_478
timestamp 1755005639
transform -1 0 9000 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_479
timestamp 1755005639
transform -1 0 8700 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_480
timestamp 1755005639
transform 1 0 300 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_481
timestamp 1755005639
transform 1 0 600 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_482
timestamp 1755005639
transform 1 0 900 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_483
timestamp 1755005639
transform 1 0 1200 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_484
timestamp 1755005639
transform 1 0 1500 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_485
timestamp 1755005639
transform 1 0 1800 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_486
timestamp 1755005639
transform 1 0 2100 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_487
timestamp 1755005639
transform 1 0 2400 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_488
timestamp 1755005639
transform 1 0 300 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_489
timestamp 1755005639
transform 1 0 600 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_490
timestamp 1755005639
transform 1 0 900 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_491
timestamp 1755005639
transform 1 0 1200 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_492
timestamp 1755005639
transform 1 0 1500 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_493
timestamp 1755005639
transform 1 0 1800 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_494
timestamp 1755005639
transform 1 0 2100 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_495
timestamp 1755005639
transform 1 0 2400 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_496
timestamp 1755005639
transform 1 0 5700 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_497
timestamp 1755005639
transform 1 0 6000 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_498
timestamp 1755005639
transform 1 0 6300 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_499
timestamp 1755005639
transform 1 0 6600 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_500
timestamp 1755005639
transform 1 0 6900 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_501
timestamp 1755005639
transform 1 0 7200 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_502
timestamp 1755005639
transform 1 0 7500 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_503
timestamp 1755005639
transform 1 0 7800 0 1 6300
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_504
timestamp 1755005639
transform 1 0 5700 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_505
timestamp 1755005639
transform 1 0 6000 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_506
timestamp 1755005639
transform 1 0 6300 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_507
timestamp 1755005639
transform 1 0 6600 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_508
timestamp 1755005639
transform 1 0 6900 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_509
timestamp 1755005639
transform 1 0 7200 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_510
timestamp 1755005639
transform 1 0 7500 0 1 7200
box -34 -34 334 934
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_511
timestamp 1755005639
transform 1 0 7800 0 1 7200
box -34 -34 334 934
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_0
timestamp 1755005639
transform -1 0 8400 0 1 450
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_1
timestamp 1755005639
transform -1 0 8400 0 1 1350
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_2
timestamp 1755005639
transform -1 0 8400 0 1 2250
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_3
timestamp 1755005639
transform -1 0 8400 0 1 3150
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_4
timestamp 1755005639
transform -1 0 8400 0 1 4050
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_5
timestamp 1755005639
transform -1 0 8400 0 1 4950
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_6
timestamp 1755005639
transform -1 0 8400 0 1 5850
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_7
timestamp 1755005639
transform -1 0 300 0 1 450
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_8
timestamp 1755005639
transform -1 0 300 0 1 1350
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_9
timestamp 1755005639
transform -1 0 300 0 1 2250
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_10
timestamp 1755005639
transform -1 0 300 0 1 5850
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_11
timestamp 1755005639
transform -1 0 300 0 1 4950
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_12
timestamp 1755005639
transform -1 0 3000 0 1 1350
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_13
timestamp 1755005639
transform -1 0 3000 0 1 2250
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_14
timestamp 1755005639
transform -1 0 3000 0 1 3150
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_15
timestamp 1755005639
transform -1 0 3000 0 1 4050
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_16
timestamp 1755005639
transform -1 0 3000 0 1 4950
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_17
timestamp 1755005639
transform -1 0 3000 0 1 5850
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_18
timestamp 1755005639
transform -1 0 300 0 1 3150
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_19
timestamp 1755005639
transform -1 0 300 0 1 4050
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_20
timestamp 1755005639
transform -1 0 3000 0 1 450
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_21
timestamp 1755005639
transform -1 0 300 0 1 8550
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_22
timestamp 1755005639
transform -1 0 300 0 1 9450
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_23
timestamp 1755005639
transform -1 0 300 0 1 12150
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_24
timestamp 1755005639
transform -1 0 300 0 1 13050
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_25
timestamp 1755005639
transform -1 0 300 0 1 13950
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_26
timestamp 1755005639
transform -1 0 3000 0 1 8550
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_27
timestamp 1755005639
transform -1 0 3000 0 1 9450
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_28
timestamp 1755005639
transform -1 0 3000 0 1 10350
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_29
timestamp 1755005639
transform -1 0 3000 0 1 11250
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_30
timestamp 1755005639
transform -1 0 3000 0 1 12150
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_31
timestamp 1755005639
transform -1 0 3000 0 1 13050
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_32
timestamp 1755005639
transform -1 0 3000 0 1 13950
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_33
timestamp 1755005639
transform -1 0 300 0 1 10350
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_34
timestamp 1755005639
transform -1 0 300 0 1 11250
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_35
timestamp 1755005639
transform -1 0 8400 0 1 8550
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_36
timestamp 1755005639
transform -1 0 8400 0 1 9450
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_37
timestamp 1755005639
transform -1 0 8400 0 1 10350
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_38
timestamp 1755005639
transform -1 0 8400 0 1 11250
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_39
timestamp 1755005639
transform -1 0 8400 0 1 12150
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_40
timestamp 1755005639
transform -1 0 8400 0 1 13050
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_41
timestamp 1755005639
transform -1 0 8400 0 1 13950
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_42
timestamp 1755005639
transform -1 0 5700 0 1 450
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_43
timestamp 1755005639
transform -1 0 5700 0 1 1350
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_44
timestamp 1755005639
transform -1 0 5700 0 1 2250
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_45
timestamp 1755005639
transform -1 0 5700 0 1 3150
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_46
timestamp 1755005639
transform -1 0 5700 0 1 4050
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_47
timestamp 1755005639
transform -1 0 5700 0 1 4950
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_48
timestamp 1755005639
transform -1 0 5700 0 1 5850
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_49
timestamp 1755005639
transform -1 0 5700 0 1 6750
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_50
timestamp 1755005639
transform -1 0 5700 0 1 7650
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_51
timestamp 1755005639
transform -1 0 5700 0 1 8550
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_52
timestamp 1755005639
transform -1 0 5700 0 1 9450
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_53
timestamp 1755005639
transform -1 0 5700 0 1 10350
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_54
timestamp 1755005639
transform -1 0 5700 0 1 11250
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_55
timestamp 1755005639
transform -1 0 5700 0 1 12150
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_56
timestamp 1755005639
transform -1 0 5700 0 1 13050
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_57
timestamp 1755005639
transform -1 0 5700 0 1 13950
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_58
timestamp 1755005639
transform -1 0 3000 0 1 6750
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_59
timestamp 1755005639
transform -1 0 3000 0 1 7650
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_60
timestamp 1755005639
transform -1 0 8400 0 1 6750
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_61
timestamp 1755005639
transform -1 0 8400 0 1 7650
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_62
timestamp 1755005639
transform -1 0 300 0 1 6750
box -34 -484 334 484
use 018SRAM_strap1_2x_256x8m81  018SRAM_strap1_2x_256x8m81_63
timestamp 1755005639
transform -1 0 300 0 1 7650
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_0
timestamp 1755005639
transform 1 0 10800 0 1 450
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_1
timestamp 1755005639
transform 1 0 10800 0 1 1350
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_2
timestamp 1755005639
transform 1 0 10800 0 1 2250
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_3
timestamp 1755005639
transform 1 0 10800 0 1 4950
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_4
timestamp 1755005639
transform 1 0 10800 0 1 5850
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_5
timestamp 1755005639
transform 1 0 10800 0 1 3150
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_6
timestamp 1755005639
transform 1 0 10800 0 1 4050
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_7
timestamp 1755005639
transform 1 0 10800 0 1 8550
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_8
timestamp 1755005639
transform 1 0 10800 0 1 9450
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_9
timestamp 1755005639
transform 1 0 10800 0 1 13050
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_10
timestamp 1755005639
transform 1 0 10800 0 1 13950
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_11
timestamp 1755005639
transform 1 0 10800 0 1 12150
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_12
timestamp 1755005639
transform 1 0 10800 0 1 10350
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_13
timestamp 1755005639
transform 1 0 10800 0 1 11250
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_14
timestamp 1755005639
transform 1 0 10800 0 1 6750
box -34 -484 334 484
use 018SRAM_strap1_2x_bndry_256x8m81  018SRAM_strap1_2x_bndry_256x8m81_15
timestamp 1755005639
transform 1 0 10800 0 1 7650
box -34 -484 334 484
<< properties >>
string GDS_END 1032710
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 997250
<< end >>
