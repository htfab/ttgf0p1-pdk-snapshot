magic
tech gf180mcuD
magscale 1 10
timestamp 1753864693
<< nwell >>
rect -86 354 2998 870
<< pwell >>
rect -86 -86 2998 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 756 68 812 268
rect 916 68 972 268
rect 1076 68 1132 268
rect 1236 68 1292 268
rect 1524 68 1580 268
rect 1684 68 1740 268
rect 1844 68 1900 268
rect 2004 68 2060 268
rect 2164 68 2220 268
rect 2324 68 2380 268
rect 2484 68 2540 268
rect 2644 68 2700 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 756 440 812 716
rect 916 440 972 716
rect 1076 440 1132 716
rect 1236 440 1292 716
rect 1524 440 1580 716
rect 1684 440 1740 716
rect 1844 440 1900 716
rect 2004 440 2060 716
rect 2164 440 2220 716
rect 2324 440 2380 716
rect 2484 440 2540 716
rect 2644 440 2700 716
<< ndiff >>
rect 28 225 116 268
rect 28 179 41 225
rect 87 179 116 225
rect 28 68 116 179
rect 172 127 276 268
rect 172 81 201 127
rect 247 81 276 127
rect 172 68 276 81
rect 332 230 436 268
rect 332 184 361 230
rect 407 184 436 230
rect 332 68 436 184
rect 492 127 596 268
rect 492 81 521 127
rect 567 81 596 127
rect 492 68 596 81
rect 652 198 756 268
rect 652 152 681 198
rect 727 152 756 198
rect 652 68 756 152
rect 812 255 916 268
rect 812 209 841 255
rect 887 209 916 255
rect 812 68 916 209
rect 972 152 1076 268
rect 972 106 1001 152
rect 1047 106 1076 152
rect 972 68 1076 106
rect 1132 244 1236 268
rect 1132 198 1161 244
rect 1207 198 1236 244
rect 1132 68 1236 198
rect 1292 152 1380 268
rect 1292 106 1321 152
rect 1367 106 1380 152
rect 1292 68 1380 106
rect 1436 152 1524 268
rect 1436 106 1449 152
rect 1495 106 1524 152
rect 1436 68 1524 106
rect 1580 244 1684 268
rect 1580 198 1609 244
rect 1655 198 1684 244
rect 1580 68 1684 198
rect 1740 152 1844 268
rect 1740 106 1769 152
rect 1815 106 1844 152
rect 1740 68 1844 106
rect 1900 244 2004 268
rect 1900 198 1929 244
rect 1975 198 2004 244
rect 1900 68 2004 198
rect 2060 210 2164 268
rect 2060 164 2089 210
rect 2135 164 2164 210
rect 2060 68 2164 164
rect 2220 127 2324 268
rect 2220 81 2249 127
rect 2295 81 2324 127
rect 2220 68 2324 81
rect 2380 244 2484 268
rect 2380 198 2409 244
rect 2455 198 2484 244
rect 2380 68 2484 198
rect 2540 127 2644 268
rect 2540 81 2569 127
rect 2615 81 2644 127
rect 2540 68 2644 81
rect 2700 223 2788 268
rect 2700 177 2729 223
rect 2775 177 2788 223
rect 2700 68 2788 177
<< pdiff >>
rect 28 667 116 716
rect 28 453 41 667
rect 87 453 116 667
rect 28 440 116 453
rect 172 586 276 716
rect 172 540 201 586
rect 247 540 276 586
rect 172 440 276 540
rect 332 678 436 716
rect 332 632 361 678
rect 407 632 436 678
rect 332 440 436 632
rect 492 586 596 716
rect 492 540 521 586
rect 567 540 596 586
rect 492 440 596 540
rect 652 678 756 716
rect 652 632 681 678
rect 727 632 756 678
rect 652 440 756 632
rect 812 586 916 716
rect 812 540 841 586
rect 887 540 916 586
rect 812 440 916 540
rect 972 678 1076 716
rect 972 632 1001 678
rect 1047 632 1076 678
rect 972 440 1076 632
rect 1132 586 1236 716
rect 1132 540 1161 586
rect 1207 540 1236 586
rect 1132 440 1236 540
rect 1292 678 1524 716
rect 1292 632 1321 678
rect 1367 632 1524 678
rect 1292 586 1524 632
rect 1292 584 1415 586
rect 1292 538 1321 584
rect 1367 540 1415 584
rect 1461 540 1524 586
rect 1367 538 1524 540
rect 1292 440 1524 538
rect 1580 703 1684 716
rect 1580 657 1609 703
rect 1655 657 1684 703
rect 1580 440 1684 657
rect 1740 586 1844 716
rect 1740 540 1769 586
rect 1815 540 1844 586
rect 1740 440 1844 540
rect 1900 703 2004 716
rect 1900 657 1929 703
rect 1975 657 2004 703
rect 1900 440 2004 657
rect 2060 586 2164 716
rect 2060 540 2089 586
rect 2135 540 2164 586
rect 2060 440 2164 540
rect 2220 703 2324 716
rect 2220 657 2249 703
rect 2295 657 2324 703
rect 2220 440 2324 657
rect 2380 586 2484 716
rect 2380 540 2409 586
rect 2455 540 2484 586
rect 2380 440 2484 540
rect 2540 703 2644 716
rect 2540 657 2569 703
rect 2615 657 2644 703
rect 2540 440 2644 657
rect 2700 667 2788 716
rect 2700 458 2729 667
rect 2775 458 2788 667
rect 2700 440 2788 458
<< ndiffc >>
rect 41 179 87 225
rect 201 81 247 127
rect 361 184 407 230
rect 521 81 567 127
rect 681 152 727 198
rect 841 209 887 255
rect 1001 106 1047 152
rect 1161 198 1207 244
rect 1321 106 1367 152
rect 1449 106 1495 152
rect 1609 198 1655 244
rect 1769 106 1815 152
rect 1929 198 1975 244
rect 2089 164 2135 210
rect 2249 81 2295 127
rect 2409 198 2455 244
rect 2569 81 2615 127
rect 2729 177 2775 223
<< pdiffc >>
rect 41 453 87 667
rect 201 540 247 586
rect 361 632 407 678
rect 521 540 567 586
rect 681 632 727 678
rect 841 540 887 586
rect 1001 632 1047 678
rect 1161 540 1207 586
rect 1321 632 1367 678
rect 1321 538 1367 584
rect 1415 540 1461 586
rect 1609 657 1655 703
rect 1769 540 1815 586
rect 1929 657 1975 703
rect 2089 540 2135 586
rect 2249 657 2295 703
rect 2409 540 2455 586
rect 2569 657 2615 703
rect 2729 458 2775 667
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 756 716 812 760
rect 916 716 972 760
rect 1076 716 1132 760
rect 1236 716 1292 760
rect 1524 716 1580 760
rect 1684 716 1740 760
rect 1844 716 1900 760
rect 2004 716 2060 760
rect 2164 716 2220 760
rect 2324 716 2380 760
rect 2484 716 2540 760
rect 2644 716 2700 760
rect 116 391 172 440
rect 276 391 332 440
rect 436 391 492 440
rect 596 391 652 440
rect 98 378 652 391
rect 98 332 111 378
rect 639 332 652 378
rect 98 319 652 332
rect 116 268 172 319
rect 276 268 332 319
rect 436 268 492 319
rect 596 268 652 319
rect 756 392 812 440
rect 916 392 972 440
rect 1076 392 1132 440
rect 1236 392 1292 440
rect 756 379 1292 392
rect 756 333 933 379
rect 1279 333 1292 379
rect 756 320 1292 333
rect 756 268 812 320
rect 916 268 972 320
rect 1076 268 1132 320
rect 1236 268 1292 320
rect 1524 392 1580 440
rect 1684 392 1740 440
rect 1844 392 1900 440
rect 2004 392 2060 440
rect 1524 379 2060 392
rect 1524 333 1537 379
rect 2047 333 2060 379
rect 1524 320 2060 333
rect 1524 268 1580 320
rect 1684 268 1740 320
rect 1844 268 1900 320
rect 2004 268 2060 320
rect 2164 392 2220 440
rect 2324 392 2380 440
rect 2484 392 2540 440
rect 2644 392 2700 440
rect 2164 379 2700 392
rect 2164 333 2177 379
rect 2687 333 2700 379
rect 2164 320 2700 333
rect 2164 268 2220 320
rect 2324 268 2380 320
rect 2484 268 2540 320
rect 2644 268 2700 320
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 756 24 812 68
rect 916 24 972 68
rect 1076 24 1132 68
rect 1236 24 1292 68
rect 1524 24 1580 68
rect 1684 24 1740 68
rect 1844 24 1900 68
rect 2004 24 2060 68
rect 2164 24 2220 68
rect 2324 24 2380 68
rect 2484 24 2540 68
rect 2644 24 2700 68
<< polycontact >>
rect 111 332 639 378
rect 933 333 1279 379
rect 1537 333 2047 379
rect 2177 333 2687 379
<< metal1 >>
rect 0 724 2912 844
rect 1609 703 1655 724
rect 41 667 361 678
rect 87 632 361 667
rect 407 632 681 678
rect 727 632 1001 678
rect 1047 632 1321 678
rect 1367 632 1378 678
rect 1609 646 1655 657
rect 1929 703 1975 724
rect 1929 646 1975 657
rect 2249 703 2295 724
rect 2249 646 2295 657
rect 2569 703 2615 724
rect 2569 646 2615 657
rect 2729 667 2775 678
rect 1321 586 1367 632
rect 183 540 201 586
rect 247 540 521 586
rect 567 540 841 586
rect 887 540 1161 586
rect 1207 540 1227 586
rect 1321 584 1415 586
rect 41 440 87 453
rect 98 378 652 384
rect 98 332 111 378
rect 639 332 652 378
rect 98 325 652 332
rect 814 255 887 540
rect 1367 540 1415 584
rect 1461 540 1769 586
rect 1815 540 2089 586
rect 2135 540 2409 586
rect 2455 540 2729 586
rect 1321 527 1367 538
rect 2729 447 2775 458
rect 933 379 1292 392
rect 1279 333 1292 379
rect 933 320 1292 333
rect 1524 379 2078 385
rect 1524 333 1537 379
rect 2047 333 2078 379
rect 1524 326 2078 333
rect 2164 379 2700 385
rect 2164 333 2177 379
rect 2687 333 2700 379
rect 2164 326 2700 333
rect 41 230 87 237
rect 41 225 361 230
rect 87 184 361 225
rect 407 198 727 230
rect 814 209 841 255
rect 887 209 1161 244
rect 814 198 1161 209
rect 1207 198 1609 244
rect 1655 198 1929 244
rect 1975 198 1988 244
rect 2089 210 2409 244
rect 407 184 681 198
rect 41 148 87 179
rect 2135 198 2409 210
rect 2455 223 2775 244
rect 2455 198 2729 223
rect 2089 152 2135 164
rect 2729 159 2775 177
rect 201 127 247 138
rect 201 60 247 81
rect 521 127 567 138
rect 681 106 1001 152
rect 1047 106 1321 152
rect 1367 106 1379 152
rect 1432 106 1449 152
rect 1495 106 1769 152
rect 1815 106 2135 152
rect 2249 127 2295 138
rect 521 60 567 81
rect 2249 60 2295 81
rect 2569 127 2615 138
rect 2569 60 2615 81
rect 0 -60 2912 60
<< labels >>
flabel metal1 s 0 724 2912 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 2912 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 814 198 887 586 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 98 325 652 384 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 933 320 1292 392 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel metal1 1524 326 2078 385 0 FreeSans 200 0 0 0 C
port 8 nsew signal input
flabel metal1 2164 326 2700 385 0 FreeSans 200 0 0 0 D
port 9 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 2912 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
