magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 453 4342 1094
<< pwell >>
rect -86 -86 4342 453
<< mvnmos >>
rect 137 159 257 319
rect 497 159 617 319
rect 721 159 841 319
rect 945 159 1065 319
rect 1169 159 1289 319
rect 1393 159 1513 319
rect 1617 159 1737 319
rect 1841 159 1961 319
rect 2252 156 2372 316
rect 2476 156 2596 316
rect 2892 156 3012 316
rect 3116 156 3236 316
rect 3340 156 3460 316
rect 3564 156 3684 316
rect 3788 156 3908 316
rect 4012 156 4132 316
<< mvpmos >>
rect 157 596 257 852
rect 429 596 529 852
rect 655 596 755 852
rect 898 596 998 852
rect 1190 596 1290 852
rect 1394 596 1494 852
rect 1686 596 1786 852
rect 1890 596 1990 852
rect 2360 596 2460 852
rect 2564 596 2664 852
rect 2920 596 3020 852
rect 3136 596 3236 852
rect 3360 596 3460 852
rect 3584 596 3684 852
rect 3788 596 3888 852
rect 4012 596 4112 852
<< mvndiff >>
rect 49 303 137 319
rect 49 257 62 303
rect 108 257 137 303
rect 49 159 137 257
rect 257 303 497 319
rect 257 257 286 303
rect 332 257 497 303
rect 257 159 497 257
rect 617 303 721 319
rect 617 257 646 303
rect 692 257 721 303
rect 617 159 721 257
rect 841 303 945 319
rect 841 257 870 303
rect 916 257 945 303
rect 841 159 945 257
rect 1065 303 1169 319
rect 1065 257 1094 303
rect 1140 257 1169 303
rect 1065 159 1169 257
rect 1289 303 1393 319
rect 1289 257 1318 303
rect 1364 257 1393 303
rect 1289 159 1393 257
rect 1513 303 1617 319
rect 1513 257 1542 303
rect 1588 257 1617 303
rect 1513 159 1617 257
rect 1737 303 1841 319
rect 1737 257 1766 303
rect 1812 257 1841 303
rect 1737 159 1841 257
rect 1961 303 2049 319
rect 1961 257 1990 303
rect 2036 257 2049 303
rect 1961 159 2049 257
rect 2161 303 2252 316
rect 2161 257 2174 303
rect 2220 257 2252 303
rect 2161 156 2252 257
rect 2372 303 2476 316
rect 2372 257 2401 303
rect 2447 257 2476 303
rect 2372 156 2476 257
rect 2596 303 2684 316
rect 2596 257 2625 303
rect 2671 257 2684 303
rect 2596 156 2684 257
rect 2804 303 2892 316
rect 2804 257 2817 303
rect 2863 257 2892 303
rect 2804 156 2892 257
rect 3012 303 3116 316
rect 3012 257 3041 303
rect 3087 257 3116 303
rect 3012 156 3116 257
rect 3236 303 3340 316
rect 3236 257 3265 303
rect 3311 257 3340 303
rect 3236 156 3340 257
rect 3460 303 3564 316
rect 3460 257 3489 303
rect 3535 257 3564 303
rect 3460 156 3564 257
rect 3684 303 3788 316
rect 3684 257 3713 303
rect 3759 257 3788 303
rect 3684 156 3788 257
rect 3908 303 4012 316
rect 3908 257 3937 303
rect 3983 257 4012 303
rect 3908 156 4012 257
rect 4132 303 4220 316
rect 4132 257 4161 303
rect 4207 257 4220 303
rect 4132 156 4220 257
<< mvpdiff >>
rect 1058 871 1130 884
rect 1058 852 1071 871
rect 69 759 157 852
rect 69 619 82 759
rect 128 619 157 759
rect 69 596 157 619
rect 257 759 429 852
rect 257 619 286 759
rect 332 619 429 759
rect 257 596 429 619
rect 529 759 655 852
rect 529 619 558 759
rect 604 619 655 759
rect 529 596 655 619
rect 755 665 898 852
rect 755 619 823 665
rect 869 619 898 665
rect 755 596 898 619
rect 998 825 1071 852
rect 1117 852 1130 871
rect 1554 871 1626 884
rect 1554 852 1567 871
rect 1117 825 1190 852
rect 998 596 1190 825
rect 1290 665 1394 852
rect 1290 619 1319 665
rect 1365 619 1394 665
rect 1290 596 1394 619
rect 1494 825 1567 852
rect 1613 852 1626 871
rect 1613 825 1686 852
rect 1494 596 1686 825
rect 1786 665 1890 852
rect 1786 619 1815 665
rect 1861 619 1890 665
rect 1786 596 1890 619
rect 1990 839 2078 852
rect 1990 699 2019 839
rect 2065 699 2078 839
rect 1990 596 2078 699
rect 2272 759 2360 852
rect 2272 619 2285 759
rect 2331 619 2360 759
rect 2272 596 2360 619
rect 2460 759 2564 852
rect 2460 619 2489 759
rect 2535 619 2564 759
rect 2460 596 2564 619
rect 2664 759 2752 852
rect 2664 619 2693 759
rect 2739 619 2752 759
rect 2664 596 2752 619
rect 2832 759 2920 852
rect 2832 619 2845 759
rect 2891 619 2920 759
rect 2832 596 2920 619
rect 3020 831 3136 852
rect 3020 691 3049 831
rect 3095 691 3136 831
rect 3020 596 3136 691
rect 3236 759 3360 852
rect 3236 619 3265 759
rect 3311 619 3360 759
rect 3236 596 3360 619
rect 3460 759 3584 852
rect 3460 619 3489 759
rect 3535 619 3584 759
rect 3460 596 3584 619
rect 3684 759 3788 852
rect 3684 619 3713 759
rect 3759 619 3788 759
rect 3684 596 3788 619
rect 3888 759 4012 852
rect 3888 619 3917 759
rect 3963 619 4012 759
rect 3888 596 4012 619
rect 4112 759 4200 852
rect 4112 619 4141 759
rect 4187 619 4200 759
rect 4112 596 4200 619
<< mvndiffc >>
rect 62 257 108 303
rect 286 257 332 303
rect 646 257 692 303
rect 870 257 916 303
rect 1094 257 1140 303
rect 1318 257 1364 303
rect 1542 257 1588 303
rect 1766 257 1812 303
rect 1990 257 2036 303
rect 2174 257 2220 303
rect 2401 257 2447 303
rect 2625 257 2671 303
rect 2817 257 2863 303
rect 3041 257 3087 303
rect 3265 257 3311 303
rect 3489 257 3535 303
rect 3713 257 3759 303
rect 3937 257 3983 303
rect 4161 257 4207 303
<< mvpdiffc >>
rect 82 619 128 759
rect 286 619 332 759
rect 558 619 604 759
rect 823 619 869 665
rect 1071 825 1117 871
rect 1319 619 1365 665
rect 1567 825 1613 871
rect 1815 619 1861 665
rect 2019 699 2065 839
rect 2285 619 2331 759
rect 2489 619 2535 759
rect 2693 619 2739 759
rect 2845 619 2891 759
rect 3049 691 3095 831
rect 3265 619 3311 759
rect 3489 619 3535 759
rect 3713 619 3759 759
rect 3917 619 3963 759
rect 4141 619 4187 759
<< polysilicon >>
rect 655 944 3460 984
rect 157 852 257 896
rect 429 852 529 896
rect 655 852 755 944
rect 898 852 998 896
rect 1190 852 1290 896
rect 1394 852 1494 896
rect 1686 852 1786 896
rect 1890 852 1990 896
rect 2360 852 2460 896
rect 2564 852 2664 896
rect 2920 852 3020 896
rect 3136 852 3236 896
rect 3360 852 3460 944
rect 3584 944 4112 984
rect 3584 852 3684 944
rect 3788 852 3888 896
rect 4012 852 4112 944
rect 157 531 257 596
rect 157 485 170 531
rect 216 485 257 531
rect 157 363 257 485
rect 429 531 529 596
rect 429 485 470 531
rect 516 485 529 531
rect 655 528 755 596
rect 429 472 529 485
rect 577 494 755 528
rect 898 531 998 596
rect 577 471 677 494
rect 898 485 926 531
rect 972 485 998 531
rect 898 472 998 485
rect 577 363 617 471
rect 718 433 841 446
rect 718 387 731 433
rect 777 387 841 433
rect 718 379 841 387
rect 137 319 257 363
rect 497 319 617 363
rect 721 319 841 379
rect 945 363 998 472
rect 1190 511 1290 596
rect 1394 536 1494 596
rect 1686 536 1786 596
rect 1394 511 1786 536
rect 1890 531 1990 596
rect 1890 511 1931 531
rect 1190 485 1931 511
rect 1977 485 1990 531
rect 2360 536 2460 596
rect 2564 555 2664 596
rect 2360 496 2516 536
rect 2564 509 2581 555
rect 2627 536 2664 555
rect 2920 552 3020 596
rect 2920 536 3012 552
rect 2627 509 3012 536
rect 2564 496 3012 509
rect 1190 472 1990 485
rect 1190 471 1961 472
rect 1190 363 1289 471
rect 945 319 1065 363
rect 1169 319 1289 363
rect 1393 319 1513 471
rect 1617 319 1737 471
rect 1841 319 1961 471
rect 2476 448 2516 496
rect 2252 435 2428 448
rect 2252 389 2369 435
rect 2415 389 2428 435
rect 2252 376 2428 389
rect 2476 435 2844 448
rect 2476 389 2785 435
rect 2831 389 2844 435
rect 2476 376 2844 389
rect 2252 316 2372 376
rect 2476 316 2596 376
rect 2892 316 3012 496
rect 3136 531 3236 596
rect 3136 485 3166 531
rect 3212 485 3236 531
rect 3136 360 3236 485
rect 3360 500 3460 596
rect 3584 552 3684 596
rect 3360 487 3740 500
rect 3360 460 3681 487
rect 3564 441 3681 460
rect 3727 441 3740 487
rect 3564 428 3740 441
rect 3116 316 3236 360
rect 3340 316 3460 360
rect 3564 316 3684 428
rect 3788 408 3888 596
rect 3788 395 3908 408
rect 3788 349 3838 395
rect 3884 349 3908 395
rect 3788 316 3908 349
rect 4012 360 4112 596
rect 4012 316 4132 360
rect 137 115 257 159
rect 497 115 617 159
rect 721 64 841 159
rect 945 115 1065 159
rect 1169 115 1289 159
rect 1393 115 1513 159
rect 1617 115 1737 159
rect 1841 115 1961 159
rect 2252 112 2372 156
rect 2476 112 2596 156
rect 2892 112 3012 156
rect 3116 112 3236 156
rect 3340 64 3460 156
rect 3564 112 3684 156
rect 3788 112 3908 156
rect 4012 64 4132 156
rect 721 24 4132 64
<< polycontact >>
rect 170 485 216 531
rect 470 485 516 531
rect 926 485 972 531
rect 731 387 777 433
rect 1931 485 1977 531
rect 2581 509 2627 555
rect 2369 389 2415 435
rect 2785 389 2831 435
rect 3166 485 3212 531
rect 3681 441 3727 487
rect 3838 349 3884 395
<< metal1 >>
rect 0 918 4256 1098
rect 82 759 128 918
rect 1071 871 1117 918
rect 1071 814 1117 825
rect 1567 871 1613 918
rect 1567 814 1613 825
rect 2019 839 2065 918
rect 82 608 128 619
rect 286 759 332 770
rect 140 531 216 542
rect 140 485 170 531
rect 140 466 216 485
rect 62 303 108 314
rect 62 90 108 257
rect 286 303 332 619
rect 378 768 604 770
rect 378 759 1973 768
rect 378 722 558 759
rect 378 303 424 722
rect 604 722 1973 759
rect 558 608 604 619
rect 823 665 869 676
rect 470 531 516 542
rect 470 444 516 485
rect 470 433 777 444
rect 470 387 731 433
rect 470 354 777 387
rect 823 385 869 619
rect 1318 665 1365 676
rect 1318 619 1319 665
rect 926 531 978 542
rect 972 485 978 531
rect 926 430 978 485
rect 1318 406 1365 619
rect 1815 665 1874 676
rect 1861 619 1874 665
rect 1815 406 1874 619
rect 1927 642 1973 722
rect 2693 816 3003 862
rect 2019 688 2065 699
rect 2285 759 2331 770
rect 2189 642 2285 654
rect 1927 619 2285 642
rect 1927 608 2331 619
rect 2489 759 2535 770
rect 1927 596 2220 608
rect 823 339 916 385
rect 870 303 916 339
rect 1318 360 1874 406
rect 1931 531 1977 542
rect 1931 406 1977 485
rect 1931 360 2128 406
rect 378 257 646 303
rect 692 257 703 303
rect 286 246 332 257
rect 870 246 916 257
rect 1094 303 1140 314
rect 1094 90 1140 257
rect 1318 303 1364 360
rect 1318 246 1364 257
rect 1542 303 1588 314
rect 1542 90 1588 257
rect 1766 303 1874 360
rect 1812 257 1874 303
rect 1766 242 1874 257
rect 1990 303 2036 314
rect 1990 90 2036 257
rect 2082 200 2128 360
rect 2174 303 2220 596
rect 2489 527 2535 619
rect 2693 759 2739 816
rect 2174 246 2220 257
rect 2266 481 2535 527
rect 2581 555 2627 566
rect 2266 200 2312 481
rect 2581 435 2627 509
rect 2358 389 2369 435
rect 2415 389 2627 435
rect 2401 303 2447 314
rect 2401 200 2447 257
rect 2494 242 2546 389
rect 2693 314 2739 619
rect 2625 303 2739 314
rect 2671 257 2739 303
rect 2625 246 2739 257
rect 2785 759 2891 770
rect 2785 619 2845 759
rect 2785 435 2891 619
rect 2957 634 3003 816
rect 3049 831 3095 918
rect 3049 680 3095 691
rect 3141 816 3535 862
rect 3141 634 3187 816
rect 2957 588 3187 634
rect 3265 759 3311 770
rect 2831 389 2891 435
rect 3166 531 3218 542
rect 3212 485 3218 531
rect 3166 430 3218 485
rect 2785 303 2891 389
rect 2785 257 2817 303
rect 2863 257 2891 303
rect 2785 246 2891 257
rect 3041 303 3087 314
rect 2082 154 2447 200
rect 3041 90 3087 257
rect 3265 303 3311 619
rect 3265 246 3311 257
rect 3489 759 3535 816
rect 3489 303 3535 619
rect 3713 759 3759 770
rect 3713 590 3759 619
rect 3917 759 3963 918
rect 3917 608 3963 619
rect 4141 759 4207 770
rect 4187 619 4207 759
rect 3589 544 3759 590
rect 3589 303 3635 544
rect 4141 498 4207 619
rect 3681 487 4207 498
rect 3727 452 4207 487
rect 3681 430 3727 441
rect 3838 395 3890 406
rect 3884 349 3890 395
rect 3589 257 3713 303
rect 3759 257 3770 303
rect 3489 246 3535 257
rect 3838 242 3890 349
rect 3937 303 3983 314
rect 3937 90 3983 257
rect 4161 303 4207 452
rect 4161 246 4207 257
rect 0 -90 4256 90
<< labels >>
flabel metal1 s 3838 242 3890 406 0 FreeSans 200 0 0 0 I0
port 1 nsew default input
flabel metal1 s 3166 430 3218 542 0 FreeSans 200 0 0 0 I1
port 2 nsew default input
flabel metal1 s 140 466 216 542 0 FreeSans 200 0 0 0 I2
port 3 nsew default input
flabel metal1 s 926 430 978 542 0 FreeSans 200 0 0 0 I3
port 4 nsew default input
flabel metal1 s 470 444 516 542 0 FreeSans 200 0 0 0 S0
port 5 nsew default input
flabel metal1 s 2581 435 2627 566 0 FreeSans 200 0 0 0 S1
port 6 nsew default input
flabel metal1 s 0 918 4256 1098 0 FreeSans 200 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 3937 90 3983 314 0 FreeSans 200 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 1815 406 1874 676 0 FreeSans 200 0 0 0 Z
port 7 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 9 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 10 nsew ground bidirectional
rlabel metal1 s 470 354 777 444 1 S0
port 5 nsew default input
rlabel metal1 s 2358 389 2627 435 1 S1
port 6 nsew default input
rlabel metal1 s 2494 242 2546 389 1 S1
port 6 nsew default input
rlabel metal1 s 1318 406 1365 676 1 Z
port 7 nsew default output
rlabel metal1 s 1318 360 1874 406 1 Z
port 7 nsew default output
rlabel metal1 s 1766 246 1874 360 1 Z
port 7 nsew default output
rlabel metal1 s 1318 246 1364 360 1 Z
port 7 nsew default output
rlabel metal1 s 1766 242 1874 246 1 Z
port 7 nsew default output
rlabel metal1 s 3917 814 3963 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3049 814 3095 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2019 814 2065 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1567 814 1613 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1071 814 1117 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 82 814 128 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3917 688 3963 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3049 688 3095 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2019 688 2065 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 82 688 128 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3917 680 3963 688 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3049 680 3095 688 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 82 680 128 688 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3917 608 3963 680 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 82 608 128 680 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3041 90 3087 314 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 1990 90 2036 314 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 1542 90 1588 314 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 1094 90 1140 314 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 62 90 108 314 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4256 90 1 VSS
port 11 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4256 1008
string GDS_END 33272
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 23692
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
