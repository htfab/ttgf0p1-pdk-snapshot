magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< nwell >>
rect -86 377 1990 870
rect -86 352 680 377
rect 904 352 1990 377
<< pwell >>
rect 680 352 904 377
rect -86 -86 1990 352
<< mvnmos >>
rect 126 68 246 232
rect 350 68 470 232
rect 574 68 694 232
rect 986 68 1106 232
rect 1210 68 1330 232
rect 1434 68 1554 232
rect 1658 68 1778 232
<< mvpmos >>
rect 175 497 275 716
rect 379 497 479 716
rect 583 497 683 716
rect 1056 480 1156 716
rect 1260 480 1360 716
rect 1464 480 1564 716
rect 1678 480 1778 716
<< mvndiff >>
rect 754 244 826 257
rect 754 232 767 244
rect 38 192 126 232
rect 38 146 51 192
rect 97 146 126 192
rect 38 68 126 146
rect 246 139 350 232
rect 246 93 275 139
rect 321 93 350 139
rect 246 68 350 93
rect 470 166 574 232
rect 470 120 499 166
rect 545 120 574 166
rect 470 68 574 120
rect 694 198 767 232
rect 813 198 826 244
rect 694 68 826 198
rect 898 152 986 232
rect 898 106 911 152
rect 957 106 986 152
rect 898 68 986 106
rect 1106 127 1210 232
rect 1106 81 1135 127
rect 1181 81 1210 127
rect 1106 68 1210 81
rect 1330 192 1434 232
rect 1330 146 1359 192
rect 1405 146 1434 192
rect 1330 68 1434 146
rect 1554 173 1658 232
rect 1554 127 1583 173
rect 1629 127 1658 173
rect 1554 68 1658 127
rect 1778 173 1866 232
rect 1778 127 1807 173
rect 1853 127 1866 173
rect 1778 68 1866 127
<< mvpdiff >>
rect 87 665 175 716
rect 87 525 100 665
rect 146 525 175 665
rect 87 497 175 525
rect 275 703 379 716
rect 275 563 304 703
rect 350 563 379 703
rect 275 497 379 563
rect 479 671 583 716
rect 479 625 508 671
rect 554 625 583 671
rect 479 497 583 625
rect 683 567 771 716
rect 683 521 712 567
rect 758 521 771 567
rect 683 497 771 521
rect 968 652 1056 716
rect 968 512 981 652
rect 1027 512 1056 652
rect 968 480 1056 512
rect 1156 635 1260 716
rect 1156 589 1185 635
rect 1231 589 1260 635
rect 1156 480 1260 589
rect 1360 544 1464 716
rect 1360 498 1389 544
rect 1435 498 1464 544
rect 1360 480 1464 498
rect 1564 653 1678 716
rect 1564 607 1593 653
rect 1639 607 1678 653
rect 1564 480 1678 607
rect 1778 665 1866 716
rect 1778 525 1807 665
rect 1853 525 1866 665
rect 1778 480 1866 525
<< mvndiffc >>
rect 51 146 97 192
rect 275 93 321 139
rect 499 120 545 166
rect 767 198 813 244
rect 911 106 957 152
rect 1135 81 1181 127
rect 1359 146 1405 192
rect 1583 127 1629 173
rect 1807 127 1853 173
<< mvpdiffc >>
rect 100 525 146 665
rect 304 563 350 703
rect 508 625 554 671
rect 712 521 758 567
rect 981 512 1027 652
rect 1185 589 1231 635
rect 1389 498 1435 544
rect 1593 607 1639 653
rect 1807 525 1853 665
<< polysilicon >>
rect 175 716 275 760
rect 379 716 479 760
rect 583 716 683 760
rect 1056 716 1156 760
rect 1260 716 1360 760
rect 1464 716 1564 760
rect 1678 716 1778 760
rect 175 412 275 497
rect 379 412 479 497
rect 583 464 683 497
rect 583 418 596 464
rect 642 418 683 464
rect 126 385 535 412
rect 583 405 683 418
rect 1056 447 1156 480
rect 126 339 165 385
rect 211 372 535 385
rect 211 339 246 372
rect 126 232 246 339
rect 495 357 535 372
rect 1056 401 1083 447
rect 1129 401 1156 447
rect 1056 388 1156 401
rect 1260 439 1360 480
rect 1260 393 1273 439
rect 1319 420 1360 439
rect 1464 420 1564 480
rect 1319 393 1564 420
rect 350 311 427 324
rect 495 317 614 357
rect 350 265 368 311
rect 414 276 427 311
rect 574 288 614 317
rect 414 265 470 276
rect 350 232 470 265
rect 574 232 694 288
rect 1056 287 1106 388
rect 1260 380 1564 393
rect 1678 400 1778 480
rect 1678 354 1698 400
rect 1744 354 1778 400
rect 986 232 1106 287
rect 1210 314 1554 332
rect 1210 268 1267 314
rect 1313 292 1554 314
rect 1313 268 1330 292
rect 1210 232 1330 268
rect 1434 232 1554 292
rect 1678 287 1778 354
rect 1658 232 1778 287
rect 126 24 246 68
rect 350 24 470 68
rect 574 24 694 68
rect 986 24 1106 68
rect 1210 24 1330 68
rect 1434 24 1554 68
rect 1658 24 1778 68
<< polycontact >>
rect 596 418 642 464
rect 165 339 211 385
rect 1083 401 1129 447
rect 1273 393 1319 439
rect 368 265 414 311
rect 1698 354 1744 400
rect 1267 268 1313 314
<< metal1 >>
rect 0 724 1904 844
rect 293 703 361 724
rect 100 665 146 676
rect 293 563 304 703
rect 350 563 361 703
rect 489 625 508 671
rect 554 652 1027 671
rect 554 625 981 652
rect 711 567 758 578
rect 100 517 146 525
rect 711 521 712 567
rect 100 471 642 517
rect 368 464 642 471
rect 82 385 318 425
rect 82 339 165 385
rect 211 339 318 385
rect 82 325 318 339
rect 368 418 596 464
rect 368 407 642 418
rect 368 311 414 407
rect 711 361 758 521
rect 368 245 414 265
rect 51 198 414 245
rect 597 315 758 361
rect 51 192 97 198
rect 597 177 643 315
rect 804 311 850 625
rect 1185 635 1231 724
rect 1185 578 1231 589
rect 1277 614 1547 660
rect 1277 532 1323 614
rect 981 493 1027 512
rect 1083 485 1323 532
rect 1376 544 1435 560
rect 1376 498 1389 544
rect 1501 550 1547 614
rect 1593 653 1639 724
rect 1593 596 1639 607
rect 1804 665 1857 676
rect 1804 550 1807 665
rect 1501 525 1807 550
rect 1853 525 1857 665
rect 1501 504 1857 525
rect 1083 447 1129 485
rect 1083 383 1129 401
rect 1175 393 1273 439
rect 1319 393 1330 439
rect 1175 311 1221 393
rect 1376 332 1435 498
rect 804 269 1221 311
rect 754 265 1221 269
rect 1267 314 1313 328
rect 754 244 850 265
rect 754 198 767 244
rect 813 198 850 244
rect 1267 219 1313 268
rect 499 166 643 177
rect 51 114 97 146
rect 275 139 321 152
rect 545 152 643 166
rect 1032 173 1313 219
rect 1359 192 1435 332
rect 1481 400 1755 438
rect 1481 354 1698 400
rect 1744 354 1755 400
rect 1481 328 1755 354
rect 1481 232 1554 328
rect 1032 152 1078 173
rect 545 120 911 152
rect 499 106 911 120
rect 957 106 1078 152
rect 1405 146 1435 192
rect 275 60 321 93
rect 1124 81 1135 127
rect 1181 81 1192 127
rect 1359 106 1435 146
rect 1583 173 1629 184
rect 1124 60 1192 81
rect 1583 60 1629 127
rect 1804 173 1857 504
rect 1804 127 1807 173
rect 1853 127 1857 173
rect 1804 116 1857 127
rect 0 -60 1904 60
<< labels >>
flabel metal1 s 0 724 1904 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 1583 152 1629 184 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 1376 332 1435 560 0 FreeSans 400 0 0 0 ZN
port 3 nsew default output
flabel metal1 s 82 325 318 425 0 FreeSans 400 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1481 328 1755 438 0 FreeSans 400 0 0 0 I
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 5 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 1481 232 1554 328 1 I
port 2 nsew default input
rlabel metal1 s 1359 106 1435 332 1 ZN
port 3 nsew default output
rlabel metal1 s 1593 596 1639 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1185 596 1231 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 293 596 361 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1185 578 1231 596 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 293 578 361 596 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 293 563 361 578 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1583 127 1629 152 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 275 127 321 152 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1583 60 1629 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1124 60 1192 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 275 60 321 127 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1904 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1904 784
string GDS_END 527620
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 522194
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
