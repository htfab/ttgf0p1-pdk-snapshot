VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tie_diff_w2
  CLASS BLOCK ;
  FOREIGN tie_diff_w2 ;
  ORIGIN 0.430 0.000 ;
  SIZE 3.140 BY 7.430 ;
  PIN vdd
    ANTENNADIFFAREA 4.682400 ;
    PORT
      LAYER Nwell ;
        RECT -0.430 3.400 2.710 7.430 ;
      LAYER Metal1 ;
        RECT 0.000 5.660 2.280 7.000 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 4.370400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 0.000 2.280 1.340 ;
    END
  END vss
END tie_diff_w2
END LIBRARY

