magic
tech gf180mcuD
magscale 1 10
timestamp 1753445457
<< nwell >>
rect -86 354 1542 870
<< pwell >>
rect -86 -86 1542 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 724 68 780 268
rect 901 68 957 268
rect 1061 68 1117 268
rect 1221 68 1277 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 724 440 780 716
rect 901 440 957 716
rect 1061 440 1117 716
rect 1221 440 1277 716
<< ndiff >>
rect 28 127 116 268
rect 28 81 41 127
rect 87 81 116 127
rect 28 68 116 81
rect 172 68 276 268
rect 332 248 436 268
rect 332 202 361 248
rect 407 202 436 248
rect 332 68 436 202
rect 492 127 724 268
rect 492 81 521 127
rect 695 81 724 127
rect 492 68 724 81
rect 780 255 901 268
rect 780 209 826 255
rect 872 209 901 255
rect 780 68 901 209
rect 957 255 1061 268
rect 957 81 986 255
rect 1032 81 1061 255
rect 957 68 1061 81
rect 1117 255 1221 268
rect 1117 209 1146 255
rect 1192 209 1221 255
rect 1117 68 1221 209
rect 1277 255 1368 268
rect 1277 81 1306 255
rect 1352 81 1368 255
rect 1277 68 1368 81
<< pdiff >>
rect 28 595 116 716
rect 28 549 41 595
rect 87 549 116 595
rect 28 440 116 549
rect 172 703 276 716
rect 172 657 201 703
rect 247 657 276 703
rect 172 440 276 657
rect 332 595 436 716
rect 332 549 361 595
rect 407 549 436 595
rect 332 440 436 549
rect 492 667 580 716
rect 492 456 521 667
rect 567 456 580 667
rect 492 440 580 456
rect 636 703 724 716
rect 636 453 649 703
rect 695 453 724 703
rect 636 440 724 453
rect 780 665 901 716
rect 780 453 826 665
rect 872 453 901 665
rect 780 440 901 453
rect 957 703 1061 716
rect 957 453 986 703
rect 1032 453 1061 703
rect 957 440 1061 453
rect 1117 665 1221 716
rect 1117 453 1146 665
rect 1192 453 1221 665
rect 1117 440 1221 453
rect 1277 703 1368 716
rect 1277 453 1306 703
rect 1352 453 1368 703
rect 1277 440 1368 453
<< ndiffc >>
rect 41 81 87 127
rect 361 202 407 248
rect 521 81 695 127
rect 826 209 872 255
rect 986 81 1032 255
rect 1146 209 1192 255
rect 1306 81 1352 255
<< pdiffc >>
rect 41 549 87 595
rect 201 657 247 703
rect 361 549 407 595
rect 521 456 567 667
rect 649 453 695 703
rect 826 453 872 665
rect 986 453 1032 703
rect 1146 453 1192 665
rect 1306 453 1352 703
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 724 716 780 760
rect 901 716 957 760
rect 1061 716 1117 760
rect 1221 716 1277 760
rect 116 393 172 440
rect 276 393 332 440
rect 436 393 492 440
rect 80 376 172 393
rect 80 330 102 376
rect 148 330 172 376
rect 80 316 172 330
rect 240 377 332 393
rect 240 331 265 377
rect 311 331 332 377
rect 240 316 332 331
rect 400 379 492 393
rect 724 391 780 440
rect 400 333 423 379
rect 469 333 492 379
rect 400 316 492 333
rect 692 377 780 391
rect 901 377 957 440
rect 692 331 714 377
rect 760 348 957 377
rect 1061 377 1117 440
rect 1221 377 1277 440
rect 1061 348 1277 377
rect 760 331 1277 348
rect 692 317 780 331
rect 116 268 172 316
rect 276 268 332 316
rect 436 268 492 316
rect 724 268 780 317
rect 901 301 1117 331
rect 901 268 957 301
rect 1061 268 1117 301
rect 1221 268 1277 331
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 724 24 780 68
rect 901 24 957 68
rect 1061 24 1117 68
rect 1221 24 1277 68
<< polycontact >>
rect 102 330 148 376
rect 265 331 311 377
rect 423 333 469 379
rect 714 331 760 377
<< metal1 >>
rect 0 724 1456 844
rect 201 703 247 724
rect 649 703 695 724
rect 201 646 247 657
rect 521 667 567 678
rect 41 595 87 620
rect 361 595 407 609
rect 87 549 361 595
rect 41 533 87 549
rect 361 534 407 549
rect 80 376 172 472
rect 567 456 585 495
rect 521 445 585 456
rect 80 330 102 376
rect 148 330 172 376
rect 80 316 172 330
rect 240 377 332 393
rect 240 331 265 377
rect 311 331 332 377
rect 240 316 332 331
rect 400 379 492 393
rect 400 333 423 379
rect 469 333 492 379
rect 400 316 492 333
rect 539 377 585 445
rect 986 703 1032 724
rect 649 429 695 453
rect 826 665 890 676
rect 872 453 890 665
rect 826 378 890 453
rect 1306 703 1352 724
rect 986 429 1032 453
rect 1146 665 1210 676
rect 1192 453 1210 665
rect 1146 378 1210 453
rect 1306 429 1352 453
rect 539 331 714 377
rect 760 331 780 377
rect 826 332 1210 378
rect 539 248 585 331
rect 349 202 361 248
rect 407 202 585 248
rect 826 255 890 332
rect 872 209 890 255
rect 826 198 890 209
rect 986 255 1032 276
rect 41 127 87 138
rect 41 60 87 81
rect 521 127 695 138
rect 521 60 695 81
rect 1146 255 1210 332
rect 1192 209 1210 255
rect 1146 198 1210 209
rect 1306 255 1352 276
rect 986 60 1032 81
rect 1306 60 1352 81
rect 0 -60 1456 60
<< labels >>
flabel metal1 s 0 724 1456 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1456 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 826 198 890 676 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 80 316 172 472 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 240 316 332 393 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel metal1 400 316 492 393 0 FreeSans 200 0 0 0 C
port 8 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1456 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
