magic
tech gf180mcuD
magscale 1 10
timestamp 1753579406
<< nwell >>
rect -86 354 1654 870
<< pwell >>
rect -86 -86 1654 354
<< nmos >>
rect 116 68 172 268
rect 276 68 332 268
rect 436 68 492 268
rect 596 68 652 268
rect 891 68 947 268
rect 1051 68 1107 268
rect 1211 68 1267 268
rect 1371 68 1427 268
<< pmos >>
rect 116 440 172 716
rect 276 440 332 716
rect 436 440 492 716
rect 596 440 652 716
rect 891 440 947 716
rect 1051 440 1107 716
rect 1211 440 1267 716
rect 1371 440 1427 716
<< ndiff >>
rect 28 189 116 268
rect 28 143 41 189
rect 87 143 116 189
rect 28 68 116 143
rect 172 127 276 268
rect 172 81 201 127
rect 247 81 276 127
rect 172 68 276 81
rect 332 198 436 268
rect 332 152 361 198
rect 407 152 436 198
rect 332 68 436 152
rect 492 248 596 268
rect 492 202 521 248
rect 567 202 596 248
rect 492 68 596 202
rect 652 152 740 268
rect 652 106 681 152
rect 727 106 740 152
rect 652 68 740 106
rect 803 156 891 268
rect 803 110 816 156
rect 862 110 891 156
rect 803 68 891 110
rect 947 248 1051 268
rect 947 202 976 248
rect 1022 202 1051 248
rect 947 68 1051 202
rect 1107 200 1211 268
rect 1107 154 1136 200
rect 1182 154 1211 200
rect 1107 68 1211 154
rect 1267 127 1371 268
rect 1267 81 1296 127
rect 1342 81 1371 127
rect 1267 68 1371 81
rect 1427 248 1540 268
rect 1427 202 1456 248
rect 1502 202 1540 248
rect 1427 68 1540 202
<< pdiff >>
rect 28 552 116 716
rect 28 506 41 552
rect 87 506 116 552
rect 28 440 116 506
rect 172 678 276 716
rect 172 632 201 678
rect 247 632 276 678
rect 172 440 276 632
rect 332 556 436 716
rect 332 510 361 556
rect 407 510 436 556
rect 332 440 436 510
rect 492 678 596 716
rect 492 632 521 678
rect 567 632 596 678
rect 492 440 596 632
rect 652 556 740 716
rect 652 510 681 556
rect 727 510 740 556
rect 652 440 740 510
rect 803 579 891 716
rect 803 533 816 579
rect 862 533 891 579
rect 803 440 891 533
rect 947 703 1051 716
rect 947 657 976 703
rect 1022 657 1051 703
rect 947 440 1051 657
rect 1107 553 1211 716
rect 1107 507 1136 553
rect 1182 507 1211 553
rect 1107 440 1211 507
rect 1267 703 1371 716
rect 1267 657 1296 703
rect 1342 657 1371 703
rect 1267 440 1371 657
rect 1427 564 1540 716
rect 1427 518 1456 564
rect 1502 518 1540 564
rect 1427 440 1540 518
<< ndiffc >>
rect 41 143 87 189
rect 201 81 247 127
rect 361 152 407 198
rect 521 202 567 248
rect 681 106 727 152
rect 816 110 862 156
rect 976 202 1022 248
rect 1136 154 1182 200
rect 1296 81 1342 127
rect 1456 202 1502 248
<< pdiffc >>
rect 41 506 87 552
rect 201 632 247 678
rect 361 510 407 556
rect 521 632 567 678
rect 681 510 727 556
rect 816 533 862 579
rect 976 657 1022 703
rect 1136 507 1182 553
rect 1296 657 1342 703
rect 1456 518 1502 564
<< polysilicon >>
rect 116 716 172 760
rect 276 716 332 760
rect 436 716 492 760
rect 596 716 652 760
rect 891 716 947 760
rect 1051 716 1107 760
rect 1211 716 1267 760
rect 1371 716 1427 760
rect 116 393 172 440
rect 276 393 332 440
rect 116 380 332 393
rect 116 334 129 380
rect 319 334 332 380
rect 116 318 332 334
rect 116 268 172 318
rect 276 268 332 318
rect 436 393 492 440
rect 596 393 652 440
rect 436 380 652 393
rect 436 334 449 380
rect 639 334 652 380
rect 436 318 652 334
rect 436 268 492 318
rect 596 268 652 318
rect 891 393 947 440
rect 1051 393 1107 440
rect 891 377 1107 393
rect 891 331 904 377
rect 1094 331 1107 377
rect 891 318 1107 331
rect 891 268 947 318
rect 1051 268 1107 318
rect 1211 393 1267 440
rect 1371 393 1427 440
rect 1211 377 1427 393
rect 1211 331 1224 377
rect 1414 331 1427 377
rect 1211 318 1427 331
rect 1211 268 1267 318
rect 1371 268 1427 318
rect 116 24 172 68
rect 276 24 332 68
rect 436 24 492 68
rect 596 24 652 68
rect 891 24 947 68
rect 1051 24 1107 68
rect 1211 24 1267 68
rect 1371 24 1427 68
<< polycontact >>
rect 129 334 319 380
rect 449 334 639 380
rect 904 331 1094 377
rect 1224 331 1414 377
<< metal1 >>
rect 0 724 1568 844
rect 976 703 1022 724
rect 187 632 201 678
rect 247 632 521 678
rect 567 632 862 678
rect 976 646 1022 657
rect 1296 703 1342 724
rect 1296 646 1342 657
rect 816 579 862 632
rect 41 552 87 563
rect 361 556 744 576
rect 87 510 361 530
rect 407 530 681 556
rect 87 506 407 510
rect 41 484 407 506
rect 727 510 744 556
rect 681 496 744 510
rect 1456 564 1502 577
rect 862 533 1136 553
rect 816 507 1136 533
rect 1182 518 1456 553
rect 1182 507 1502 518
rect 698 467 744 496
rect 116 380 328 393
rect 116 334 129 380
rect 319 334 328 380
rect 116 318 328 334
rect 436 380 652 393
rect 436 334 449 380
rect 639 334 652 380
rect 436 318 652 334
rect 698 248 786 467
rect 891 377 1107 393
rect 891 331 904 377
rect 1094 331 1107 377
rect 891 318 1107 331
rect 1211 377 1427 393
rect 1211 331 1224 377
rect 1414 331 1427 377
rect 1211 318 1427 331
rect 41 200 407 246
rect 494 202 521 248
rect 567 202 976 248
rect 1022 202 1038 248
rect 1136 202 1456 248
rect 1502 202 1513 248
rect 41 189 87 200
rect 41 107 87 143
rect 361 198 407 200
rect 1136 200 1182 202
rect 201 127 247 138
rect 361 106 681 152
rect 727 106 738 152
rect 803 110 816 156
rect 862 154 1136 156
rect 862 110 1182 154
rect 1296 127 1342 138
rect 201 60 247 81
rect 1296 60 1342 81
rect 0 -60 1568 60
<< labels >>
flabel metal1 s 0 724 1568 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 1568 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 698 202 786 467 0 FreeSans 200 0 0 0 Y
port 5 nsew signal output
flabel metal1 116 318 328 393 0 FreeSans 200 0 0 0 A
port 6 nsew signal input
flabel metal1 436 318 652 393 0 FreeSans 200 0 0 0 B
port 7 nsew signal input
flabel metal1 891 318 1107 393 0 FreeSans 200 0 0 0 C
port 8 nsew signal input
flabel metal1 1211 318 1427 393 0 FreeSans 200 0 0 0 D
port 9 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1568 784
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y
<< end >>
