magic
tech gf180mcuD
magscale 1 10
timestamp 1755005639
<< metal1 >>
rect 14757 50970 14833 50982
rect 14757 50918 14769 50970
rect 14821 50918 14833 50970
rect 14757 50862 14833 50918
rect 14757 50810 14769 50862
rect 14821 50810 14833 50862
rect 14757 50754 14833 50810
rect 14757 50702 14769 50754
rect 14821 50702 14833 50754
rect 14757 50646 14833 50702
rect 14757 50594 14769 50646
rect 14821 50594 14833 50646
rect 14757 50538 14833 50594
rect 14757 50486 14769 50538
rect 14821 50486 14833 50538
rect 14757 50430 14833 50486
rect 14757 50378 14769 50430
rect 14821 50378 14833 50430
rect 14757 50322 14833 50378
rect 14757 50270 14769 50322
rect 14821 50270 14833 50322
rect 14757 50214 14833 50270
rect 14757 50162 14769 50214
rect 14821 50162 14833 50214
rect 14757 50106 14833 50162
rect 14757 50054 14769 50106
rect 14821 50054 14833 50106
rect 14757 49998 14833 50054
rect 14757 49946 14769 49998
rect 14821 49946 14833 49998
rect 14757 49890 14833 49946
rect 14757 49838 14769 49890
rect 14821 49838 14833 49890
rect 14757 49782 14833 49838
rect 14757 49730 14769 49782
rect 14821 49730 14833 49782
rect 14757 49674 14833 49730
rect 14757 49622 14769 49674
rect 14821 49622 14833 49674
rect 14757 49610 14833 49622
rect 14757 36570 14833 36582
rect 14757 36518 14769 36570
rect 14821 36518 14833 36570
rect 14757 36462 14833 36518
rect 14757 36410 14769 36462
rect 14821 36410 14833 36462
rect 14757 36354 14833 36410
rect 14757 36302 14769 36354
rect 14821 36302 14833 36354
rect 14757 36246 14833 36302
rect 14757 36194 14769 36246
rect 14821 36194 14833 36246
rect 14757 36138 14833 36194
rect 14757 36086 14769 36138
rect 14821 36086 14833 36138
rect 14757 36030 14833 36086
rect 14757 35978 14769 36030
rect 14821 35978 14833 36030
rect 14757 35922 14833 35978
rect 14757 35870 14769 35922
rect 14821 35870 14833 35922
rect 14757 35814 14833 35870
rect 14757 35762 14769 35814
rect 14821 35762 14833 35814
rect 14757 35706 14833 35762
rect 14757 35654 14769 35706
rect 14821 35654 14833 35706
rect 14757 35598 14833 35654
rect 14757 35546 14769 35598
rect 14821 35546 14833 35598
rect 14757 35490 14833 35546
rect 14757 35438 14769 35490
rect 14821 35438 14833 35490
rect 14757 35382 14833 35438
rect 14757 35330 14769 35382
rect 14821 35330 14833 35382
rect 14757 35274 14833 35330
rect 14757 35222 14769 35274
rect 14821 35222 14833 35274
rect 14757 35210 14833 35222
<< via1 >>
rect 14769 50918 14821 50970
rect 14769 50810 14821 50862
rect 14769 50702 14821 50754
rect 14769 50594 14821 50646
rect 14769 50486 14821 50538
rect 14769 50378 14821 50430
rect 14769 50270 14821 50322
rect 14769 50162 14821 50214
rect 14769 50054 14821 50106
rect 14769 49946 14821 49998
rect 14769 49838 14821 49890
rect 14769 49730 14821 49782
rect 14769 49622 14821 49674
rect 14769 36518 14821 36570
rect 14769 36410 14821 36462
rect 14769 36302 14821 36354
rect 14769 36194 14821 36246
rect 14769 36086 14821 36138
rect 14769 35978 14821 36030
rect 14769 35870 14821 35922
rect 14769 35762 14821 35814
rect 14769 35654 14821 35706
rect 14769 35546 14821 35598
rect 14769 35438 14821 35490
rect 14769 35330 14821 35382
rect 14769 35222 14821 35274
<< metal2 >>
rect 7640 56433 8460 56443
rect 6182 56422 7002 56432
rect 6182 56366 6192 56422
rect 6248 56366 6316 56422
rect 6372 56366 6440 56422
rect 6496 56366 6564 56422
rect 6620 56366 6688 56422
rect 6744 56366 6812 56422
rect 6868 56366 6936 56422
rect 6992 56366 7002 56422
rect 6182 56298 7002 56366
rect 6182 56242 6192 56298
rect 6248 56242 6316 56298
rect 6372 56242 6440 56298
rect 6496 56242 6564 56298
rect 6620 56242 6688 56298
rect 6744 56242 6812 56298
rect 6868 56242 6936 56298
rect 6992 56242 7002 56298
rect 6182 56174 7002 56242
rect 6182 56118 6192 56174
rect 6248 56118 6316 56174
rect 6372 56118 6440 56174
rect 6496 56118 6564 56174
rect 6620 56118 6688 56174
rect 6744 56118 6812 56174
rect 6868 56118 6936 56174
rect 6992 56118 7002 56174
rect 6182 56050 7002 56118
rect 6182 55994 6192 56050
rect 6248 55994 6316 56050
rect 6372 55994 6440 56050
rect 6496 55994 6564 56050
rect 6620 55994 6688 56050
rect 6744 55994 6812 56050
rect 6868 55994 6936 56050
rect 6992 55994 7002 56050
rect 6182 55926 7002 55994
rect 6182 55870 6192 55926
rect 6248 55870 6316 55926
rect 6372 55870 6440 55926
rect 6496 55870 6564 55926
rect 6620 55870 6688 55926
rect 6744 55870 6812 55926
rect 6868 55870 6936 55926
rect 6992 55870 7002 55926
rect 6182 55802 7002 55870
rect 6182 55746 6192 55802
rect 6248 55746 6316 55802
rect 6372 55746 6440 55802
rect 6496 55746 6564 55802
rect 6620 55746 6688 55802
rect 6744 55746 6812 55802
rect 6868 55746 6936 55802
rect 6992 55746 7002 55802
rect 6182 55678 7002 55746
rect 6182 55622 6192 55678
rect 6248 55622 6316 55678
rect 6372 55622 6440 55678
rect 6496 55622 6564 55678
rect 6620 55622 6688 55678
rect 6744 55622 6812 55678
rect 6868 55622 6936 55678
rect 6992 55622 7002 55678
rect 6182 55554 7002 55622
rect 6182 55498 6192 55554
rect 6248 55498 6316 55554
rect 6372 55498 6440 55554
rect 6496 55498 6564 55554
rect 6620 55498 6688 55554
rect 6744 55498 6812 55554
rect 6868 55498 6936 55554
rect 6992 55498 7002 55554
rect 6182 55430 7002 55498
rect 6182 55374 6192 55430
rect 6248 55374 6316 55430
rect 6372 55374 6440 55430
rect 6496 55374 6564 55430
rect 6620 55374 6688 55430
rect 6744 55374 6812 55430
rect 6868 55374 6936 55430
rect 6992 55374 7002 55430
rect 6182 55306 7002 55374
rect 6182 55250 6192 55306
rect 6248 55250 6316 55306
rect 6372 55250 6440 55306
rect 6496 55250 6564 55306
rect 6620 55250 6688 55306
rect 6744 55250 6812 55306
rect 6868 55250 6936 55306
rect 6992 55250 7002 55306
rect 6182 55182 7002 55250
rect 6182 55126 6192 55182
rect 6248 55126 6316 55182
rect 6372 55126 6440 55182
rect 6496 55126 6564 55182
rect 6620 55126 6688 55182
rect 6744 55126 6812 55182
rect 6868 55126 6936 55182
rect 6992 55126 7002 55182
rect 6182 55058 7002 55126
rect 6182 55002 6192 55058
rect 6248 55002 6316 55058
rect 6372 55002 6440 55058
rect 6496 55002 6564 55058
rect 6620 55002 6688 55058
rect 6744 55002 6812 55058
rect 6868 55002 6936 55058
rect 6992 55002 7002 55058
rect 6182 54934 7002 55002
rect 6182 54878 6192 54934
rect 6248 54878 6316 54934
rect 6372 54878 6440 54934
rect 6496 54878 6564 54934
rect 6620 54878 6688 54934
rect 6744 54878 6812 54934
rect 6868 54878 6936 54934
rect 6992 54878 7002 54934
rect 6182 54810 7002 54878
rect 6182 54754 6192 54810
rect 6248 54754 6316 54810
rect 6372 54754 6440 54810
rect 6496 54754 6564 54810
rect 6620 54754 6688 54810
rect 6744 54754 6812 54810
rect 6868 54754 6936 54810
rect 6992 54754 7002 54810
rect 6182 54686 7002 54754
rect 6182 54630 6192 54686
rect 6248 54630 6316 54686
rect 6372 54630 6440 54686
rect 6496 54630 6564 54686
rect 6620 54630 6688 54686
rect 6744 54630 6812 54686
rect 6868 54630 6936 54686
rect 6992 54630 7002 54686
rect 6182 54562 7002 54630
rect 6182 54506 6192 54562
rect 6248 54506 6316 54562
rect 6372 54506 6440 54562
rect 6496 54506 6564 54562
rect 6620 54506 6688 54562
rect 6744 54506 6812 54562
rect 6868 54506 6936 54562
rect 6992 54506 7002 54562
rect 6182 54438 7002 54506
rect 6182 54382 6192 54438
rect 6248 54382 6316 54438
rect 6372 54382 6440 54438
rect 6496 54382 6564 54438
rect 6620 54382 6688 54438
rect 6744 54382 6812 54438
rect 6868 54382 6936 54438
rect 6992 54382 7002 54438
rect 6182 54314 7002 54382
rect 6182 54258 6192 54314
rect 6248 54258 6316 54314
rect 6372 54258 6440 54314
rect 6496 54258 6564 54314
rect 6620 54258 6688 54314
rect 6744 54258 6812 54314
rect 6868 54258 6936 54314
rect 6992 54258 7002 54314
rect 6182 54190 7002 54258
rect 6182 54134 6192 54190
rect 6248 54134 6316 54190
rect 6372 54134 6440 54190
rect 6496 54134 6564 54190
rect 6620 54134 6688 54190
rect 6744 54134 6812 54190
rect 6868 54134 6936 54190
rect 6992 54134 7002 54190
rect 6182 54066 7002 54134
rect 6182 54010 6192 54066
rect 6248 54010 6316 54066
rect 6372 54010 6440 54066
rect 6496 54010 6564 54066
rect 6620 54010 6688 54066
rect 6744 54010 6812 54066
rect 6868 54010 6936 54066
rect 6992 54010 7002 54066
rect 6182 53942 7002 54010
rect 6182 53886 6192 53942
rect 6248 53886 6316 53942
rect 6372 53886 6440 53942
rect 6496 53886 6564 53942
rect 6620 53886 6688 53942
rect 6744 53886 6812 53942
rect 6868 53886 6936 53942
rect 6992 53886 7002 53942
rect 6182 53818 7002 53886
rect 6182 53762 6192 53818
rect 6248 53762 6316 53818
rect 6372 53762 6440 53818
rect 6496 53762 6564 53818
rect 6620 53762 6688 53818
rect 6744 53762 6812 53818
rect 6868 53762 6936 53818
rect 6992 53762 7002 53818
rect 6182 53694 7002 53762
rect 6182 53638 6192 53694
rect 6248 53638 6316 53694
rect 6372 53638 6440 53694
rect 6496 53638 6564 53694
rect 6620 53638 6688 53694
rect 6744 53638 6812 53694
rect 6868 53638 6936 53694
rect 6992 53638 7002 53694
rect 6182 53570 7002 53638
rect 6182 53514 6192 53570
rect 6248 53514 6316 53570
rect 6372 53514 6440 53570
rect 6496 53514 6564 53570
rect 6620 53514 6688 53570
rect 6744 53514 6812 53570
rect 6868 53514 6936 53570
rect 6992 53514 7002 53570
rect 6182 53446 7002 53514
rect 6182 53390 6192 53446
rect 6248 53390 6316 53446
rect 6372 53390 6440 53446
rect 6496 53390 6564 53446
rect 6620 53390 6688 53446
rect 6744 53390 6812 53446
rect 6868 53390 6936 53446
rect 6992 53390 7002 53446
rect 6182 53322 7002 53390
rect 6182 53266 6192 53322
rect 6248 53266 6316 53322
rect 6372 53266 6440 53322
rect 6496 53266 6564 53322
rect 6620 53266 6688 53322
rect 6744 53266 6812 53322
rect 6868 53266 6936 53322
rect 6992 53266 7002 53322
rect 6182 53256 7002 53266
rect 7640 56377 7650 56433
rect 7706 56377 7774 56433
rect 7830 56377 7898 56433
rect 7954 56377 8022 56433
rect 8078 56377 8146 56433
rect 8202 56377 8270 56433
rect 8326 56377 8394 56433
rect 8450 56377 8460 56433
rect 7640 56309 8460 56377
rect 7640 56253 7650 56309
rect 7706 56253 7774 56309
rect 7830 56253 7898 56309
rect 7954 56253 8022 56309
rect 8078 56253 8146 56309
rect 8202 56253 8270 56309
rect 8326 56253 8394 56309
rect 8450 56253 8460 56309
rect 7640 56185 8460 56253
rect 7640 56129 7650 56185
rect 7706 56129 7774 56185
rect 7830 56129 7898 56185
rect 7954 56129 8022 56185
rect 8078 56129 8146 56185
rect 8202 56129 8270 56185
rect 8326 56129 8394 56185
rect 8450 56129 8460 56185
rect 7640 56061 8460 56129
rect 7640 56005 7650 56061
rect 7706 56005 7774 56061
rect 7830 56005 7898 56061
rect 7954 56005 8022 56061
rect 8078 56005 8146 56061
rect 8202 56005 8270 56061
rect 8326 56005 8394 56061
rect 8450 56005 8460 56061
rect 7640 55937 8460 56005
rect 7640 55881 7650 55937
rect 7706 55881 7774 55937
rect 7830 55881 7898 55937
rect 7954 55881 8022 55937
rect 8078 55881 8146 55937
rect 8202 55881 8270 55937
rect 8326 55881 8394 55937
rect 8450 55881 8460 55937
rect 7640 55813 8460 55881
rect 7640 55757 7650 55813
rect 7706 55757 7774 55813
rect 7830 55757 7898 55813
rect 7954 55757 8022 55813
rect 8078 55757 8146 55813
rect 8202 55757 8270 55813
rect 8326 55757 8394 55813
rect 8450 55757 8460 55813
rect 7640 55689 8460 55757
rect 7640 55633 7650 55689
rect 7706 55633 7774 55689
rect 7830 55633 7898 55689
rect 7954 55633 8022 55689
rect 8078 55633 8146 55689
rect 8202 55633 8270 55689
rect 8326 55633 8394 55689
rect 8450 55633 8460 55689
rect 7640 55565 8460 55633
rect 7640 55509 7650 55565
rect 7706 55509 7774 55565
rect 7830 55509 7898 55565
rect 7954 55509 8022 55565
rect 8078 55509 8146 55565
rect 8202 55509 8270 55565
rect 8326 55509 8394 55565
rect 8450 55509 8460 55565
rect 7640 55441 8460 55509
rect 7640 55385 7650 55441
rect 7706 55385 7774 55441
rect 7830 55385 7898 55441
rect 7954 55385 8022 55441
rect 8078 55385 8146 55441
rect 8202 55385 8270 55441
rect 8326 55385 8394 55441
rect 8450 55385 8460 55441
rect 7640 55317 8460 55385
rect 7640 55261 7650 55317
rect 7706 55261 7774 55317
rect 7830 55261 7898 55317
rect 7954 55261 8022 55317
rect 8078 55261 8146 55317
rect 8202 55261 8270 55317
rect 8326 55261 8394 55317
rect 8450 55261 8460 55317
rect 7640 55193 8460 55261
rect 7640 55137 7650 55193
rect 7706 55137 7774 55193
rect 7830 55137 7898 55193
rect 7954 55137 8022 55193
rect 8078 55137 8146 55193
rect 8202 55137 8270 55193
rect 8326 55137 8394 55193
rect 8450 55137 8460 55193
rect 7640 55069 8460 55137
rect 7640 55013 7650 55069
rect 7706 55013 7774 55069
rect 7830 55013 7898 55069
rect 7954 55013 8022 55069
rect 8078 55013 8146 55069
rect 8202 55013 8270 55069
rect 8326 55013 8394 55069
rect 8450 55013 8460 55069
rect 7640 54945 8460 55013
rect 7640 54889 7650 54945
rect 7706 54889 7774 54945
rect 7830 54889 7898 54945
rect 7954 54889 8022 54945
rect 8078 54889 8146 54945
rect 8202 54889 8270 54945
rect 8326 54889 8394 54945
rect 8450 54889 8460 54945
rect 7640 54821 8460 54889
rect 7640 54765 7650 54821
rect 7706 54765 7774 54821
rect 7830 54765 7898 54821
rect 7954 54765 8022 54821
rect 8078 54765 8146 54821
rect 8202 54765 8270 54821
rect 8326 54765 8394 54821
rect 8450 54765 8460 54821
rect 7640 54697 8460 54765
rect 7640 54641 7650 54697
rect 7706 54641 7774 54697
rect 7830 54641 7898 54697
rect 7954 54641 8022 54697
rect 8078 54641 8146 54697
rect 8202 54641 8270 54697
rect 8326 54641 8394 54697
rect 8450 54641 8460 54697
rect 7640 54573 8460 54641
rect 7640 54517 7650 54573
rect 7706 54517 7774 54573
rect 7830 54517 7898 54573
rect 7954 54517 8022 54573
rect 8078 54517 8146 54573
rect 8202 54517 8270 54573
rect 8326 54517 8394 54573
rect 8450 54517 8460 54573
rect 7640 54449 8460 54517
rect 7640 54393 7650 54449
rect 7706 54393 7774 54449
rect 7830 54393 7898 54449
rect 7954 54393 8022 54449
rect 8078 54393 8146 54449
rect 8202 54393 8270 54449
rect 8326 54393 8394 54449
rect 8450 54393 8460 54449
rect 7640 54325 8460 54393
rect 7640 54269 7650 54325
rect 7706 54269 7774 54325
rect 7830 54269 7898 54325
rect 7954 54269 8022 54325
rect 8078 54269 8146 54325
rect 8202 54269 8270 54325
rect 8326 54269 8394 54325
rect 8450 54269 8460 54325
rect 7640 54201 8460 54269
rect 7640 54145 7650 54201
rect 7706 54145 7774 54201
rect 7830 54145 7898 54201
rect 7954 54145 8022 54201
rect 8078 54145 8146 54201
rect 8202 54145 8270 54201
rect 8326 54145 8394 54201
rect 8450 54145 8460 54201
rect 7640 54077 8460 54145
rect 7640 54021 7650 54077
rect 7706 54021 7774 54077
rect 7830 54021 7898 54077
rect 7954 54021 8022 54077
rect 8078 54021 8146 54077
rect 8202 54021 8270 54077
rect 8326 54021 8394 54077
rect 8450 54021 8460 54077
rect 7640 53953 8460 54021
rect 7640 53897 7650 53953
rect 7706 53897 7774 53953
rect 7830 53897 7898 53953
rect 7954 53897 8022 53953
rect 8078 53897 8146 53953
rect 8202 53897 8270 53953
rect 8326 53897 8394 53953
rect 8450 53897 8460 53953
rect 7640 53829 8460 53897
rect 7640 53773 7650 53829
rect 7706 53773 7774 53829
rect 7830 53773 7898 53829
rect 7954 53773 8022 53829
rect 8078 53773 8146 53829
rect 8202 53773 8270 53829
rect 8326 53773 8394 53829
rect 8450 53773 8460 53829
rect 7640 53705 8460 53773
rect 7640 53649 7650 53705
rect 7706 53649 7774 53705
rect 7830 53649 7898 53705
rect 7954 53649 8022 53705
rect 8078 53649 8146 53705
rect 8202 53649 8270 53705
rect 8326 53649 8394 53705
rect 8450 53649 8460 53705
rect 7640 53581 8460 53649
rect 7640 53525 7650 53581
rect 7706 53525 7774 53581
rect 7830 53525 7898 53581
rect 7954 53525 8022 53581
rect 8078 53525 8146 53581
rect 8202 53525 8270 53581
rect 8326 53525 8394 53581
rect 8450 53525 8460 53581
rect 7640 53457 8460 53525
rect 7640 53401 7650 53457
rect 7706 53401 7774 53457
rect 7830 53401 7898 53457
rect 7954 53401 8022 53457
rect 8078 53401 8146 53457
rect 8202 53401 8270 53457
rect 8326 53401 8394 53457
rect 8450 53401 8460 53457
rect 7640 53333 8460 53401
rect 7640 53277 7650 53333
rect 7706 53277 7774 53333
rect 7830 53277 7898 53333
rect 7954 53277 8022 53333
rect 8078 53277 8146 53333
rect 8202 53277 8270 53333
rect 8326 53277 8394 53333
rect 8450 53277 8460 53333
rect 7640 53209 8460 53277
rect 7640 53153 7650 53209
rect 7706 53153 7774 53209
rect 7830 53153 7898 53209
rect 7954 53153 8022 53209
rect 8078 53153 8146 53209
rect 8202 53153 8270 53209
rect 8326 53153 8394 53209
rect 8450 53153 8460 53209
rect 7640 53085 8460 53153
rect 7640 53029 7650 53085
rect 7706 53029 7774 53085
rect 7830 53029 7898 53085
rect 7954 53029 8022 53085
rect 8078 53029 8146 53085
rect 8202 53029 8270 53085
rect 8326 53029 8394 53085
rect 8450 53029 8460 53085
rect 7640 52961 8460 53029
rect 7640 52905 7650 52961
rect 7706 52905 7774 52961
rect 7830 52905 7898 52961
rect 7954 52905 8022 52961
rect 8078 52905 8146 52961
rect 8202 52905 8270 52961
rect 8326 52905 8394 52961
rect 8450 52905 8460 52961
rect 7640 52837 8460 52905
rect 7640 52781 7650 52837
rect 7706 52781 7774 52837
rect 7830 52781 7898 52837
rect 7954 52781 8022 52837
rect 8078 52781 8146 52837
rect 8202 52781 8270 52837
rect 8326 52781 8394 52837
rect 8450 52781 8460 52837
rect 7640 52771 8460 52781
rect 8733 52737 9612 52826
rect 8733 52681 8812 52737
rect 8868 52681 8936 52737
rect 8992 52681 9060 52737
rect 9116 52681 9184 52737
rect 9240 52681 9308 52737
rect 9364 52681 9432 52737
rect 9488 52681 9612 52737
rect 8733 52613 9612 52681
rect 8733 52557 8812 52613
rect 8868 52557 8936 52613
rect 8992 52557 9060 52613
rect 9116 52557 9184 52613
rect 9240 52557 9308 52613
rect 9364 52557 9432 52613
rect 9488 52557 9612 52613
rect 8733 52489 9612 52557
rect 8733 52433 8812 52489
rect 8868 52433 8936 52489
rect 8992 52433 9060 52489
rect 9116 52433 9184 52489
rect 9240 52433 9308 52489
rect 9364 52433 9432 52489
rect 9488 52433 9612 52489
rect 8733 52365 9612 52433
rect 8733 52309 8812 52365
rect 8868 52309 8936 52365
rect 8992 52309 9060 52365
rect 9116 52309 9184 52365
rect 9240 52309 9308 52365
rect 9364 52309 9432 52365
rect 9488 52309 9612 52365
rect 8733 52241 9612 52309
rect 8733 52185 8812 52241
rect 8868 52185 8936 52241
rect 8992 52185 9060 52241
rect 9116 52185 9184 52241
rect 9240 52185 9308 52241
rect 9364 52185 9432 52241
rect 9488 52185 9612 52241
rect 8733 52117 9612 52185
rect 8733 52061 8812 52117
rect 8868 52061 8936 52117
rect 8992 52061 9060 52117
rect 9116 52061 9184 52117
rect 9240 52061 9308 52117
rect 9364 52061 9432 52117
rect 9488 52061 9612 52117
rect 8733 51993 9612 52061
rect 8733 51937 8812 51993
rect 8868 51937 8936 51993
rect 8992 51937 9060 51993
rect 9116 51937 9184 51993
rect 9240 51937 9308 51993
rect 9364 51937 9432 51993
rect 9488 51937 9612 51993
rect 8733 51869 9612 51937
rect 8733 51813 8812 51869
rect 8868 51813 8936 51869
rect 8992 51813 9060 51869
rect 9116 51813 9184 51869
rect 9240 51813 9308 51869
rect 9364 51813 9432 51869
rect 9488 51813 9612 51869
rect 8733 51745 9612 51813
rect 8733 51689 8812 51745
rect 8868 51689 8936 51745
rect 8992 51689 9060 51745
rect 9116 51689 9184 51745
rect 9240 51689 9308 51745
rect 9364 51689 9432 51745
rect 9488 51689 9612 51745
rect 8733 51621 9612 51689
rect 8733 51565 8812 51621
rect 8868 51565 8936 51621
rect 8992 51565 9060 51621
rect 9116 51565 9184 51621
rect 9240 51565 9308 51621
rect 9364 51565 9432 51621
rect 9488 51565 9612 51621
rect 7640 51452 8460 51462
rect 7640 51396 7650 51452
rect 7706 51396 7774 51452
rect 7830 51396 7898 51452
rect 7954 51396 8022 51452
rect 8078 51396 8146 51452
rect 8202 51396 8270 51452
rect 8326 51396 8394 51452
rect 8450 51396 8460 51452
rect 7640 51328 8460 51396
rect 7640 51272 7650 51328
rect 7706 51272 7774 51328
rect 7830 51272 7898 51328
rect 7954 51272 8022 51328
rect 8078 51272 8146 51328
rect 8202 51272 8270 51328
rect 8326 51272 8394 51328
rect 8450 51272 8460 51328
rect 7640 51204 8460 51272
rect 7640 51148 7650 51204
rect 7706 51148 7774 51204
rect 7830 51148 7898 51204
rect 7954 51148 8022 51204
rect 8078 51148 8146 51204
rect 8202 51148 8270 51204
rect 8326 51148 8394 51204
rect 8450 51148 8460 51204
rect 7640 51080 8460 51148
rect 7640 51024 7650 51080
rect 7706 51024 7774 51080
rect 7830 51024 7898 51080
rect 7954 51024 8022 51080
rect 8078 51024 8146 51080
rect 8202 51024 8270 51080
rect 8326 51024 8394 51080
rect 8450 51024 8460 51080
rect 7640 50956 8460 51024
rect 7640 50900 7650 50956
rect 7706 50900 7774 50956
rect 7830 50900 7898 50956
rect 7954 50900 8022 50956
rect 8078 50900 8146 50956
rect 8202 50900 8270 50956
rect 8326 50900 8394 50956
rect 8450 50900 8460 50956
rect 7640 50832 8460 50900
rect 7640 50776 7650 50832
rect 7706 50776 7774 50832
rect 7830 50776 7898 50832
rect 7954 50776 8022 50832
rect 8078 50776 8146 50832
rect 8202 50776 8270 50832
rect 8326 50776 8394 50832
rect 8450 50776 8460 50832
rect 7640 50708 8460 50776
rect 7640 50652 7650 50708
rect 7706 50652 7774 50708
rect 7830 50652 7898 50708
rect 7954 50652 8022 50708
rect 8078 50652 8146 50708
rect 8202 50652 8270 50708
rect 8326 50652 8394 50708
rect 8450 50652 8460 50708
rect 7640 50584 8460 50652
rect 7640 50528 7650 50584
rect 7706 50528 7774 50584
rect 7830 50528 7898 50584
rect 7954 50528 8022 50584
rect 8078 50528 8146 50584
rect 8202 50528 8270 50584
rect 8326 50528 8394 50584
rect 8450 50528 8460 50584
rect 7640 50518 8460 50528
rect 1094 42890 1170 42900
rect 1094 42834 1104 42890
rect 1160 42834 1170 42890
rect 1094 42766 1170 42834
rect 1094 42710 1104 42766
rect 1160 42710 1170 42766
rect 1094 42642 1170 42710
rect 1094 42586 1104 42642
rect 1160 42586 1170 42642
rect 1094 42518 1170 42586
rect 1094 42462 1104 42518
rect 1160 42462 1170 42518
rect 1094 42394 1170 42462
rect 1094 42338 1104 42394
rect 1160 42338 1170 42394
rect 1094 42270 1170 42338
rect 1094 42214 1104 42270
rect 1160 42214 1170 42270
rect 1094 42146 1170 42214
rect 1094 42090 1104 42146
rect 1160 42090 1170 42146
rect 1094 42022 1170 42090
rect 1094 41966 1104 42022
rect 1160 41966 1170 42022
rect 1094 41898 1170 41966
rect 1094 41842 1104 41898
rect 1160 41842 1170 41898
rect 1094 41774 1170 41842
rect 1094 41718 1104 41774
rect 1160 41718 1170 41774
rect 1094 41650 1170 41718
rect 1094 41594 1104 41650
rect 1160 41594 1170 41650
rect 1094 41526 1170 41594
rect 1094 41470 1104 41526
rect 1160 41470 1170 41526
rect 1094 41402 1170 41470
rect 1094 41346 1104 41402
rect 1160 41346 1170 41402
rect 1094 41278 1170 41346
rect 1094 41222 1104 41278
rect 1160 41222 1170 41278
rect 1094 41212 1170 41222
rect 1218 42766 1294 42776
rect 1218 42710 1228 42766
rect 1284 42710 1294 42766
rect 1218 42642 1294 42710
rect 1218 42586 1228 42642
rect 1284 42586 1294 42642
rect 1218 42518 1294 42586
rect 1218 42462 1228 42518
rect 1284 42462 1294 42518
rect 1218 42394 1294 42462
rect 1218 42338 1228 42394
rect 1284 42338 1294 42394
rect 1218 42270 1294 42338
rect 1218 42214 1228 42270
rect 1284 42214 1294 42270
rect 1218 42146 1294 42214
rect 1218 42090 1228 42146
rect 1284 42090 1294 42146
rect 1218 42022 1294 42090
rect 1218 41966 1228 42022
rect 1284 41966 1294 42022
rect 1218 41898 1294 41966
rect 1218 41842 1228 41898
rect 1284 41842 1294 41898
rect 1218 41774 1294 41842
rect 1218 41718 1228 41774
rect 1284 41718 1294 41774
rect 1218 41650 1294 41718
rect 1218 41594 1228 41650
rect 1284 41594 1294 41650
rect 1218 41526 1294 41594
rect 1218 41470 1228 41526
rect 1284 41470 1294 41526
rect 1218 41402 1294 41470
rect 1218 41346 1228 41402
rect 1284 41346 1294 41402
rect 1218 41278 1294 41346
rect 1218 41222 1228 41278
rect 1284 41222 1294 41278
rect 1218 41154 1294 41222
rect 1218 41098 1228 41154
rect 1284 41098 1294 41154
rect 1218 41088 1294 41098
rect 1342 42642 1418 42652
rect 1342 42586 1352 42642
rect 1408 42586 1418 42642
rect 1342 42518 1418 42586
rect 1342 42462 1352 42518
rect 1408 42462 1418 42518
rect 1342 42394 1418 42462
rect 1342 42338 1352 42394
rect 1408 42338 1418 42394
rect 1342 42270 1418 42338
rect 1342 42214 1352 42270
rect 1408 42214 1418 42270
rect 1342 42146 1418 42214
rect 1342 42090 1352 42146
rect 1408 42090 1418 42146
rect 1342 42022 1418 42090
rect 1342 41966 1352 42022
rect 1408 41966 1418 42022
rect 1342 41898 1418 41966
rect 1342 41842 1352 41898
rect 1408 41842 1418 41898
rect 1342 41774 1418 41842
rect 1342 41718 1352 41774
rect 1408 41718 1418 41774
rect 1342 41650 1418 41718
rect 1342 41594 1352 41650
rect 1408 41594 1418 41650
rect 1342 41526 1418 41594
rect 1342 41470 1352 41526
rect 1408 41470 1418 41526
rect 1342 41402 1418 41470
rect 1342 41346 1352 41402
rect 1408 41346 1418 41402
rect 1342 41278 1418 41346
rect 1342 41222 1352 41278
rect 1408 41222 1418 41278
rect 1342 41154 1418 41222
rect 1342 41098 1352 41154
rect 1408 41098 1418 41154
rect 1342 41030 1418 41098
rect 1342 40974 1352 41030
rect 1408 40974 1418 41030
rect 1342 40964 1418 40974
rect 1466 42518 1542 42528
rect 1466 42462 1476 42518
rect 1532 42462 1542 42518
rect 1466 42394 1542 42462
rect 1466 42338 1476 42394
rect 1532 42338 1542 42394
rect 1466 42270 1542 42338
rect 1466 42214 1476 42270
rect 1532 42214 1542 42270
rect 1466 42146 1542 42214
rect 1466 42090 1476 42146
rect 1532 42090 1542 42146
rect 1466 42022 1542 42090
rect 1466 41966 1476 42022
rect 1532 41966 1542 42022
rect 1466 41898 1542 41966
rect 1466 41842 1476 41898
rect 1532 41842 1542 41898
rect 1466 41774 1542 41842
rect 1466 41718 1476 41774
rect 1532 41718 1542 41774
rect 1466 41650 1542 41718
rect 1466 41594 1476 41650
rect 1532 41594 1542 41650
rect 1466 41526 1542 41594
rect 1466 41470 1476 41526
rect 1532 41470 1542 41526
rect 1466 41402 1542 41470
rect 1466 41346 1476 41402
rect 1532 41346 1542 41402
rect 1466 41278 1542 41346
rect 1466 41222 1476 41278
rect 1532 41222 1542 41278
rect 1466 41154 1542 41222
rect 1466 41098 1476 41154
rect 1532 41098 1542 41154
rect 1466 41030 1542 41098
rect 1466 40974 1476 41030
rect 1532 40974 1542 41030
rect 1466 40906 1542 40974
rect 1466 40850 1476 40906
rect 1532 40850 1542 40906
rect 1466 40840 1542 40850
rect 1590 42394 1666 42404
rect 1590 42338 1600 42394
rect 1656 42338 1666 42394
rect 1590 42270 1666 42338
rect 1590 42214 1600 42270
rect 1656 42214 1666 42270
rect 1590 42146 1666 42214
rect 1590 42090 1600 42146
rect 1656 42090 1666 42146
rect 1590 42022 1666 42090
rect 1590 41966 1600 42022
rect 1656 41966 1666 42022
rect 1590 41898 1666 41966
rect 1590 41842 1600 41898
rect 1656 41842 1666 41898
rect 1590 41774 1666 41842
rect 1590 41718 1600 41774
rect 1656 41718 1666 41774
rect 1590 41650 1666 41718
rect 1590 41594 1600 41650
rect 1656 41594 1666 41650
rect 1590 41526 1666 41594
rect 1590 41470 1600 41526
rect 1656 41470 1666 41526
rect 1590 41402 1666 41470
rect 1590 41346 1600 41402
rect 1656 41346 1666 41402
rect 1590 41278 1666 41346
rect 1590 41222 1600 41278
rect 1656 41222 1666 41278
rect 1590 41154 1666 41222
rect 1590 41098 1600 41154
rect 1656 41098 1666 41154
rect 1590 41030 1666 41098
rect 1590 40974 1600 41030
rect 1656 40974 1666 41030
rect 1590 40906 1666 40974
rect 1590 40850 1600 40906
rect 1656 40850 1666 40906
rect 1590 40782 1666 40850
rect 1590 40726 1600 40782
rect 1656 40726 1666 40782
rect 1590 40716 1666 40726
rect 1714 42270 1790 42280
rect 1714 42214 1724 42270
rect 1780 42214 1790 42270
rect 1714 42146 1790 42214
rect 1714 42090 1724 42146
rect 1780 42090 1790 42146
rect 1714 42022 1790 42090
rect 1714 41966 1724 42022
rect 1780 41966 1790 42022
rect 1714 41898 1790 41966
rect 1714 41842 1724 41898
rect 1780 41842 1790 41898
rect 1714 41774 1790 41842
rect 1714 41718 1724 41774
rect 1780 41718 1790 41774
rect 1714 41650 1790 41718
rect 1714 41594 1724 41650
rect 1780 41594 1790 41650
rect 1714 41526 1790 41594
rect 1714 41470 1724 41526
rect 1780 41470 1790 41526
rect 1714 41402 1790 41470
rect 1714 41346 1724 41402
rect 1780 41346 1790 41402
rect 1714 41278 1790 41346
rect 1714 41222 1724 41278
rect 1780 41222 1790 41278
rect 1714 41154 1790 41222
rect 1714 41098 1724 41154
rect 1780 41098 1790 41154
rect 1714 41030 1790 41098
rect 1714 40974 1724 41030
rect 1780 40974 1790 41030
rect 1714 40906 1790 40974
rect 1714 40850 1724 40906
rect 1780 40850 1790 40906
rect 1714 40782 1790 40850
rect 1714 40726 1724 40782
rect 1780 40726 1790 40782
rect 1714 40658 1790 40726
rect 1714 40602 1724 40658
rect 1780 40602 1790 40658
rect 1714 40592 1790 40602
rect 1838 42146 1914 42156
rect 1838 42090 1848 42146
rect 1904 42090 1914 42146
rect 1838 42022 1914 42090
rect 1838 41966 1848 42022
rect 1904 41966 1914 42022
rect 1838 41898 1914 41966
rect 1838 41842 1848 41898
rect 1904 41842 1914 41898
rect 1838 41774 1914 41842
rect 1838 41718 1848 41774
rect 1904 41718 1914 41774
rect 1838 41650 1914 41718
rect 1838 41594 1848 41650
rect 1904 41594 1914 41650
rect 1838 41526 1914 41594
rect 1838 41470 1848 41526
rect 1904 41470 1914 41526
rect 1838 41402 1914 41470
rect 1838 41346 1848 41402
rect 1904 41346 1914 41402
rect 1838 41278 1914 41346
rect 1838 41222 1848 41278
rect 1904 41222 1914 41278
rect 1838 41154 1914 41222
rect 1838 41098 1848 41154
rect 1904 41098 1914 41154
rect 1838 41030 1914 41098
rect 1838 40974 1848 41030
rect 1904 40974 1914 41030
rect 1838 40906 1914 40974
rect 1838 40850 1848 40906
rect 1904 40850 1914 40906
rect 1838 40782 1914 40850
rect 1838 40726 1848 40782
rect 1904 40726 1914 40782
rect 1838 40658 1914 40726
rect 1838 40602 1848 40658
rect 1904 40602 1914 40658
rect 1838 40534 1914 40602
rect 1838 40478 1848 40534
rect 1904 40478 1914 40534
rect 1838 40468 1914 40478
rect 1962 42022 2038 42032
rect 1962 41966 1972 42022
rect 2028 41966 2038 42022
rect 1962 41898 2038 41966
rect 1962 41842 1972 41898
rect 2028 41842 2038 41898
rect 1962 41774 2038 41842
rect 1962 41718 1972 41774
rect 2028 41718 2038 41774
rect 1962 41650 2038 41718
rect 8733 41714 9612 51565
rect 13707 50948 13910 50992
rect 12842 50938 13910 50948
rect 12842 50882 12852 50938
rect 12908 50882 12976 50938
rect 13032 50882 13100 50938
rect 13156 50882 13224 50938
rect 13280 50882 13348 50938
rect 13404 50882 13472 50938
rect 13528 50882 13596 50938
rect 13652 50882 13720 50938
rect 13776 50882 13844 50938
rect 13900 50882 13910 50938
rect 12842 50814 13910 50882
rect 12842 50758 12852 50814
rect 12908 50758 12976 50814
rect 13032 50758 13100 50814
rect 13156 50758 13224 50814
rect 13280 50758 13348 50814
rect 13404 50758 13472 50814
rect 13528 50758 13596 50814
rect 13652 50758 13720 50814
rect 13776 50758 13844 50814
rect 13900 50758 13910 50814
rect 12842 50690 13910 50758
rect 12842 50634 12852 50690
rect 12908 50634 12976 50690
rect 13032 50634 13100 50690
rect 13156 50634 13224 50690
rect 13280 50634 13348 50690
rect 13404 50634 13472 50690
rect 13528 50634 13596 50690
rect 13652 50634 13720 50690
rect 13776 50634 13844 50690
rect 13900 50634 13910 50690
rect 12842 50566 13910 50634
rect 12842 50510 12852 50566
rect 12908 50510 12976 50566
rect 13032 50510 13100 50566
rect 13156 50510 13224 50566
rect 13280 50510 13348 50566
rect 13404 50510 13472 50566
rect 13528 50510 13596 50566
rect 13652 50510 13720 50566
rect 13776 50510 13844 50566
rect 13900 50510 13910 50566
rect 12842 50442 13910 50510
rect 12842 50386 12852 50442
rect 12908 50386 12976 50442
rect 13032 50386 13100 50442
rect 13156 50386 13224 50442
rect 13280 50386 13348 50442
rect 13404 50386 13472 50442
rect 13528 50386 13596 50442
rect 13652 50386 13720 50442
rect 13776 50386 13844 50442
rect 13900 50386 13910 50442
rect 12842 50318 13910 50386
rect 12842 50262 12852 50318
rect 12908 50262 12976 50318
rect 13032 50262 13100 50318
rect 13156 50262 13224 50318
rect 13280 50262 13348 50318
rect 13404 50262 13472 50318
rect 13528 50262 13596 50318
rect 13652 50262 13720 50318
rect 13776 50262 13844 50318
rect 13900 50262 13910 50318
rect 12842 50194 13910 50262
rect 12842 50138 12852 50194
rect 12908 50138 12976 50194
rect 13032 50138 13100 50194
rect 13156 50138 13224 50194
rect 13280 50138 13348 50194
rect 13404 50138 13472 50194
rect 13528 50138 13596 50194
rect 13652 50138 13720 50194
rect 13776 50138 13844 50194
rect 13900 50138 13910 50194
rect 12842 50070 13910 50138
rect 12842 50014 12852 50070
rect 12908 50014 12976 50070
rect 13032 50014 13100 50070
rect 13156 50014 13224 50070
rect 13280 50014 13348 50070
rect 13404 50014 13472 50070
rect 13528 50014 13596 50070
rect 13652 50014 13720 50070
rect 13776 50014 13844 50070
rect 13900 50014 13910 50070
rect 12842 49946 13910 50014
rect 12842 49890 12852 49946
rect 12908 49890 12976 49946
rect 13032 49890 13100 49946
rect 13156 49890 13224 49946
rect 13280 49890 13348 49946
rect 13404 49890 13472 49946
rect 13528 49890 13596 49946
rect 13652 49890 13720 49946
rect 13776 49890 13844 49946
rect 13900 49890 13910 49946
rect 12842 49822 13910 49890
rect 12842 49766 12852 49822
rect 12908 49766 12976 49822
rect 13032 49766 13100 49822
rect 13156 49766 13224 49822
rect 13280 49766 13348 49822
rect 13404 49766 13472 49822
rect 13528 49766 13596 49822
rect 13652 49766 13720 49822
rect 13776 49766 13844 49822
rect 13900 49766 13910 49822
rect 12842 49698 13910 49766
rect 12842 49642 12852 49698
rect 12908 49642 12976 49698
rect 13032 49642 13100 49698
rect 13156 49642 13224 49698
rect 13280 49642 13348 49698
rect 13404 49642 13472 49698
rect 13528 49642 13596 49698
rect 13652 49642 13720 49698
rect 13776 49642 13844 49698
rect 13900 49642 13910 49698
rect 12842 49632 13910 49642
rect 13707 49592 13910 49632
rect 14757 50972 14833 50982
rect 14757 49620 14767 50972
rect 14823 49620 14833 50972
rect 14757 49610 14833 49620
rect 10638 49356 10996 49392
rect 10638 49346 12481 49356
rect 10638 49290 10679 49346
rect 10735 49290 10803 49346
rect 10859 49290 10927 49346
rect 10983 49290 11051 49346
rect 11107 49290 11175 49346
rect 11231 49290 11299 49346
rect 11355 49290 11423 49346
rect 11479 49290 11547 49346
rect 11603 49290 11671 49346
rect 11727 49290 11795 49346
rect 11851 49290 11919 49346
rect 11975 49290 12043 49346
rect 12099 49290 12167 49346
rect 12223 49290 12291 49346
rect 12347 49290 12415 49346
rect 12471 49290 12481 49346
rect 10638 49222 12481 49290
rect 10638 49166 10679 49222
rect 10735 49166 10803 49222
rect 10859 49166 10927 49222
rect 10983 49166 11051 49222
rect 11107 49166 11175 49222
rect 11231 49166 11299 49222
rect 11355 49166 11423 49222
rect 11479 49166 11547 49222
rect 11603 49166 11671 49222
rect 11727 49166 11795 49222
rect 11851 49166 11919 49222
rect 11975 49166 12043 49222
rect 12099 49166 12167 49222
rect 12223 49166 12291 49222
rect 12347 49166 12415 49222
rect 12471 49166 12481 49222
rect 10638 49098 12481 49166
rect 10638 49042 10679 49098
rect 10735 49042 10803 49098
rect 10859 49042 10927 49098
rect 10983 49042 11051 49098
rect 11107 49042 11175 49098
rect 11231 49042 11299 49098
rect 11355 49042 11423 49098
rect 11479 49042 11547 49098
rect 11603 49042 11671 49098
rect 11727 49042 11795 49098
rect 11851 49042 11919 49098
rect 11975 49042 12043 49098
rect 12099 49042 12167 49098
rect 12223 49042 12291 49098
rect 12347 49042 12415 49098
rect 12471 49042 12481 49098
rect 10638 48974 12481 49042
rect 10638 48918 10679 48974
rect 10735 48918 10803 48974
rect 10859 48918 10927 48974
rect 10983 48918 11051 48974
rect 11107 48918 11175 48974
rect 11231 48918 11299 48974
rect 11355 48918 11423 48974
rect 11479 48918 11547 48974
rect 11603 48918 11671 48974
rect 11727 48918 11795 48974
rect 11851 48918 11919 48974
rect 11975 48918 12043 48974
rect 12099 48918 12167 48974
rect 12223 48918 12291 48974
rect 12347 48918 12415 48974
rect 12471 48918 12481 48974
rect 10638 48850 12481 48918
rect 10638 48794 10679 48850
rect 10735 48794 10803 48850
rect 10859 48794 10927 48850
rect 10983 48794 11051 48850
rect 11107 48794 11175 48850
rect 11231 48794 11299 48850
rect 11355 48794 11423 48850
rect 11479 48794 11547 48850
rect 11603 48794 11671 48850
rect 11727 48794 11795 48850
rect 11851 48794 11919 48850
rect 11975 48794 12043 48850
rect 12099 48794 12167 48850
rect 12223 48794 12291 48850
rect 12347 48794 12415 48850
rect 12471 48794 12481 48850
rect 10638 48726 12481 48794
rect 10638 48670 10679 48726
rect 10735 48670 10803 48726
rect 10859 48670 10927 48726
rect 10983 48670 11051 48726
rect 11107 48670 11175 48726
rect 11231 48670 11299 48726
rect 11355 48670 11423 48726
rect 11479 48670 11547 48726
rect 11603 48670 11671 48726
rect 11727 48670 11795 48726
rect 11851 48670 11919 48726
rect 11975 48670 12043 48726
rect 12099 48670 12167 48726
rect 12223 48670 12291 48726
rect 12347 48670 12415 48726
rect 12471 48670 12481 48726
rect 10638 48602 12481 48670
rect 10638 48546 10679 48602
rect 10735 48546 10803 48602
rect 10859 48546 10927 48602
rect 10983 48546 11051 48602
rect 11107 48546 11175 48602
rect 11231 48546 11299 48602
rect 11355 48546 11423 48602
rect 11479 48546 11547 48602
rect 11603 48546 11671 48602
rect 11727 48546 11795 48602
rect 11851 48546 11919 48602
rect 11975 48546 12043 48602
rect 12099 48546 12167 48602
rect 12223 48546 12291 48602
rect 12347 48546 12415 48602
rect 12471 48546 12481 48602
rect 10638 48478 12481 48546
rect 10638 48422 10679 48478
rect 10735 48422 10803 48478
rect 10859 48422 10927 48478
rect 10983 48422 11051 48478
rect 11107 48422 11175 48478
rect 11231 48422 11299 48478
rect 11355 48422 11423 48478
rect 11479 48422 11547 48478
rect 11603 48422 11671 48478
rect 11727 48422 11795 48478
rect 11851 48422 11919 48478
rect 11975 48422 12043 48478
rect 12099 48422 12167 48478
rect 12223 48422 12291 48478
rect 12347 48422 12415 48478
rect 12471 48422 12481 48478
rect 10638 48354 12481 48422
rect 10638 48298 10679 48354
rect 10735 48298 10803 48354
rect 10859 48298 10927 48354
rect 10983 48298 11051 48354
rect 11107 48298 11175 48354
rect 11231 48298 11299 48354
rect 11355 48298 11423 48354
rect 11479 48298 11547 48354
rect 11603 48298 11671 48354
rect 11727 48298 11795 48354
rect 11851 48298 11919 48354
rect 11975 48298 12043 48354
rect 12099 48298 12167 48354
rect 12223 48298 12291 48354
rect 12347 48298 12415 48354
rect 12471 48298 12481 48354
rect 10638 48230 12481 48298
rect 10638 48174 10679 48230
rect 10735 48174 10803 48230
rect 10859 48174 10927 48230
rect 10983 48174 11051 48230
rect 11107 48174 11175 48230
rect 11231 48174 11299 48230
rect 11355 48174 11423 48230
rect 11479 48174 11547 48230
rect 11603 48174 11671 48230
rect 11727 48174 11795 48230
rect 11851 48174 11919 48230
rect 11975 48174 12043 48230
rect 12099 48174 12167 48230
rect 12223 48174 12291 48230
rect 12347 48174 12415 48230
rect 12471 48174 12481 48230
rect 10638 48106 12481 48174
rect 10638 48050 10679 48106
rect 10735 48050 10803 48106
rect 10859 48050 10927 48106
rect 10983 48050 11051 48106
rect 11107 48050 11175 48106
rect 11231 48050 11299 48106
rect 11355 48050 11423 48106
rect 11479 48050 11547 48106
rect 11603 48050 11671 48106
rect 11727 48050 11795 48106
rect 11851 48050 11919 48106
rect 11975 48050 12043 48106
rect 12099 48050 12167 48106
rect 12223 48050 12291 48106
rect 12347 48050 12415 48106
rect 12471 48050 12481 48106
rect 10638 48040 12481 48050
rect 10638 47992 10996 48040
rect 1962 41594 1972 41650
rect 2028 41594 2038 41650
rect 1962 41526 2038 41594
rect 1962 41470 1972 41526
rect 2028 41470 2038 41526
rect 1962 41402 2038 41470
rect 1962 41346 1972 41402
rect 2028 41346 2038 41402
rect 1962 41278 2038 41346
rect 1962 41222 1972 41278
rect 2028 41222 2038 41278
rect 1962 41154 2038 41222
rect 1962 41098 1972 41154
rect 2028 41098 2038 41154
rect 1962 41030 2038 41098
rect 1962 40974 1972 41030
rect 2028 40974 2038 41030
rect 1962 40906 2038 40974
rect 1962 40850 1972 40906
rect 2028 40850 2038 40906
rect 1962 40782 2038 40850
rect 1962 40726 1972 40782
rect 2028 40726 2038 40782
rect 1962 40658 2038 40726
rect 1962 40602 1972 40658
rect 2028 40602 2038 40658
rect 1962 40534 2038 40602
rect 1962 40478 1972 40534
rect 2028 40478 2038 40534
rect 1962 40410 2038 40478
rect 1962 40354 1972 40410
rect 2028 40354 2038 40410
rect 1962 40344 2038 40354
rect 4460 39524 4536 39534
rect 4460 39468 4470 39524
rect 4526 39468 4536 39524
rect 4460 39400 4536 39468
rect 4460 39344 4470 39400
rect 4526 39344 4536 39400
rect 4460 39276 4536 39344
rect 4460 39220 4470 39276
rect 4526 39220 4536 39276
rect 2517 39205 2593 39215
rect 2517 39149 2527 39205
rect 2583 39149 2593 39205
rect 2517 39081 2593 39149
rect 4460 39152 4536 39220
rect 4460 39096 4470 39152
rect 4526 39096 4536 39152
rect 2517 39025 2527 39081
rect 2583 39025 2593 39081
rect 2517 38957 2593 39025
rect 2517 38901 2527 38957
rect 2583 38901 2593 38957
rect 2517 38833 2593 38901
rect 2517 38777 2527 38833
rect 2583 38777 2593 38833
rect 2517 38709 2593 38777
rect 2517 38653 2527 38709
rect 2583 38653 2593 38709
rect 2517 38585 2593 38653
rect 2517 38529 2527 38585
rect 2583 38529 2593 38585
rect 2517 38461 2593 38529
rect 2517 38405 2527 38461
rect 2583 38405 2593 38461
rect 2517 38337 2593 38405
rect 2517 38281 2527 38337
rect 2583 38281 2593 38337
rect 2517 38213 2593 38281
rect 2517 38157 2527 38213
rect 2583 38157 2593 38213
rect 2517 38089 2593 38157
rect 2517 38033 2527 38089
rect 2583 38033 2593 38089
rect 2517 37965 2593 38033
rect 2517 37909 2527 37965
rect 2583 37909 2593 37965
rect 2517 37841 2593 37909
rect 2517 37785 2527 37841
rect 2583 37785 2593 37841
rect 2517 37717 2593 37785
rect 2517 37661 2527 37717
rect 2583 37661 2593 37717
rect 2517 37593 2593 37661
rect 2517 37537 2527 37593
rect 2583 37537 2593 37593
rect 2517 37527 2593 37537
rect 2641 39081 2717 39091
rect 2641 39025 2651 39081
rect 2707 39025 2717 39081
rect 2641 38957 2717 39025
rect 4460 39028 4536 39096
rect 4460 38972 4470 39028
rect 4526 38972 4536 39028
rect 2641 38901 2651 38957
rect 2707 38901 2717 38957
rect 2641 38833 2717 38901
rect 2641 38777 2651 38833
rect 2707 38777 2717 38833
rect 2641 38709 2717 38777
rect 2641 38653 2651 38709
rect 2707 38653 2717 38709
rect 2641 38585 2717 38653
rect 2641 38529 2651 38585
rect 2707 38529 2717 38585
rect 2641 38461 2717 38529
rect 2641 38405 2651 38461
rect 2707 38405 2717 38461
rect 2641 38337 2717 38405
rect 2641 38281 2651 38337
rect 2707 38281 2717 38337
rect 2641 38213 2717 38281
rect 2641 38157 2651 38213
rect 2707 38157 2717 38213
rect 2641 38089 2717 38157
rect 2641 38033 2651 38089
rect 2707 38033 2717 38089
rect 2641 37965 2717 38033
rect 2641 37909 2651 37965
rect 2707 37909 2717 37965
rect 2641 37841 2717 37909
rect 2641 37785 2651 37841
rect 2707 37785 2717 37841
rect 2641 37717 2717 37785
rect 2641 37661 2651 37717
rect 2707 37661 2717 37717
rect 2641 37593 2717 37661
rect 2641 37537 2651 37593
rect 2707 37537 2717 37593
rect 2641 37469 2717 37537
rect 2641 37413 2651 37469
rect 2707 37413 2717 37469
rect 2641 37403 2717 37413
rect 2765 38957 2841 38967
rect 2765 38901 2775 38957
rect 2831 38901 2841 38957
rect 2765 38833 2841 38901
rect 4460 38904 4536 38972
rect 4460 38848 4470 38904
rect 4526 38848 4536 38904
rect 2765 38777 2775 38833
rect 2831 38777 2841 38833
rect 2765 38709 2841 38777
rect 2765 38653 2775 38709
rect 2831 38653 2841 38709
rect 2765 38585 2841 38653
rect 2765 38529 2775 38585
rect 2831 38529 2841 38585
rect 2765 38461 2841 38529
rect 2765 38405 2775 38461
rect 2831 38405 2841 38461
rect 2765 38337 2841 38405
rect 2765 38281 2775 38337
rect 2831 38281 2841 38337
rect 2765 38213 2841 38281
rect 2765 38157 2775 38213
rect 2831 38157 2841 38213
rect 2765 38089 2841 38157
rect 2765 38033 2775 38089
rect 2831 38033 2841 38089
rect 2765 37965 2841 38033
rect 2765 37909 2775 37965
rect 2831 37909 2841 37965
rect 2765 37841 2841 37909
rect 2765 37785 2775 37841
rect 2831 37785 2841 37841
rect 2765 37717 2841 37785
rect 2765 37661 2775 37717
rect 2831 37661 2841 37717
rect 2765 37593 2841 37661
rect 2765 37537 2775 37593
rect 2831 37537 2841 37593
rect 2765 37469 2841 37537
rect 2765 37413 2775 37469
rect 2831 37413 2841 37469
rect 2765 37345 2841 37413
rect 2765 37289 2775 37345
rect 2831 37289 2841 37345
rect 2765 37279 2841 37289
rect 2889 38833 2965 38843
rect 2889 38777 2899 38833
rect 2955 38777 2965 38833
rect 2889 38709 2965 38777
rect 4460 38780 4536 38848
rect 4460 38724 4470 38780
rect 4526 38724 4536 38780
rect 2889 38653 2899 38709
rect 2955 38653 2965 38709
rect 2889 38585 2965 38653
rect 2889 38529 2899 38585
rect 2955 38529 2965 38585
rect 2889 38461 2965 38529
rect 2889 38405 2899 38461
rect 2955 38405 2965 38461
rect 2889 38337 2965 38405
rect 2889 38281 2899 38337
rect 2955 38281 2965 38337
rect 2889 38213 2965 38281
rect 2889 38157 2899 38213
rect 2955 38157 2965 38213
rect 2889 38089 2965 38157
rect 2889 38033 2899 38089
rect 2955 38033 2965 38089
rect 2889 37965 2965 38033
rect 2889 37909 2899 37965
rect 2955 37909 2965 37965
rect 2889 37841 2965 37909
rect 2889 37785 2899 37841
rect 2955 37785 2965 37841
rect 2889 37717 2965 37785
rect 2889 37661 2899 37717
rect 2955 37661 2965 37717
rect 2889 37593 2965 37661
rect 2889 37537 2899 37593
rect 2955 37537 2965 37593
rect 2889 37469 2965 37537
rect 2889 37413 2899 37469
rect 2955 37413 2965 37469
rect 2889 37345 2965 37413
rect 2889 37289 2899 37345
rect 2955 37289 2965 37345
rect 2889 37221 2965 37289
rect 2889 37165 2899 37221
rect 2955 37165 2965 37221
rect 2889 37155 2965 37165
rect 3013 38709 3089 38719
rect 3013 38653 3023 38709
rect 3079 38653 3089 38709
rect 3013 38585 3089 38653
rect 4460 38656 4536 38724
rect 4460 38600 4470 38656
rect 4526 38600 4536 38656
rect 3013 38529 3023 38585
rect 3079 38529 3089 38585
rect 3013 38461 3089 38529
rect 3013 38405 3023 38461
rect 3079 38405 3089 38461
rect 3013 38337 3089 38405
rect 3013 38281 3023 38337
rect 3079 38281 3089 38337
rect 3013 38213 3089 38281
rect 3013 38157 3023 38213
rect 3079 38157 3089 38213
rect 3013 38089 3089 38157
rect 3013 38033 3023 38089
rect 3079 38033 3089 38089
rect 3013 37965 3089 38033
rect 3013 37909 3023 37965
rect 3079 37909 3089 37965
rect 3013 37841 3089 37909
rect 3013 37785 3023 37841
rect 3079 37785 3089 37841
rect 3013 37717 3089 37785
rect 3013 37661 3023 37717
rect 3079 37661 3089 37717
rect 3013 37593 3089 37661
rect 3013 37537 3023 37593
rect 3079 37537 3089 37593
rect 3013 37469 3089 37537
rect 3013 37413 3023 37469
rect 3079 37413 3089 37469
rect 3013 37345 3089 37413
rect 3013 37289 3023 37345
rect 3079 37289 3089 37345
rect 3013 37221 3089 37289
rect 3013 37165 3023 37221
rect 3079 37165 3089 37221
rect 3013 37097 3089 37165
rect 3013 37041 3023 37097
rect 3079 37041 3089 37097
rect 3013 37031 3089 37041
rect 3137 38585 3213 38595
rect 3137 38529 3147 38585
rect 3203 38529 3213 38585
rect 3137 38461 3213 38529
rect 4460 38532 4536 38600
rect 4460 38476 4470 38532
rect 4526 38476 4536 38532
rect 3137 38405 3147 38461
rect 3203 38405 3213 38461
rect 3137 38337 3213 38405
rect 3137 38281 3147 38337
rect 3203 38281 3213 38337
rect 3137 38213 3213 38281
rect 3137 38157 3147 38213
rect 3203 38157 3213 38213
rect 3137 38089 3213 38157
rect 3137 38033 3147 38089
rect 3203 38033 3213 38089
rect 3137 37965 3213 38033
rect 3137 37909 3147 37965
rect 3203 37909 3213 37965
rect 3137 37841 3213 37909
rect 3137 37785 3147 37841
rect 3203 37785 3213 37841
rect 3137 37717 3213 37785
rect 3137 37661 3147 37717
rect 3203 37661 3213 37717
rect 3137 37593 3213 37661
rect 3137 37537 3147 37593
rect 3203 37537 3213 37593
rect 3137 37469 3213 37537
rect 3137 37413 3147 37469
rect 3203 37413 3213 37469
rect 3137 37345 3213 37413
rect 3137 37289 3147 37345
rect 3203 37289 3213 37345
rect 3137 37221 3213 37289
rect 3137 37165 3147 37221
rect 3203 37165 3213 37221
rect 3137 37097 3213 37165
rect 3137 37041 3147 37097
rect 3203 37041 3213 37097
rect 3137 36973 3213 37041
rect 3137 36917 3147 36973
rect 3203 36917 3213 36973
rect 3137 36907 3213 36917
rect 3261 38461 3337 38471
rect 3261 38405 3271 38461
rect 3327 38405 3337 38461
rect 3261 38337 3337 38405
rect 4460 38408 4536 38476
rect 4460 38352 4470 38408
rect 4526 38352 4536 38408
rect 3261 38281 3271 38337
rect 3327 38281 3337 38337
rect 3261 38213 3337 38281
rect 3261 38157 3271 38213
rect 3327 38157 3337 38213
rect 3261 38089 3337 38157
rect 3261 38033 3271 38089
rect 3327 38033 3337 38089
rect 3261 37965 3337 38033
rect 3261 37909 3271 37965
rect 3327 37909 3337 37965
rect 3261 37841 3337 37909
rect 3261 37785 3271 37841
rect 3327 37785 3337 37841
rect 3261 37717 3337 37785
rect 3261 37661 3271 37717
rect 3327 37661 3337 37717
rect 3261 37593 3337 37661
rect 3261 37537 3271 37593
rect 3327 37537 3337 37593
rect 3261 37469 3337 37537
rect 3261 37413 3271 37469
rect 3327 37413 3337 37469
rect 3261 37345 3337 37413
rect 3261 37289 3271 37345
rect 3327 37289 3337 37345
rect 3261 37221 3337 37289
rect 3261 37165 3271 37221
rect 3327 37165 3337 37221
rect 3261 37097 3337 37165
rect 3261 37041 3271 37097
rect 3327 37041 3337 37097
rect 3261 36973 3337 37041
rect 3261 36917 3271 36973
rect 3327 36917 3337 36973
rect 3261 36849 3337 36917
rect 3261 36793 3271 36849
rect 3327 36793 3337 36849
rect 3261 36783 3337 36793
rect 3385 38337 3461 38347
rect 3385 38281 3395 38337
rect 3451 38281 3461 38337
rect 3385 38213 3461 38281
rect 4460 38284 4536 38352
rect 4460 38228 4470 38284
rect 4526 38228 4536 38284
rect 3385 38157 3395 38213
rect 3451 38157 3461 38213
rect 3385 38089 3461 38157
rect 3385 38033 3395 38089
rect 3451 38033 3461 38089
rect 3385 37965 3461 38033
rect 3385 37909 3395 37965
rect 3451 37909 3461 37965
rect 3385 37841 3461 37909
rect 3385 37785 3395 37841
rect 3451 37785 3461 37841
rect 3385 37717 3461 37785
rect 3385 37661 3395 37717
rect 3451 37661 3461 37717
rect 3385 37593 3461 37661
rect 3385 37537 3395 37593
rect 3451 37537 3461 37593
rect 3385 37469 3461 37537
rect 3385 37413 3395 37469
rect 3451 37413 3461 37469
rect 3385 37345 3461 37413
rect 3385 37289 3395 37345
rect 3451 37289 3461 37345
rect 3385 37221 3461 37289
rect 3385 37165 3395 37221
rect 3451 37165 3461 37221
rect 3385 37097 3461 37165
rect 3385 37041 3395 37097
rect 3451 37041 3461 37097
rect 3385 36973 3461 37041
rect 3385 36917 3395 36973
rect 3451 36917 3461 36973
rect 3385 36849 3461 36917
rect 3385 36793 3395 36849
rect 3451 36793 3461 36849
rect 3385 36725 3461 36793
rect 3385 36669 3395 36725
rect 3451 36669 3461 36725
rect 3385 36659 3461 36669
rect 3509 38213 3585 38223
rect 3509 38157 3519 38213
rect 3575 38157 3585 38213
rect 3509 38089 3585 38157
rect 4460 38160 4536 38228
rect 4460 38104 4470 38160
rect 4526 38104 4536 38160
rect 3509 38033 3519 38089
rect 3575 38033 3585 38089
rect 3509 37965 3585 38033
rect 3509 37909 3519 37965
rect 3575 37909 3585 37965
rect 3509 37841 3585 37909
rect 3509 37785 3519 37841
rect 3575 37785 3585 37841
rect 3509 37717 3585 37785
rect 3509 37661 3519 37717
rect 3575 37661 3585 37717
rect 3509 37593 3585 37661
rect 3509 37537 3519 37593
rect 3575 37537 3585 37593
rect 3509 37469 3585 37537
rect 3509 37413 3519 37469
rect 3575 37413 3585 37469
rect 3509 37345 3585 37413
rect 3509 37289 3519 37345
rect 3575 37289 3585 37345
rect 3509 37221 3585 37289
rect 3509 37165 3519 37221
rect 3575 37165 3585 37221
rect 3509 37097 3585 37165
rect 3509 37041 3519 37097
rect 3575 37041 3585 37097
rect 3509 36973 3585 37041
rect 3509 36917 3519 36973
rect 3575 36917 3585 36973
rect 3509 36849 3585 36917
rect 3509 36793 3519 36849
rect 3575 36793 3585 36849
rect 3509 36725 3585 36793
rect 3509 36669 3519 36725
rect 3575 36669 3585 36725
rect 3509 36601 3585 36669
rect 3509 36545 3519 36601
rect 3575 36545 3585 36601
rect 3509 36535 3585 36545
rect 3633 38089 3709 38099
rect 3633 38033 3643 38089
rect 3699 38033 3709 38089
rect 3633 37965 3709 38033
rect 4460 38036 4536 38104
rect 4460 37980 4470 38036
rect 4526 37980 4536 38036
rect 3633 37909 3643 37965
rect 3699 37909 3709 37965
rect 3633 37841 3709 37909
rect 3633 37785 3643 37841
rect 3699 37785 3709 37841
rect 3633 37717 3709 37785
rect 3633 37661 3643 37717
rect 3699 37661 3709 37717
rect 3633 37593 3709 37661
rect 3633 37537 3643 37593
rect 3699 37537 3709 37593
rect 3633 37469 3709 37537
rect 3633 37413 3643 37469
rect 3699 37413 3709 37469
rect 3633 37345 3709 37413
rect 3633 37289 3643 37345
rect 3699 37289 3709 37345
rect 3633 37221 3709 37289
rect 3633 37165 3643 37221
rect 3699 37165 3709 37221
rect 3633 37097 3709 37165
rect 3633 37041 3643 37097
rect 3699 37041 3709 37097
rect 3633 36973 3709 37041
rect 3633 36917 3643 36973
rect 3699 36917 3709 36973
rect 3633 36849 3709 36917
rect 3633 36793 3643 36849
rect 3699 36793 3709 36849
rect 3633 36725 3709 36793
rect 3633 36669 3643 36725
rect 3699 36669 3709 36725
rect 3633 36601 3709 36669
rect 3633 36545 3643 36601
rect 3699 36545 3709 36601
rect 3633 36477 3709 36545
rect 3633 36421 3643 36477
rect 3699 36421 3709 36477
rect 3633 36411 3709 36421
rect 3757 37965 3833 37975
rect 3757 37909 3767 37965
rect 3823 37909 3833 37965
rect 3757 37841 3833 37909
rect 4460 37912 4536 37980
rect 4460 37856 4470 37912
rect 4526 37856 4536 37912
rect 3757 37785 3767 37841
rect 3823 37785 3833 37841
rect 3757 37717 3833 37785
rect 3757 37661 3767 37717
rect 3823 37661 3833 37717
rect 3757 37593 3833 37661
rect 3757 37537 3767 37593
rect 3823 37537 3833 37593
rect 3757 37469 3833 37537
rect 3757 37413 3767 37469
rect 3823 37413 3833 37469
rect 3757 37345 3833 37413
rect 3757 37289 3767 37345
rect 3823 37289 3833 37345
rect 3757 37221 3833 37289
rect 3757 37165 3767 37221
rect 3823 37165 3833 37221
rect 3757 37097 3833 37165
rect 3757 37041 3767 37097
rect 3823 37041 3833 37097
rect 3757 36973 3833 37041
rect 3757 36917 3767 36973
rect 3823 36917 3833 36973
rect 3757 36849 3833 36917
rect 3757 36793 3767 36849
rect 3823 36793 3833 36849
rect 3757 36725 3833 36793
rect 3757 36669 3767 36725
rect 3823 36669 3833 36725
rect 3757 36601 3833 36669
rect 3757 36545 3767 36601
rect 3823 36545 3833 36601
rect 3757 36477 3833 36545
rect 3757 36421 3767 36477
rect 3823 36421 3833 36477
rect 3757 36353 3833 36421
rect 3757 36297 3767 36353
rect 3823 36297 3833 36353
rect 3757 36287 3833 36297
rect 3881 37841 3957 37851
rect 4460 37846 4536 37856
rect 4584 39400 4660 39410
rect 4584 39344 4594 39400
rect 4650 39344 4660 39400
rect 4584 39276 4660 39344
rect 4584 39220 4594 39276
rect 4650 39220 4660 39276
rect 4584 39152 4660 39220
rect 4584 39096 4594 39152
rect 4650 39096 4660 39152
rect 4584 39028 4660 39096
rect 4584 38972 4594 39028
rect 4650 38972 4660 39028
rect 4584 38904 4660 38972
rect 4584 38848 4594 38904
rect 4650 38848 4660 38904
rect 4584 38780 4660 38848
rect 4584 38724 4594 38780
rect 4650 38724 4660 38780
rect 4584 38656 4660 38724
rect 4584 38600 4594 38656
rect 4650 38600 4660 38656
rect 4584 38532 4660 38600
rect 4584 38476 4594 38532
rect 4650 38476 4660 38532
rect 4584 38408 4660 38476
rect 4584 38352 4594 38408
rect 4650 38352 4660 38408
rect 4584 38284 4660 38352
rect 4584 38228 4594 38284
rect 4650 38228 4660 38284
rect 4584 38160 4660 38228
rect 4584 38104 4594 38160
rect 4650 38104 4660 38160
rect 4584 38036 4660 38104
rect 4584 37980 4594 38036
rect 4650 37980 4660 38036
rect 4584 37912 4660 37980
rect 4584 37856 4594 37912
rect 4650 37856 4660 37912
rect 3881 37785 3891 37841
rect 3947 37785 3957 37841
rect 3881 37717 3957 37785
rect 4584 37788 4660 37856
rect 4584 37732 4594 37788
rect 4650 37732 4660 37788
rect 3881 37661 3891 37717
rect 3947 37661 3957 37717
rect 3881 37593 3957 37661
rect 3881 37537 3891 37593
rect 3947 37537 3957 37593
rect 3881 37469 3957 37537
rect 3881 37413 3891 37469
rect 3947 37413 3957 37469
rect 3881 37345 3957 37413
rect 3881 37289 3891 37345
rect 3947 37289 3957 37345
rect 3881 37221 3957 37289
rect 3881 37165 3891 37221
rect 3947 37165 3957 37221
rect 3881 37097 3957 37165
rect 3881 37041 3891 37097
rect 3947 37041 3957 37097
rect 3881 36973 3957 37041
rect 3881 36917 3891 36973
rect 3947 36917 3957 36973
rect 3881 36849 3957 36917
rect 3881 36793 3891 36849
rect 3947 36793 3957 36849
rect 3881 36725 3957 36793
rect 3881 36669 3891 36725
rect 3947 36669 3957 36725
rect 3881 36601 3957 36669
rect 3881 36545 3891 36601
rect 3947 36545 3957 36601
rect 3881 36477 3957 36545
rect 3881 36421 3891 36477
rect 3947 36421 3957 36477
rect 3881 36353 3957 36421
rect 3881 36297 3891 36353
rect 3947 36297 3957 36353
rect 3881 36229 3957 36297
rect 3881 36173 3891 36229
rect 3947 36173 3957 36229
rect 3881 36163 3957 36173
rect 4005 37717 4081 37727
rect 4584 37722 4660 37732
rect 4708 39276 4784 39286
rect 4708 39220 4718 39276
rect 4774 39220 4784 39276
rect 4708 39152 4784 39220
rect 4708 39096 4718 39152
rect 4774 39096 4784 39152
rect 4708 39028 4784 39096
rect 4708 38972 4718 39028
rect 4774 38972 4784 39028
rect 4708 38904 4784 38972
rect 4708 38848 4718 38904
rect 4774 38848 4784 38904
rect 4708 38780 4784 38848
rect 4708 38724 4718 38780
rect 4774 38724 4784 38780
rect 4708 38656 4784 38724
rect 4708 38600 4718 38656
rect 4774 38600 4784 38656
rect 4708 38532 4784 38600
rect 4708 38476 4718 38532
rect 4774 38476 4784 38532
rect 4708 38408 4784 38476
rect 4708 38352 4718 38408
rect 4774 38352 4784 38408
rect 4708 38284 4784 38352
rect 4708 38228 4718 38284
rect 4774 38228 4784 38284
rect 4708 38160 4784 38228
rect 4708 38104 4718 38160
rect 4774 38104 4784 38160
rect 4708 38036 4784 38104
rect 4708 37980 4718 38036
rect 4774 37980 4784 38036
rect 4708 37912 4784 37980
rect 4708 37856 4718 37912
rect 4774 37856 4784 37912
rect 4708 37788 4784 37856
rect 4708 37732 4718 37788
rect 4774 37732 4784 37788
rect 4005 37661 4015 37717
rect 4071 37661 4081 37717
rect 4005 37593 4081 37661
rect 4708 37664 4784 37732
rect 4708 37608 4718 37664
rect 4774 37608 4784 37664
rect 4005 37537 4015 37593
rect 4071 37537 4081 37593
rect 4005 37469 4081 37537
rect 4005 37413 4015 37469
rect 4071 37413 4081 37469
rect 4005 37345 4081 37413
rect 4005 37289 4015 37345
rect 4071 37289 4081 37345
rect 4005 37221 4081 37289
rect 4005 37165 4015 37221
rect 4071 37165 4081 37221
rect 4005 37097 4081 37165
rect 4005 37041 4015 37097
rect 4071 37041 4081 37097
rect 4005 36973 4081 37041
rect 4005 36917 4015 36973
rect 4071 36917 4081 36973
rect 4005 36849 4081 36917
rect 4005 36793 4015 36849
rect 4071 36793 4081 36849
rect 4005 36725 4081 36793
rect 4005 36669 4015 36725
rect 4071 36669 4081 36725
rect 4005 36601 4081 36669
rect 4005 36545 4015 36601
rect 4071 36545 4081 36601
rect 4005 36477 4081 36545
rect 4005 36421 4015 36477
rect 4071 36421 4081 36477
rect 4005 36353 4081 36421
rect 4005 36297 4015 36353
rect 4071 36297 4081 36353
rect 4005 36229 4081 36297
rect 4005 36173 4015 36229
rect 4071 36173 4081 36229
rect 4005 36105 4081 36173
rect 4005 36049 4015 36105
rect 4071 36049 4081 36105
rect 4005 36039 4081 36049
rect 4129 37593 4205 37603
rect 4708 37598 4784 37608
rect 4832 39152 4908 39162
rect 4832 39096 4842 39152
rect 4898 39096 4908 39152
rect 4832 39028 4908 39096
rect 4832 38972 4842 39028
rect 4898 38972 4908 39028
rect 4832 38904 4908 38972
rect 4832 38848 4842 38904
rect 4898 38848 4908 38904
rect 4832 38780 4908 38848
rect 4832 38724 4842 38780
rect 4898 38724 4908 38780
rect 4832 38656 4908 38724
rect 4832 38600 4842 38656
rect 4898 38600 4908 38656
rect 4832 38532 4908 38600
rect 4832 38476 4842 38532
rect 4898 38476 4908 38532
rect 4832 38408 4908 38476
rect 4832 38352 4842 38408
rect 4898 38352 4908 38408
rect 4832 38284 4908 38352
rect 4832 38228 4842 38284
rect 4898 38228 4908 38284
rect 4832 38160 4908 38228
rect 4832 38104 4842 38160
rect 4898 38104 4908 38160
rect 4832 38036 4908 38104
rect 4832 37980 4842 38036
rect 4898 37980 4908 38036
rect 4832 37912 4908 37980
rect 4832 37856 4842 37912
rect 4898 37856 4908 37912
rect 4832 37788 4908 37856
rect 4832 37732 4842 37788
rect 4898 37732 4908 37788
rect 4832 37664 4908 37732
rect 4832 37608 4842 37664
rect 4898 37608 4908 37664
rect 4129 37537 4139 37593
rect 4195 37537 4205 37593
rect 4129 37469 4205 37537
rect 4832 37540 4908 37608
rect 4832 37484 4842 37540
rect 4898 37484 4908 37540
rect 4832 37474 4908 37484
rect 4956 39028 5032 39038
rect 4956 38972 4966 39028
rect 5022 38972 5032 39028
rect 4956 38904 5032 38972
rect 4956 38848 4966 38904
rect 5022 38848 5032 38904
rect 4956 38780 5032 38848
rect 4956 38724 4966 38780
rect 5022 38724 5032 38780
rect 4956 38656 5032 38724
rect 4956 38600 4966 38656
rect 5022 38600 5032 38656
rect 4956 38532 5032 38600
rect 4956 38476 4966 38532
rect 5022 38476 5032 38532
rect 4956 38408 5032 38476
rect 4956 38352 4966 38408
rect 5022 38352 5032 38408
rect 4956 38284 5032 38352
rect 4956 38228 4966 38284
rect 5022 38228 5032 38284
rect 4956 38160 5032 38228
rect 4956 38104 4966 38160
rect 5022 38104 5032 38160
rect 4956 38036 5032 38104
rect 4956 37980 4966 38036
rect 5022 37980 5032 38036
rect 4956 37912 5032 37980
rect 4956 37856 4966 37912
rect 5022 37856 5032 37912
rect 4956 37788 5032 37856
rect 4956 37732 4966 37788
rect 5022 37732 5032 37788
rect 4956 37664 5032 37732
rect 4956 37608 4966 37664
rect 5022 37608 5032 37664
rect 4956 37540 5032 37608
rect 4956 37484 4966 37540
rect 5022 37484 5032 37540
rect 4129 37413 4139 37469
rect 4195 37413 4205 37469
rect 4129 37345 4205 37413
rect 4956 37416 5032 37484
rect 4956 37360 4966 37416
rect 5022 37360 5032 37416
rect 4956 37350 5032 37360
rect 5080 38904 5156 38914
rect 5080 38848 5090 38904
rect 5146 38848 5156 38904
rect 5080 38780 5156 38848
rect 5080 38724 5090 38780
rect 5146 38724 5156 38780
rect 5080 38656 5156 38724
rect 5080 38600 5090 38656
rect 5146 38600 5156 38656
rect 5080 38532 5156 38600
rect 5080 38476 5090 38532
rect 5146 38476 5156 38532
rect 5080 38408 5156 38476
rect 5080 38352 5090 38408
rect 5146 38352 5156 38408
rect 5080 38284 5156 38352
rect 5080 38228 5090 38284
rect 5146 38228 5156 38284
rect 5080 38160 5156 38228
rect 5080 38104 5090 38160
rect 5146 38104 5156 38160
rect 5080 38036 5156 38104
rect 5080 37980 5090 38036
rect 5146 37980 5156 38036
rect 5080 37912 5156 37980
rect 5080 37856 5090 37912
rect 5146 37856 5156 37912
rect 5080 37788 5156 37856
rect 5080 37732 5090 37788
rect 5146 37732 5156 37788
rect 5080 37664 5156 37732
rect 5080 37608 5090 37664
rect 5146 37608 5156 37664
rect 5080 37540 5156 37608
rect 5080 37484 5090 37540
rect 5146 37484 5156 37540
rect 5080 37416 5156 37484
rect 5080 37360 5090 37416
rect 5146 37360 5156 37416
rect 4129 37289 4139 37345
rect 4195 37289 4205 37345
rect 4129 37221 4205 37289
rect 5080 37292 5156 37360
rect 5080 37236 5090 37292
rect 5146 37236 5156 37292
rect 5080 37226 5156 37236
rect 5204 38780 5280 38790
rect 5204 38724 5214 38780
rect 5270 38724 5280 38780
rect 5204 38656 5280 38724
rect 5204 38600 5214 38656
rect 5270 38600 5280 38656
rect 5204 38532 5280 38600
rect 5204 38476 5214 38532
rect 5270 38476 5280 38532
rect 5204 38408 5280 38476
rect 5204 38352 5214 38408
rect 5270 38352 5280 38408
rect 5204 38284 5280 38352
rect 5204 38228 5214 38284
rect 5270 38228 5280 38284
rect 5204 38160 5280 38228
rect 5204 38104 5214 38160
rect 5270 38104 5280 38160
rect 5204 38036 5280 38104
rect 5204 37980 5214 38036
rect 5270 37980 5280 38036
rect 5204 37912 5280 37980
rect 5204 37856 5214 37912
rect 5270 37856 5280 37912
rect 5204 37788 5280 37856
rect 5204 37732 5214 37788
rect 5270 37732 5280 37788
rect 5204 37664 5280 37732
rect 5204 37608 5214 37664
rect 5270 37608 5280 37664
rect 5204 37540 5280 37608
rect 5204 37484 5214 37540
rect 5270 37484 5280 37540
rect 5204 37416 5280 37484
rect 5204 37360 5214 37416
rect 5270 37360 5280 37416
rect 5204 37292 5280 37360
rect 5204 37236 5214 37292
rect 5270 37236 5280 37292
rect 4129 37165 4139 37221
rect 4195 37165 4205 37221
rect 4129 37097 4205 37165
rect 5204 37168 5280 37236
rect 5204 37112 5214 37168
rect 5270 37112 5280 37168
rect 5204 37102 5280 37112
rect 5328 38656 5404 38666
rect 5328 38600 5338 38656
rect 5394 38600 5404 38656
rect 5328 38532 5404 38600
rect 5328 38476 5338 38532
rect 5394 38476 5404 38532
rect 5328 38408 5404 38476
rect 5328 38352 5338 38408
rect 5394 38352 5404 38408
rect 5328 38284 5404 38352
rect 5328 38228 5338 38284
rect 5394 38228 5404 38284
rect 5328 38160 5404 38228
rect 5328 38104 5338 38160
rect 5394 38104 5404 38160
rect 5328 38036 5404 38104
rect 5328 37980 5338 38036
rect 5394 37980 5404 38036
rect 5328 37912 5404 37980
rect 5328 37856 5338 37912
rect 5394 37856 5404 37912
rect 5328 37788 5404 37856
rect 5328 37732 5338 37788
rect 5394 37732 5404 37788
rect 5328 37664 5404 37732
rect 5328 37608 5338 37664
rect 5394 37608 5404 37664
rect 5328 37540 5404 37608
rect 5328 37484 5338 37540
rect 5394 37484 5404 37540
rect 5328 37416 5404 37484
rect 5328 37360 5338 37416
rect 5394 37360 5404 37416
rect 5328 37292 5404 37360
rect 5328 37236 5338 37292
rect 5394 37236 5404 37292
rect 5328 37168 5404 37236
rect 5328 37112 5338 37168
rect 5394 37112 5404 37168
rect 4129 37041 4139 37097
rect 4195 37041 4205 37097
rect 4129 36973 4205 37041
rect 5328 37044 5404 37112
rect 5328 36988 5338 37044
rect 5394 36988 5404 37044
rect 5328 36978 5404 36988
rect 5452 38532 5528 38542
rect 5452 38476 5462 38532
rect 5518 38476 5528 38532
rect 5452 38408 5528 38476
rect 5452 38352 5462 38408
rect 5518 38352 5528 38408
rect 5452 38284 5528 38352
rect 5452 38228 5462 38284
rect 5518 38228 5528 38284
rect 5452 38160 5528 38228
rect 5452 38104 5462 38160
rect 5518 38104 5528 38160
rect 5452 38036 5528 38104
rect 5452 37980 5462 38036
rect 5518 37980 5528 38036
rect 5452 37912 5528 37980
rect 5452 37856 5462 37912
rect 5518 37856 5528 37912
rect 5452 37788 5528 37856
rect 5452 37732 5462 37788
rect 5518 37732 5528 37788
rect 5452 37664 5528 37732
rect 5452 37608 5462 37664
rect 5518 37608 5528 37664
rect 5452 37540 5528 37608
rect 5452 37484 5462 37540
rect 5518 37484 5528 37540
rect 5452 37416 5528 37484
rect 5452 37360 5462 37416
rect 5518 37360 5528 37416
rect 5452 37292 5528 37360
rect 5452 37236 5462 37292
rect 5518 37236 5528 37292
rect 5452 37168 5528 37236
rect 5452 37112 5462 37168
rect 5518 37112 5528 37168
rect 5452 37044 5528 37112
rect 5452 36988 5462 37044
rect 5518 36988 5528 37044
rect 4129 36917 4139 36973
rect 4195 36917 4205 36973
rect 4129 36849 4205 36917
rect 5452 36920 5528 36988
rect 5452 36864 5462 36920
rect 5518 36864 5528 36920
rect 5452 36854 5528 36864
rect 5576 38402 5652 38412
rect 5576 38346 5586 38402
rect 5642 38346 5652 38402
rect 5576 38278 5652 38346
rect 5576 38222 5586 38278
rect 5642 38222 5652 38278
rect 5576 38154 5652 38222
rect 5576 38098 5586 38154
rect 5642 38098 5652 38154
rect 5576 38030 5652 38098
rect 5576 37974 5586 38030
rect 5642 37974 5652 38030
rect 5576 37906 5652 37974
rect 5576 37850 5586 37906
rect 5642 37850 5652 37906
rect 5576 37782 5652 37850
rect 5576 37726 5586 37782
rect 5642 37726 5652 37782
rect 5576 37658 5652 37726
rect 5576 37602 5586 37658
rect 5642 37602 5652 37658
rect 5576 37534 5652 37602
rect 5576 37478 5586 37534
rect 5642 37478 5652 37534
rect 5576 37410 5652 37478
rect 5576 37354 5586 37410
rect 5642 37354 5652 37410
rect 5576 37286 5652 37354
rect 5576 37230 5586 37286
rect 5642 37230 5652 37286
rect 5576 37162 5652 37230
rect 5576 37106 5586 37162
rect 5642 37106 5652 37162
rect 5576 37038 5652 37106
rect 5576 36982 5586 37038
rect 5642 36982 5652 37038
rect 5576 36914 5652 36982
rect 5576 36858 5586 36914
rect 5642 36858 5652 36914
rect 4129 36793 4139 36849
rect 4195 36793 4205 36849
rect 5576 36848 5652 36858
rect 5700 38273 5776 38283
rect 5700 38217 5710 38273
rect 5766 38217 5776 38273
rect 5700 38149 5776 38217
rect 5700 38093 5710 38149
rect 5766 38093 5776 38149
rect 5700 38025 5776 38093
rect 5700 37969 5710 38025
rect 5766 37969 5776 38025
rect 5700 37901 5776 37969
rect 5700 37845 5710 37901
rect 5766 37845 5776 37901
rect 5700 37777 5776 37845
rect 5700 37721 5710 37777
rect 5766 37721 5776 37777
rect 5700 37653 5776 37721
rect 5700 37597 5710 37653
rect 5766 37597 5776 37653
rect 5700 37529 5776 37597
rect 5700 37473 5710 37529
rect 5766 37473 5776 37529
rect 5700 37405 5776 37473
rect 5700 37349 5710 37405
rect 5766 37349 5776 37405
rect 5700 37281 5776 37349
rect 5700 37225 5710 37281
rect 5766 37225 5776 37281
rect 5700 37157 5776 37225
rect 5700 37101 5710 37157
rect 5766 37101 5776 37157
rect 5700 37033 5776 37101
rect 5700 36977 5710 37033
rect 5766 36977 5776 37033
rect 5700 36909 5776 36977
rect 5700 36853 5710 36909
rect 5766 36853 5776 36909
rect 5824 38162 5900 38172
rect 5824 38106 5834 38162
rect 5890 38106 5900 38162
rect 5824 38038 5900 38106
rect 5824 37982 5834 38038
rect 5890 37982 5900 38038
rect 5824 37914 5900 37982
rect 5824 37858 5834 37914
rect 5890 37858 5900 37914
rect 5824 37790 5900 37858
rect 5824 37734 5834 37790
rect 5890 37734 5900 37790
rect 5824 37666 5900 37734
rect 5824 37610 5834 37666
rect 5890 37610 5900 37666
rect 5824 37542 5900 37610
rect 5824 37486 5834 37542
rect 5890 37486 5900 37542
rect 5824 37418 5900 37486
rect 5824 37362 5834 37418
rect 5890 37362 5900 37418
rect 5824 37294 5900 37362
rect 5824 37238 5834 37294
rect 5890 37238 5900 37294
rect 5824 37170 5900 37238
rect 5824 37114 5834 37170
rect 5890 37114 5900 37170
rect 5824 37046 5900 37114
rect 5824 36990 5834 37046
rect 5890 36990 5900 37046
rect 5824 36922 5900 36990
rect 5824 36866 5834 36922
rect 5890 36866 5900 36922
rect 5824 36856 5900 36866
rect 5948 38141 6024 38151
rect 5948 38085 5958 38141
rect 6014 38085 6024 38141
rect 5948 38017 6024 38085
rect 5948 37961 5958 38017
rect 6014 37961 6024 38017
rect 5948 37893 6024 37961
rect 5948 37837 5958 37893
rect 6014 37837 6024 37893
rect 5948 37769 6024 37837
rect 5948 37713 5958 37769
rect 6014 37713 6024 37769
rect 5948 37645 6024 37713
rect 5948 37589 5958 37645
rect 6014 37589 6024 37645
rect 5948 37521 6024 37589
rect 5948 37465 5958 37521
rect 6014 37465 6024 37521
rect 5948 37397 6024 37465
rect 5948 37341 5958 37397
rect 6014 37341 6024 37397
rect 5948 37273 6024 37341
rect 5948 37217 5958 37273
rect 6014 37217 6024 37273
rect 5948 37149 6024 37217
rect 5948 37093 5958 37149
rect 6014 37093 6024 37149
rect 5948 37025 6024 37093
rect 5948 36969 5958 37025
rect 6014 36969 6024 37025
rect 5948 36901 6024 36969
rect 5700 36843 5776 36853
rect 5948 36845 5958 36901
rect 6014 36845 6024 36901
rect 5948 36835 6024 36845
rect 6072 38140 6148 38150
rect 6072 38084 6082 38140
rect 6138 38084 6148 38140
rect 6072 38016 6148 38084
rect 6072 37960 6082 38016
rect 6138 37960 6148 38016
rect 6072 37892 6148 37960
rect 6072 37836 6082 37892
rect 6138 37836 6148 37892
rect 6072 37768 6148 37836
rect 6072 37712 6082 37768
rect 6138 37712 6148 37768
rect 6072 37644 6148 37712
rect 6072 37588 6082 37644
rect 6138 37588 6148 37644
rect 6072 37520 6148 37588
rect 6072 37464 6082 37520
rect 6138 37464 6148 37520
rect 6072 37396 6148 37464
rect 6072 37340 6082 37396
rect 6138 37340 6148 37396
rect 6072 37272 6148 37340
rect 6072 37216 6082 37272
rect 6138 37216 6148 37272
rect 6072 37148 6148 37216
rect 6072 37092 6082 37148
rect 6138 37092 6148 37148
rect 6072 37024 6148 37092
rect 6072 36968 6082 37024
rect 6138 36968 6148 37024
rect 6072 36900 6148 36968
rect 6072 36844 6082 36900
rect 6138 36844 6148 36900
rect 6072 36834 6148 36844
rect 7552 38144 8620 38154
rect 7552 38088 7562 38144
rect 7618 38088 7686 38144
rect 7742 38088 7810 38144
rect 7866 38088 7934 38144
rect 7990 38088 8058 38144
rect 8114 38088 8182 38144
rect 8238 38088 8306 38144
rect 8362 38088 8430 38144
rect 8486 38088 8554 38144
rect 8610 38088 8620 38144
rect 7552 38020 8620 38088
rect 7552 37964 7562 38020
rect 7618 37964 7686 38020
rect 7742 37964 7810 38020
rect 7866 37964 7934 38020
rect 7990 37964 8058 38020
rect 8114 37964 8182 38020
rect 8238 37964 8306 38020
rect 8362 37964 8430 38020
rect 8486 37964 8554 38020
rect 8610 37964 8620 38020
rect 7552 37896 8620 37964
rect 7552 37840 7562 37896
rect 7618 37840 7686 37896
rect 7742 37840 7810 37896
rect 7866 37840 7934 37896
rect 7990 37840 8058 37896
rect 8114 37840 8182 37896
rect 8238 37840 8306 37896
rect 8362 37840 8430 37896
rect 8486 37840 8554 37896
rect 8610 37840 8620 37896
rect 7552 37772 8620 37840
rect 7552 37716 7562 37772
rect 7618 37716 7686 37772
rect 7742 37716 7810 37772
rect 7866 37716 7934 37772
rect 7990 37716 8058 37772
rect 8114 37716 8182 37772
rect 8238 37716 8306 37772
rect 8362 37716 8430 37772
rect 8486 37716 8554 37772
rect 8610 37716 8620 37772
rect 7552 37648 8620 37716
rect 7552 37592 7562 37648
rect 7618 37592 7686 37648
rect 7742 37592 7810 37648
rect 7866 37592 7934 37648
rect 7990 37592 8058 37648
rect 8114 37592 8182 37648
rect 8238 37592 8306 37648
rect 8362 37592 8430 37648
rect 8486 37592 8554 37648
rect 8610 37592 8620 37648
rect 7552 37524 8620 37592
rect 7552 37468 7562 37524
rect 7618 37468 7686 37524
rect 7742 37468 7810 37524
rect 7866 37468 7934 37524
rect 7990 37468 8058 37524
rect 8114 37468 8182 37524
rect 8238 37468 8306 37524
rect 8362 37468 8430 37524
rect 8486 37468 8554 37524
rect 8610 37468 8620 37524
rect 7552 37400 8620 37468
rect 7552 37344 7562 37400
rect 7618 37344 7686 37400
rect 7742 37344 7810 37400
rect 7866 37344 7934 37400
rect 7990 37344 8058 37400
rect 8114 37344 8182 37400
rect 8238 37344 8306 37400
rect 8362 37344 8430 37400
rect 8486 37344 8554 37400
rect 8610 37344 8620 37400
rect 7552 37276 8620 37344
rect 7552 37220 7562 37276
rect 7618 37220 7686 37276
rect 7742 37220 7810 37276
rect 7866 37220 7934 37276
rect 7990 37220 8058 37276
rect 8114 37220 8182 37276
rect 8238 37220 8306 37276
rect 8362 37220 8430 37276
rect 8486 37220 8554 37276
rect 8610 37220 8620 37276
rect 7552 37152 8620 37220
rect 7552 37096 7562 37152
rect 7618 37096 7686 37152
rect 7742 37096 7810 37152
rect 7866 37096 7934 37152
rect 7990 37096 8058 37152
rect 8114 37096 8182 37152
rect 8238 37096 8306 37152
rect 8362 37096 8430 37152
rect 8486 37096 8554 37152
rect 8610 37096 8620 37152
rect 7552 37028 8620 37096
rect 7552 36972 7562 37028
rect 7618 36972 7686 37028
rect 7742 36972 7810 37028
rect 7866 36972 7934 37028
rect 7990 36972 8058 37028
rect 8114 36972 8182 37028
rect 8238 36972 8306 37028
rect 8362 36972 8430 37028
rect 8486 36972 8554 37028
rect 8610 36972 8620 37028
rect 7552 36904 8620 36972
rect 7552 36848 7562 36904
rect 7618 36848 7686 36904
rect 7742 36848 7810 36904
rect 7866 36848 7934 36904
rect 7990 36848 8058 36904
rect 8114 36848 8182 36904
rect 8238 36848 8306 36904
rect 8362 36848 8430 36904
rect 8486 36848 8554 36904
rect 8610 36848 8620 36904
rect 7552 36838 8620 36848
rect 10669 38144 12481 38154
rect 10669 38088 10679 38144
rect 10735 38088 10803 38144
rect 10859 38088 10927 38144
rect 10983 38088 11051 38144
rect 11107 38088 11175 38144
rect 11231 38088 11299 38144
rect 11355 38088 11423 38144
rect 11479 38088 11547 38144
rect 11603 38088 11671 38144
rect 11727 38088 11795 38144
rect 11851 38088 11919 38144
rect 11975 38088 12043 38144
rect 12099 38088 12167 38144
rect 12223 38088 12291 38144
rect 12347 38088 12415 38144
rect 12471 38088 12481 38144
rect 10669 38020 12481 38088
rect 10669 37964 10679 38020
rect 10735 37964 10803 38020
rect 10859 37964 10927 38020
rect 10983 37964 11051 38020
rect 11107 37964 11175 38020
rect 11231 37964 11299 38020
rect 11355 37964 11423 38020
rect 11479 37964 11547 38020
rect 11603 37964 11671 38020
rect 11727 37964 11795 38020
rect 11851 37964 11919 38020
rect 11975 37964 12043 38020
rect 12099 37964 12167 38020
rect 12223 37964 12291 38020
rect 12347 37964 12415 38020
rect 12471 37964 12481 38020
rect 10669 37896 12481 37964
rect 10669 37840 10679 37896
rect 10735 37840 10803 37896
rect 10859 37840 10927 37896
rect 10983 37840 11051 37896
rect 11107 37840 11175 37896
rect 11231 37840 11299 37896
rect 11355 37840 11423 37896
rect 11479 37840 11547 37896
rect 11603 37840 11671 37896
rect 11727 37840 11795 37896
rect 11851 37840 11919 37896
rect 11975 37840 12043 37896
rect 12099 37840 12167 37896
rect 12223 37840 12291 37896
rect 12347 37840 12415 37896
rect 12471 37840 12481 37896
rect 10669 37772 12481 37840
rect 10669 37716 10679 37772
rect 10735 37716 10803 37772
rect 10859 37716 10927 37772
rect 10983 37716 11051 37772
rect 11107 37716 11175 37772
rect 11231 37716 11299 37772
rect 11355 37716 11423 37772
rect 11479 37716 11547 37772
rect 11603 37716 11671 37772
rect 11727 37716 11795 37772
rect 11851 37716 11919 37772
rect 11975 37716 12043 37772
rect 12099 37716 12167 37772
rect 12223 37716 12291 37772
rect 12347 37716 12415 37772
rect 12471 37716 12481 37772
rect 10669 37648 12481 37716
rect 10669 37592 10679 37648
rect 10735 37592 10803 37648
rect 10859 37592 10927 37648
rect 10983 37592 11051 37648
rect 11107 37592 11175 37648
rect 11231 37592 11299 37648
rect 11355 37592 11423 37648
rect 11479 37592 11547 37648
rect 11603 37592 11671 37648
rect 11727 37592 11795 37648
rect 11851 37592 11919 37648
rect 11975 37592 12043 37648
rect 12099 37592 12167 37648
rect 12223 37592 12291 37648
rect 12347 37592 12415 37648
rect 12471 37592 12481 37648
rect 10669 37524 12481 37592
rect 10669 37468 10679 37524
rect 10735 37468 10803 37524
rect 10859 37468 10927 37524
rect 10983 37468 11051 37524
rect 11107 37468 11175 37524
rect 11231 37468 11299 37524
rect 11355 37468 11423 37524
rect 11479 37468 11547 37524
rect 11603 37468 11671 37524
rect 11727 37468 11795 37524
rect 11851 37468 11919 37524
rect 11975 37468 12043 37524
rect 12099 37468 12167 37524
rect 12223 37468 12291 37524
rect 12347 37468 12415 37524
rect 12471 37468 12481 37524
rect 10669 37400 12481 37468
rect 10669 37344 10679 37400
rect 10735 37344 10803 37400
rect 10859 37344 10927 37400
rect 10983 37344 11051 37400
rect 11107 37344 11175 37400
rect 11231 37344 11299 37400
rect 11355 37344 11423 37400
rect 11479 37344 11547 37400
rect 11603 37344 11671 37400
rect 11727 37344 11795 37400
rect 11851 37344 11919 37400
rect 11975 37344 12043 37400
rect 12099 37344 12167 37400
rect 12223 37344 12291 37400
rect 12347 37344 12415 37400
rect 12471 37344 12481 37400
rect 10669 37276 12481 37344
rect 10669 37220 10679 37276
rect 10735 37220 10803 37276
rect 10859 37220 10927 37276
rect 10983 37220 11051 37276
rect 11107 37220 11175 37276
rect 11231 37220 11299 37276
rect 11355 37220 11423 37276
rect 11479 37220 11547 37276
rect 11603 37220 11671 37276
rect 11727 37220 11795 37276
rect 11851 37220 11919 37276
rect 11975 37220 12043 37276
rect 12099 37220 12167 37276
rect 12223 37220 12291 37276
rect 12347 37220 12415 37276
rect 12471 37220 12481 37276
rect 10669 37152 12481 37220
rect 10669 37096 10679 37152
rect 10735 37096 10803 37152
rect 10859 37096 10927 37152
rect 10983 37096 11051 37152
rect 11107 37096 11175 37152
rect 11231 37096 11299 37152
rect 11355 37096 11423 37152
rect 11479 37096 11547 37152
rect 11603 37096 11671 37152
rect 11727 37096 11795 37152
rect 11851 37096 11919 37152
rect 11975 37096 12043 37152
rect 12099 37096 12167 37152
rect 12223 37096 12291 37152
rect 12347 37096 12415 37152
rect 12471 37096 12481 37152
rect 10669 37028 12481 37096
rect 10669 36972 10679 37028
rect 10735 36972 10803 37028
rect 10859 36972 10927 37028
rect 10983 36972 11051 37028
rect 11107 36972 11175 37028
rect 11231 36972 11299 37028
rect 11355 36972 11423 37028
rect 11479 36972 11547 37028
rect 11603 36972 11671 37028
rect 11727 36972 11795 37028
rect 11851 36972 11919 37028
rect 11975 36972 12043 37028
rect 12099 36972 12167 37028
rect 12223 36972 12291 37028
rect 12347 36972 12415 37028
rect 12471 36972 12481 37028
rect 10669 36904 12481 36972
rect 10669 36848 10679 36904
rect 10735 36848 10803 36904
rect 10859 36848 10927 36904
rect 10983 36848 11051 36904
rect 11107 36848 11175 36904
rect 11231 36848 11299 36904
rect 11355 36848 11423 36904
rect 11479 36848 11547 36904
rect 11603 36848 11671 36904
rect 11727 36848 11795 36904
rect 11851 36848 11919 36904
rect 11975 36848 12043 36904
rect 12099 36848 12167 36904
rect 12223 36848 12291 36904
rect 12347 36848 12415 36904
rect 12471 36848 12481 36904
rect 10669 36838 12481 36848
rect 4129 36725 4205 36793
rect 4129 36669 4139 36725
rect 4195 36669 4205 36725
rect 4129 36601 4205 36669
rect 4129 36545 4139 36601
rect 4195 36545 4205 36601
rect 14757 36572 14833 36582
rect 4129 36477 4205 36545
rect 4129 36421 4139 36477
rect 4195 36421 4205 36477
rect 4129 36353 4205 36421
rect 4129 36297 4139 36353
rect 4195 36297 4205 36353
rect 4129 36229 4205 36297
rect 4129 36173 4139 36229
rect 4195 36173 4205 36229
rect 4129 36105 4205 36173
rect 4129 36049 4139 36105
rect 4195 36049 4205 36105
rect 4129 35981 4205 36049
rect 4129 35925 4139 35981
rect 4195 35925 4205 35981
rect 4129 35915 4205 35925
rect 6358 36544 7426 36554
rect 6358 36488 6368 36544
rect 6424 36488 6492 36544
rect 6548 36488 6616 36544
rect 6672 36488 6740 36544
rect 6796 36488 6864 36544
rect 6920 36488 6988 36544
rect 7044 36488 7112 36544
rect 7168 36488 7236 36544
rect 7292 36488 7360 36544
rect 7416 36488 7426 36544
rect 6358 36420 7426 36488
rect 6358 36364 6368 36420
rect 6424 36364 6492 36420
rect 6548 36364 6616 36420
rect 6672 36364 6740 36420
rect 6796 36364 6864 36420
rect 6920 36364 6988 36420
rect 7044 36364 7112 36420
rect 7168 36364 7236 36420
rect 7292 36364 7360 36420
rect 7416 36364 7426 36420
rect 6358 36296 7426 36364
rect 6358 36240 6368 36296
rect 6424 36240 6492 36296
rect 6548 36240 6616 36296
rect 6672 36240 6740 36296
rect 6796 36240 6864 36296
rect 6920 36240 6988 36296
rect 7044 36240 7112 36296
rect 7168 36240 7236 36296
rect 7292 36240 7360 36296
rect 7416 36240 7426 36296
rect 6358 36172 7426 36240
rect 6358 36116 6368 36172
rect 6424 36116 6492 36172
rect 6548 36116 6616 36172
rect 6672 36116 6740 36172
rect 6796 36116 6864 36172
rect 6920 36116 6988 36172
rect 7044 36116 7112 36172
rect 7168 36116 7236 36172
rect 7292 36116 7360 36172
rect 7416 36116 7426 36172
rect 6358 36048 7426 36116
rect 6358 35992 6368 36048
rect 6424 35992 6492 36048
rect 6548 35992 6616 36048
rect 6672 35992 6740 36048
rect 6796 35992 6864 36048
rect 6920 35992 6988 36048
rect 7044 35992 7112 36048
rect 7168 35992 7236 36048
rect 7292 35992 7360 36048
rect 7416 35992 7426 36048
rect 6358 35924 7426 35992
rect 6358 35868 6368 35924
rect 6424 35868 6492 35924
rect 6548 35868 6616 35924
rect 6672 35868 6740 35924
rect 6796 35868 6864 35924
rect 6920 35868 6988 35924
rect 7044 35868 7112 35924
rect 7168 35868 7236 35924
rect 7292 35868 7360 35924
rect 7416 35868 7426 35924
rect 6358 35800 7426 35868
rect 6358 35744 6368 35800
rect 6424 35744 6492 35800
rect 6548 35744 6616 35800
rect 6672 35744 6740 35800
rect 6796 35744 6864 35800
rect 6920 35744 6988 35800
rect 7044 35744 7112 35800
rect 7168 35744 7236 35800
rect 7292 35744 7360 35800
rect 7416 35744 7426 35800
rect 6358 35676 7426 35744
rect 6358 35620 6368 35676
rect 6424 35620 6492 35676
rect 6548 35620 6616 35676
rect 6672 35620 6740 35676
rect 6796 35620 6864 35676
rect 6920 35620 6988 35676
rect 7044 35620 7112 35676
rect 7168 35620 7236 35676
rect 7292 35620 7360 35676
rect 7416 35620 7426 35676
rect 6358 35552 7426 35620
rect 6358 35496 6368 35552
rect 6424 35496 6492 35552
rect 6548 35496 6616 35552
rect 6672 35496 6740 35552
rect 6796 35496 6864 35552
rect 6920 35496 6988 35552
rect 7044 35496 7112 35552
rect 7168 35496 7236 35552
rect 7292 35496 7360 35552
rect 7416 35496 7426 35552
rect 6358 35428 7426 35496
rect 6358 35372 6368 35428
rect 6424 35372 6492 35428
rect 6548 35372 6616 35428
rect 6672 35372 6740 35428
rect 6796 35372 6864 35428
rect 6920 35372 6988 35428
rect 7044 35372 7112 35428
rect 7168 35372 7236 35428
rect 7292 35372 7360 35428
rect 7416 35372 7426 35428
rect 6358 35304 7426 35372
rect 6358 35248 6368 35304
rect 6424 35248 6492 35304
rect 6548 35248 6616 35304
rect 6672 35248 6740 35304
rect 6796 35248 6864 35304
rect 6920 35248 6988 35304
rect 7044 35248 7112 35304
rect 7168 35248 7236 35304
rect 7292 35248 7360 35304
rect 7416 35248 7426 35304
rect 6358 35238 7426 35248
rect 8741 36544 10553 36554
rect 8741 36488 8751 36544
rect 8807 36488 8875 36544
rect 8931 36488 8999 36544
rect 9055 36488 9123 36544
rect 9179 36488 9247 36544
rect 9303 36488 9371 36544
rect 9427 36488 9495 36544
rect 9551 36488 9619 36544
rect 9675 36488 9743 36544
rect 9799 36488 9867 36544
rect 9923 36488 9991 36544
rect 10047 36488 10115 36544
rect 10171 36488 10239 36544
rect 10295 36488 10363 36544
rect 10419 36488 10487 36544
rect 10543 36488 10553 36544
rect 8741 36420 10553 36488
rect 8741 36364 8751 36420
rect 8807 36364 8875 36420
rect 8931 36364 8999 36420
rect 9055 36364 9123 36420
rect 9179 36364 9247 36420
rect 9303 36364 9371 36420
rect 9427 36364 9495 36420
rect 9551 36364 9619 36420
rect 9675 36364 9743 36420
rect 9799 36364 9867 36420
rect 9923 36364 9991 36420
rect 10047 36364 10115 36420
rect 10171 36364 10239 36420
rect 10295 36364 10363 36420
rect 10419 36364 10487 36420
rect 10543 36364 10553 36420
rect 8741 36296 10553 36364
rect 8741 36240 8751 36296
rect 8807 36240 8875 36296
rect 8931 36240 8999 36296
rect 9055 36240 9123 36296
rect 9179 36240 9247 36296
rect 9303 36240 9371 36296
rect 9427 36240 9495 36296
rect 9551 36240 9619 36296
rect 9675 36240 9743 36296
rect 9799 36240 9867 36296
rect 9923 36240 9991 36296
rect 10047 36240 10115 36296
rect 10171 36240 10239 36296
rect 10295 36240 10363 36296
rect 10419 36240 10487 36296
rect 10543 36240 10553 36296
rect 8741 36172 10553 36240
rect 8741 36116 8751 36172
rect 8807 36116 8875 36172
rect 8931 36116 8999 36172
rect 9055 36116 9123 36172
rect 9179 36116 9247 36172
rect 9303 36116 9371 36172
rect 9427 36116 9495 36172
rect 9551 36116 9619 36172
rect 9675 36116 9743 36172
rect 9799 36116 9867 36172
rect 9923 36116 9991 36172
rect 10047 36116 10115 36172
rect 10171 36116 10239 36172
rect 10295 36116 10363 36172
rect 10419 36116 10487 36172
rect 10543 36116 10553 36172
rect 8741 36048 10553 36116
rect 8741 35992 8751 36048
rect 8807 35992 8875 36048
rect 8931 35992 8999 36048
rect 9055 35992 9123 36048
rect 9179 35992 9247 36048
rect 9303 35992 9371 36048
rect 9427 35992 9495 36048
rect 9551 35992 9619 36048
rect 9675 35992 9743 36048
rect 9799 35992 9867 36048
rect 9923 35992 9991 36048
rect 10047 35992 10115 36048
rect 10171 35992 10239 36048
rect 10295 35992 10363 36048
rect 10419 35992 10487 36048
rect 10543 35992 10553 36048
rect 8741 35924 10553 35992
rect 8741 35868 8751 35924
rect 8807 35868 8875 35924
rect 8931 35868 8999 35924
rect 9055 35868 9123 35924
rect 9179 35868 9247 35924
rect 9303 35868 9371 35924
rect 9427 35868 9495 35924
rect 9551 35868 9619 35924
rect 9675 35868 9743 35924
rect 9799 35868 9867 35924
rect 9923 35868 9991 35924
rect 10047 35868 10115 35924
rect 10171 35868 10239 35924
rect 10295 35868 10363 35924
rect 10419 35868 10487 35924
rect 10543 35868 10553 35924
rect 8741 35800 10553 35868
rect 8741 35744 8751 35800
rect 8807 35744 8875 35800
rect 8931 35744 8999 35800
rect 9055 35744 9123 35800
rect 9179 35744 9247 35800
rect 9303 35744 9371 35800
rect 9427 35744 9495 35800
rect 9551 35744 9619 35800
rect 9675 35744 9743 35800
rect 9799 35744 9867 35800
rect 9923 35744 9991 35800
rect 10047 35744 10115 35800
rect 10171 35744 10239 35800
rect 10295 35744 10363 35800
rect 10419 35744 10487 35800
rect 10543 35744 10553 35800
rect 8741 35676 10553 35744
rect 8741 35620 8751 35676
rect 8807 35620 8875 35676
rect 8931 35620 8999 35676
rect 9055 35620 9123 35676
rect 9179 35620 9247 35676
rect 9303 35620 9371 35676
rect 9427 35620 9495 35676
rect 9551 35620 9619 35676
rect 9675 35620 9743 35676
rect 9799 35620 9867 35676
rect 9923 35620 9991 35676
rect 10047 35620 10115 35676
rect 10171 35620 10239 35676
rect 10295 35620 10363 35676
rect 10419 35620 10487 35676
rect 10543 35620 10553 35676
rect 8741 35552 10553 35620
rect 8741 35496 8751 35552
rect 8807 35496 8875 35552
rect 8931 35496 8999 35552
rect 9055 35496 9123 35552
rect 9179 35496 9247 35552
rect 9303 35496 9371 35552
rect 9427 35496 9495 35552
rect 9551 35496 9619 35552
rect 9675 35496 9743 35552
rect 9799 35496 9867 35552
rect 9923 35496 9991 35552
rect 10047 35496 10115 35552
rect 10171 35496 10239 35552
rect 10295 35496 10363 35552
rect 10419 35496 10487 35552
rect 10543 35496 10553 35552
rect 8741 35428 10553 35496
rect 8741 35372 8751 35428
rect 8807 35372 8875 35428
rect 8931 35372 8999 35428
rect 9055 35372 9123 35428
rect 9179 35372 9247 35428
rect 9303 35372 9371 35428
rect 9427 35372 9495 35428
rect 9551 35372 9619 35428
rect 9675 35372 9743 35428
rect 9799 35372 9867 35428
rect 9923 35372 9991 35428
rect 10047 35372 10115 35428
rect 10171 35372 10239 35428
rect 10295 35372 10363 35428
rect 10419 35372 10487 35428
rect 10543 35372 10553 35428
rect 8741 35304 10553 35372
rect 8741 35248 8751 35304
rect 8807 35248 8875 35304
rect 8931 35248 8999 35304
rect 9055 35248 9123 35304
rect 9179 35248 9247 35304
rect 9303 35248 9371 35304
rect 9427 35248 9495 35304
rect 9551 35248 9619 35304
rect 9675 35248 9743 35304
rect 9799 35248 9867 35304
rect 9923 35248 9991 35304
rect 10047 35248 10115 35304
rect 10171 35248 10239 35304
rect 10295 35248 10363 35304
rect 10419 35248 10487 35304
rect 10543 35248 10553 35304
rect 8741 35238 10553 35248
rect 12842 36544 13910 36554
rect 12842 36488 12852 36544
rect 12908 36488 12976 36544
rect 13032 36488 13100 36544
rect 13156 36488 13224 36544
rect 13280 36488 13348 36544
rect 13404 36488 13472 36544
rect 13528 36488 13596 36544
rect 13652 36488 13720 36544
rect 13776 36488 13844 36544
rect 13900 36488 13910 36544
rect 12842 36420 13910 36488
rect 12842 36364 12852 36420
rect 12908 36364 12976 36420
rect 13032 36364 13100 36420
rect 13156 36364 13224 36420
rect 13280 36364 13348 36420
rect 13404 36364 13472 36420
rect 13528 36364 13596 36420
rect 13652 36364 13720 36420
rect 13776 36364 13844 36420
rect 13900 36364 13910 36420
rect 12842 36296 13910 36364
rect 12842 36240 12852 36296
rect 12908 36240 12976 36296
rect 13032 36240 13100 36296
rect 13156 36240 13224 36296
rect 13280 36240 13348 36296
rect 13404 36240 13472 36296
rect 13528 36240 13596 36296
rect 13652 36240 13720 36296
rect 13776 36240 13844 36296
rect 13900 36240 13910 36296
rect 12842 36172 13910 36240
rect 12842 36116 12852 36172
rect 12908 36116 12976 36172
rect 13032 36116 13100 36172
rect 13156 36116 13224 36172
rect 13280 36116 13348 36172
rect 13404 36116 13472 36172
rect 13528 36116 13596 36172
rect 13652 36116 13720 36172
rect 13776 36116 13844 36172
rect 13900 36116 13910 36172
rect 12842 36048 13910 36116
rect 12842 35992 12852 36048
rect 12908 35992 12976 36048
rect 13032 35992 13100 36048
rect 13156 35992 13224 36048
rect 13280 35992 13348 36048
rect 13404 35992 13472 36048
rect 13528 35992 13596 36048
rect 13652 35992 13720 36048
rect 13776 35992 13844 36048
rect 13900 35992 13910 36048
rect 12842 35924 13910 35992
rect 12842 35868 12852 35924
rect 12908 35868 12976 35924
rect 13032 35868 13100 35924
rect 13156 35868 13224 35924
rect 13280 35868 13348 35924
rect 13404 35868 13472 35924
rect 13528 35868 13596 35924
rect 13652 35868 13720 35924
rect 13776 35868 13844 35924
rect 13900 35868 13910 35924
rect 12842 35800 13910 35868
rect 12842 35744 12852 35800
rect 12908 35744 12976 35800
rect 13032 35744 13100 35800
rect 13156 35744 13224 35800
rect 13280 35744 13348 35800
rect 13404 35744 13472 35800
rect 13528 35744 13596 35800
rect 13652 35744 13720 35800
rect 13776 35744 13844 35800
rect 13900 35744 13910 35800
rect 12842 35676 13910 35744
rect 12842 35620 12852 35676
rect 12908 35620 12976 35676
rect 13032 35620 13100 35676
rect 13156 35620 13224 35676
rect 13280 35620 13348 35676
rect 13404 35620 13472 35676
rect 13528 35620 13596 35676
rect 13652 35620 13720 35676
rect 13776 35620 13844 35676
rect 13900 35620 13910 35676
rect 12842 35552 13910 35620
rect 12842 35496 12852 35552
rect 12908 35496 12976 35552
rect 13032 35496 13100 35552
rect 13156 35496 13224 35552
rect 13280 35496 13348 35552
rect 13404 35496 13472 35552
rect 13528 35496 13596 35552
rect 13652 35496 13720 35552
rect 13776 35496 13844 35552
rect 13900 35496 13910 35552
rect 12842 35428 13910 35496
rect 12842 35372 12852 35428
rect 12908 35372 12976 35428
rect 13032 35372 13100 35428
rect 13156 35372 13224 35428
rect 13280 35372 13348 35428
rect 13404 35372 13472 35428
rect 13528 35372 13596 35428
rect 13652 35372 13720 35428
rect 13776 35372 13844 35428
rect 13900 35372 13910 35428
rect 12842 35304 13910 35372
rect 12842 35248 12852 35304
rect 12908 35248 12976 35304
rect 13032 35248 13100 35304
rect 13156 35248 13224 35304
rect 13280 35248 13348 35304
rect 13404 35248 13472 35304
rect 13528 35248 13596 35304
rect 13652 35248 13720 35304
rect 13776 35248 13844 35304
rect 13900 35248 13910 35304
rect 12842 35238 13910 35248
rect 14757 35220 14767 36572
rect 14823 35220 14833 36572
rect 14757 35210 14833 35220
<< via2 >>
rect 6192 56366 6248 56422
rect 6316 56366 6372 56422
rect 6440 56366 6496 56422
rect 6564 56366 6620 56422
rect 6688 56366 6744 56422
rect 6812 56366 6868 56422
rect 6936 56366 6992 56422
rect 6192 56242 6248 56298
rect 6316 56242 6372 56298
rect 6440 56242 6496 56298
rect 6564 56242 6620 56298
rect 6688 56242 6744 56298
rect 6812 56242 6868 56298
rect 6936 56242 6992 56298
rect 6192 56118 6248 56174
rect 6316 56118 6372 56174
rect 6440 56118 6496 56174
rect 6564 56118 6620 56174
rect 6688 56118 6744 56174
rect 6812 56118 6868 56174
rect 6936 56118 6992 56174
rect 6192 55994 6248 56050
rect 6316 55994 6372 56050
rect 6440 55994 6496 56050
rect 6564 55994 6620 56050
rect 6688 55994 6744 56050
rect 6812 55994 6868 56050
rect 6936 55994 6992 56050
rect 6192 55870 6248 55926
rect 6316 55870 6372 55926
rect 6440 55870 6496 55926
rect 6564 55870 6620 55926
rect 6688 55870 6744 55926
rect 6812 55870 6868 55926
rect 6936 55870 6992 55926
rect 6192 55746 6248 55802
rect 6316 55746 6372 55802
rect 6440 55746 6496 55802
rect 6564 55746 6620 55802
rect 6688 55746 6744 55802
rect 6812 55746 6868 55802
rect 6936 55746 6992 55802
rect 6192 55622 6248 55678
rect 6316 55622 6372 55678
rect 6440 55622 6496 55678
rect 6564 55622 6620 55678
rect 6688 55622 6744 55678
rect 6812 55622 6868 55678
rect 6936 55622 6992 55678
rect 6192 55498 6248 55554
rect 6316 55498 6372 55554
rect 6440 55498 6496 55554
rect 6564 55498 6620 55554
rect 6688 55498 6744 55554
rect 6812 55498 6868 55554
rect 6936 55498 6992 55554
rect 6192 55374 6248 55430
rect 6316 55374 6372 55430
rect 6440 55374 6496 55430
rect 6564 55374 6620 55430
rect 6688 55374 6744 55430
rect 6812 55374 6868 55430
rect 6936 55374 6992 55430
rect 6192 55250 6248 55306
rect 6316 55250 6372 55306
rect 6440 55250 6496 55306
rect 6564 55250 6620 55306
rect 6688 55250 6744 55306
rect 6812 55250 6868 55306
rect 6936 55250 6992 55306
rect 6192 55126 6248 55182
rect 6316 55126 6372 55182
rect 6440 55126 6496 55182
rect 6564 55126 6620 55182
rect 6688 55126 6744 55182
rect 6812 55126 6868 55182
rect 6936 55126 6992 55182
rect 6192 55002 6248 55058
rect 6316 55002 6372 55058
rect 6440 55002 6496 55058
rect 6564 55002 6620 55058
rect 6688 55002 6744 55058
rect 6812 55002 6868 55058
rect 6936 55002 6992 55058
rect 6192 54878 6248 54934
rect 6316 54878 6372 54934
rect 6440 54878 6496 54934
rect 6564 54878 6620 54934
rect 6688 54878 6744 54934
rect 6812 54878 6868 54934
rect 6936 54878 6992 54934
rect 6192 54754 6248 54810
rect 6316 54754 6372 54810
rect 6440 54754 6496 54810
rect 6564 54754 6620 54810
rect 6688 54754 6744 54810
rect 6812 54754 6868 54810
rect 6936 54754 6992 54810
rect 6192 54630 6248 54686
rect 6316 54630 6372 54686
rect 6440 54630 6496 54686
rect 6564 54630 6620 54686
rect 6688 54630 6744 54686
rect 6812 54630 6868 54686
rect 6936 54630 6992 54686
rect 6192 54506 6248 54562
rect 6316 54506 6372 54562
rect 6440 54506 6496 54562
rect 6564 54506 6620 54562
rect 6688 54506 6744 54562
rect 6812 54506 6868 54562
rect 6936 54506 6992 54562
rect 6192 54382 6248 54438
rect 6316 54382 6372 54438
rect 6440 54382 6496 54438
rect 6564 54382 6620 54438
rect 6688 54382 6744 54438
rect 6812 54382 6868 54438
rect 6936 54382 6992 54438
rect 6192 54258 6248 54314
rect 6316 54258 6372 54314
rect 6440 54258 6496 54314
rect 6564 54258 6620 54314
rect 6688 54258 6744 54314
rect 6812 54258 6868 54314
rect 6936 54258 6992 54314
rect 6192 54134 6248 54190
rect 6316 54134 6372 54190
rect 6440 54134 6496 54190
rect 6564 54134 6620 54190
rect 6688 54134 6744 54190
rect 6812 54134 6868 54190
rect 6936 54134 6992 54190
rect 6192 54010 6248 54066
rect 6316 54010 6372 54066
rect 6440 54010 6496 54066
rect 6564 54010 6620 54066
rect 6688 54010 6744 54066
rect 6812 54010 6868 54066
rect 6936 54010 6992 54066
rect 6192 53886 6248 53942
rect 6316 53886 6372 53942
rect 6440 53886 6496 53942
rect 6564 53886 6620 53942
rect 6688 53886 6744 53942
rect 6812 53886 6868 53942
rect 6936 53886 6992 53942
rect 6192 53762 6248 53818
rect 6316 53762 6372 53818
rect 6440 53762 6496 53818
rect 6564 53762 6620 53818
rect 6688 53762 6744 53818
rect 6812 53762 6868 53818
rect 6936 53762 6992 53818
rect 6192 53638 6248 53694
rect 6316 53638 6372 53694
rect 6440 53638 6496 53694
rect 6564 53638 6620 53694
rect 6688 53638 6744 53694
rect 6812 53638 6868 53694
rect 6936 53638 6992 53694
rect 6192 53514 6248 53570
rect 6316 53514 6372 53570
rect 6440 53514 6496 53570
rect 6564 53514 6620 53570
rect 6688 53514 6744 53570
rect 6812 53514 6868 53570
rect 6936 53514 6992 53570
rect 6192 53390 6248 53446
rect 6316 53390 6372 53446
rect 6440 53390 6496 53446
rect 6564 53390 6620 53446
rect 6688 53390 6744 53446
rect 6812 53390 6868 53446
rect 6936 53390 6992 53446
rect 6192 53266 6248 53322
rect 6316 53266 6372 53322
rect 6440 53266 6496 53322
rect 6564 53266 6620 53322
rect 6688 53266 6744 53322
rect 6812 53266 6868 53322
rect 6936 53266 6992 53322
rect 7650 56377 7706 56433
rect 7774 56377 7830 56433
rect 7898 56377 7954 56433
rect 8022 56377 8078 56433
rect 8146 56377 8202 56433
rect 8270 56377 8326 56433
rect 8394 56377 8450 56433
rect 7650 56253 7706 56309
rect 7774 56253 7830 56309
rect 7898 56253 7954 56309
rect 8022 56253 8078 56309
rect 8146 56253 8202 56309
rect 8270 56253 8326 56309
rect 8394 56253 8450 56309
rect 7650 56129 7706 56185
rect 7774 56129 7830 56185
rect 7898 56129 7954 56185
rect 8022 56129 8078 56185
rect 8146 56129 8202 56185
rect 8270 56129 8326 56185
rect 8394 56129 8450 56185
rect 7650 56005 7706 56061
rect 7774 56005 7830 56061
rect 7898 56005 7954 56061
rect 8022 56005 8078 56061
rect 8146 56005 8202 56061
rect 8270 56005 8326 56061
rect 8394 56005 8450 56061
rect 7650 55881 7706 55937
rect 7774 55881 7830 55937
rect 7898 55881 7954 55937
rect 8022 55881 8078 55937
rect 8146 55881 8202 55937
rect 8270 55881 8326 55937
rect 8394 55881 8450 55937
rect 7650 55757 7706 55813
rect 7774 55757 7830 55813
rect 7898 55757 7954 55813
rect 8022 55757 8078 55813
rect 8146 55757 8202 55813
rect 8270 55757 8326 55813
rect 8394 55757 8450 55813
rect 7650 55633 7706 55689
rect 7774 55633 7830 55689
rect 7898 55633 7954 55689
rect 8022 55633 8078 55689
rect 8146 55633 8202 55689
rect 8270 55633 8326 55689
rect 8394 55633 8450 55689
rect 7650 55509 7706 55565
rect 7774 55509 7830 55565
rect 7898 55509 7954 55565
rect 8022 55509 8078 55565
rect 8146 55509 8202 55565
rect 8270 55509 8326 55565
rect 8394 55509 8450 55565
rect 7650 55385 7706 55441
rect 7774 55385 7830 55441
rect 7898 55385 7954 55441
rect 8022 55385 8078 55441
rect 8146 55385 8202 55441
rect 8270 55385 8326 55441
rect 8394 55385 8450 55441
rect 7650 55261 7706 55317
rect 7774 55261 7830 55317
rect 7898 55261 7954 55317
rect 8022 55261 8078 55317
rect 8146 55261 8202 55317
rect 8270 55261 8326 55317
rect 8394 55261 8450 55317
rect 7650 55137 7706 55193
rect 7774 55137 7830 55193
rect 7898 55137 7954 55193
rect 8022 55137 8078 55193
rect 8146 55137 8202 55193
rect 8270 55137 8326 55193
rect 8394 55137 8450 55193
rect 7650 55013 7706 55069
rect 7774 55013 7830 55069
rect 7898 55013 7954 55069
rect 8022 55013 8078 55069
rect 8146 55013 8202 55069
rect 8270 55013 8326 55069
rect 8394 55013 8450 55069
rect 7650 54889 7706 54945
rect 7774 54889 7830 54945
rect 7898 54889 7954 54945
rect 8022 54889 8078 54945
rect 8146 54889 8202 54945
rect 8270 54889 8326 54945
rect 8394 54889 8450 54945
rect 7650 54765 7706 54821
rect 7774 54765 7830 54821
rect 7898 54765 7954 54821
rect 8022 54765 8078 54821
rect 8146 54765 8202 54821
rect 8270 54765 8326 54821
rect 8394 54765 8450 54821
rect 7650 54641 7706 54697
rect 7774 54641 7830 54697
rect 7898 54641 7954 54697
rect 8022 54641 8078 54697
rect 8146 54641 8202 54697
rect 8270 54641 8326 54697
rect 8394 54641 8450 54697
rect 7650 54517 7706 54573
rect 7774 54517 7830 54573
rect 7898 54517 7954 54573
rect 8022 54517 8078 54573
rect 8146 54517 8202 54573
rect 8270 54517 8326 54573
rect 8394 54517 8450 54573
rect 7650 54393 7706 54449
rect 7774 54393 7830 54449
rect 7898 54393 7954 54449
rect 8022 54393 8078 54449
rect 8146 54393 8202 54449
rect 8270 54393 8326 54449
rect 8394 54393 8450 54449
rect 7650 54269 7706 54325
rect 7774 54269 7830 54325
rect 7898 54269 7954 54325
rect 8022 54269 8078 54325
rect 8146 54269 8202 54325
rect 8270 54269 8326 54325
rect 8394 54269 8450 54325
rect 7650 54145 7706 54201
rect 7774 54145 7830 54201
rect 7898 54145 7954 54201
rect 8022 54145 8078 54201
rect 8146 54145 8202 54201
rect 8270 54145 8326 54201
rect 8394 54145 8450 54201
rect 7650 54021 7706 54077
rect 7774 54021 7830 54077
rect 7898 54021 7954 54077
rect 8022 54021 8078 54077
rect 8146 54021 8202 54077
rect 8270 54021 8326 54077
rect 8394 54021 8450 54077
rect 7650 53897 7706 53953
rect 7774 53897 7830 53953
rect 7898 53897 7954 53953
rect 8022 53897 8078 53953
rect 8146 53897 8202 53953
rect 8270 53897 8326 53953
rect 8394 53897 8450 53953
rect 7650 53773 7706 53829
rect 7774 53773 7830 53829
rect 7898 53773 7954 53829
rect 8022 53773 8078 53829
rect 8146 53773 8202 53829
rect 8270 53773 8326 53829
rect 8394 53773 8450 53829
rect 7650 53649 7706 53705
rect 7774 53649 7830 53705
rect 7898 53649 7954 53705
rect 8022 53649 8078 53705
rect 8146 53649 8202 53705
rect 8270 53649 8326 53705
rect 8394 53649 8450 53705
rect 7650 53525 7706 53581
rect 7774 53525 7830 53581
rect 7898 53525 7954 53581
rect 8022 53525 8078 53581
rect 8146 53525 8202 53581
rect 8270 53525 8326 53581
rect 8394 53525 8450 53581
rect 7650 53401 7706 53457
rect 7774 53401 7830 53457
rect 7898 53401 7954 53457
rect 8022 53401 8078 53457
rect 8146 53401 8202 53457
rect 8270 53401 8326 53457
rect 8394 53401 8450 53457
rect 7650 53277 7706 53333
rect 7774 53277 7830 53333
rect 7898 53277 7954 53333
rect 8022 53277 8078 53333
rect 8146 53277 8202 53333
rect 8270 53277 8326 53333
rect 8394 53277 8450 53333
rect 7650 53153 7706 53209
rect 7774 53153 7830 53209
rect 7898 53153 7954 53209
rect 8022 53153 8078 53209
rect 8146 53153 8202 53209
rect 8270 53153 8326 53209
rect 8394 53153 8450 53209
rect 7650 53029 7706 53085
rect 7774 53029 7830 53085
rect 7898 53029 7954 53085
rect 8022 53029 8078 53085
rect 8146 53029 8202 53085
rect 8270 53029 8326 53085
rect 8394 53029 8450 53085
rect 7650 52905 7706 52961
rect 7774 52905 7830 52961
rect 7898 52905 7954 52961
rect 8022 52905 8078 52961
rect 8146 52905 8202 52961
rect 8270 52905 8326 52961
rect 8394 52905 8450 52961
rect 7650 52781 7706 52837
rect 7774 52781 7830 52837
rect 7898 52781 7954 52837
rect 8022 52781 8078 52837
rect 8146 52781 8202 52837
rect 8270 52781 8326 52837
rect 8394 52781 8450 52837
rect 8812 52681 8868 52737
rect 8936 52681 8992 52737
rect 9060 52681 9116 52737
rect 9184 52681 9240 52737
rect 9308 52681 9364 52737
rect 9432 52681 9488 52737
rect 8812 52557 8868 52613
rect 8936 52557 8992 52613
rect 9060 52557 9116 52613
rect 9184 52557 9240 52613
rect 9308 52557 9364 52613
rect 9432 52557 9488 52613
rect 8812 52433 8868 52489
rect 8936 52433 8992 52489
rect 9060 52433 9116 52489
rect 9184 52433 9240 52489
rect 9308 52433 9364 52489
rect 9432 52433 9488 52489
rect 8812 52309 8868 52365
rect 8936 52309 8992 52365
rect 9060 52309 9116 52365
rect 9184 52309 9240 52365
rect 9308 52309 9364 52365
rect 9432 52309 9488 52365
rect 8812 52185 8868 52241
rect 8936 52185 8992 52241
rect 9060 52185 9116 52241
rect 9184 52185 9240 52241
rect 9308 52185 9364 52241
rect 9432 52185 9488 52241
rect 8812 52061 8868 52117
rect 8936 52061 8992 52117
rect 9060 52061 9116 52117
rect 9184 52061 9240 52117
rect 9308 52061 9364 52117
rect 9432 52061 9488 52117
rect 8812 51937 8868 51993
rect 8936 51937 8992 51993
rect 9060 51937 9116 51993
rect 9184 51937 9240 51993
rect 9308 51937 9364 51993
rect 9432 51937 9488 51993
rect 8812 51813 8868 51869
rect 8936 51813 8992 51869
rect 9060 51813 9116 51869
rect 9184 51813 9240 51869
rect 9308 51813 9364 51869
rect 9432 51813 9488 51869
rect 8812 51689 8868 51745
rect 8936 51689 8992 51745
rect 9060 51689 9116 51745
rect 9184 51689 9240 51745
rect 9308 51689 9364 51745
rect 9432 51689 9488 51745
rect 8812 51565 8868 51621
rect 8936 51565 8992 51621
rect 9060 51565 9116 51621
rect 9184 51565 9240 51621
rect 9308 51565 9364 51621
rect 9432 51565 9488 51621
rect 7650 51396 7706 51452
rect 7774 51396 7830 51452
rect 7898 51396 7954 51452
rect 8022 51396 8078 51452
rect 8146 51396 8202 51452
rect 8270 51396 8326 51452
rect 8394 51396 8450 51452
rect 7650 51272 7706 51328
rect 7774 51272 7830 51328
rect 7898 51272 7954 51328
rect 8022 51272 8078 51328
rect 8146 51272 8202 51328
rect 8270 51272 8326 51328
rect 8394 51272 8450 51328
rect 7650 51148 7706 51204
rect 7774 51148 7830 51204
rect 7898 51148 7954 51204
rect 8022 51148 8078 51204
rect 8146 51148 8202 51204
rect 8270 51148 8326 51204
rect 8394 51148 8450 51204
rect 7650 51024 7706 51080
rect 7774 51024 7830 51080
rect 7898 51024 7954 51080
rect 8022 51024 8078 51080
rect 8146 51024 8202 51080
rect 8270 51024 8326 51080
rect 8394 51024 8450 51080
rect 7650 50900 7706 50956
rect 7774 50900 7830 50956
rect 7898 50900 7954 50956
rect 8022 50900 8078 50956
rect 8146 50900 8202 50956
rect 8270 50900 8326 50956
rect 8394 50900 8450 50956
rect 7650 50776 7706 50832
rect 7774 50776 7830 50832
rect 7898 50776 7954 50832
rect 8022 50776 8078 50832
rect 8146 50776 8202 50832
rect 8270 50776 8326 50832
rect 8394 50776 8450 50832
rect 7650 50652 7706 50708
rect 7774 50652 7830 50708
rect 7898 50652 7954 50708
rect 8022 50652 8078 50708
rect 8146 50652 8202 50708
rect 8270 50652 8326 50708
rect 8394 50652 8450 50708
rect 7650 50528 7706 50584
rect 7774 50528 7830 50584
rect 7898 50528 7954 50584
rect 8022 50528 8078 50584
rect 8146 50528 8202 50584
rect 8270 50528 8326 50584
rect 8394 50528 8450 50584
rect 1104 42834 1160 42890
rect 1104 42710 1160 42766
rect 1104 42586 1160 42642
rect 1104 42462 1160 42518
rect 1104 42338 1160 42394
rect 1104 42214 1160 42270
rect 1104 42090 1160 42146
rect 1104 41966 1160 42022
rect 1104 41842 1160 41898
rect 1104 41718 1160 41774
rect 1104 41594 1160 41650
rect 1104 41470 1160 41526
rect 1104 41346 1160 41402
rect 1104 41222 1160 41278
rect 1228 42710 1284 42766
rect 1228 42586 1284 42642
rect 1228 42462 1284 42518
rect 1228 42338 1284 42394
rect 1228 42214 1284 42270
rect 1228 42090 1284 42146
rect 1228 41966 1284 42022
rect 1228 41842 1284 41898
rect 1228 41718 1284 41774
rect 1228 41594 1284 41650
rect 1228 41470 1284 41526
rect 1228 41346 1284 41402
rect 1228 41222 1284 41278
rect 1228 41098 1284 41154
rect 1352 42586 1408 42642
rect 1352 42462 1408 42518
rect 1352 42338 1408 42394
rect 1352 42214 1408 42270
rect 1352 42090 1408 42146
rect 1352 41966 1408 42022
rect 1352 41842 1408 41898
rect 1352 41718 1408 41774
rect 1352 41594 1408 41650
rect 1352 41470 1408 41526
rect 1352 41346 1408 41402
rect 1352 41222 1408 41278
rect 1352 41098 1408 41154
rect 1352 40974 1408 41030
rect 1476 42462 1532 42518
rect 1476 42338 1532 42394
rect 1476 42214 1532 42270
rect 1476 42090 1532 42146
rect 1476 41966 1532 42022
rect 1476 41842 1532 41898
rect 1476 41718 1532 41774
rect 1476 41594 1532 41650
rect 1476 41470 1532 41526
rect 1476 41346 1532 41402
rect 1476 41222 1532 41278
rect 1476 41098 1532 41154
rect 1476 40974 1532 41030
rect 1476 40850 1532 40906
rect 1600 42338 1656 42394
rect 1600 42214 1656 42270
rect 1600 42090 1656 42146
rect 1600 41966 1656 42022
rect 1600 41842 1656 41898
rect 1600 41718 1656 41774
rect 1600 41594 1656 41650
rect 1600 41470 1656 41526
rect 1600 41346 1656 41402
rect 1600 41222 1656 41278
rect 1600 41098 1656 41154
rect 1600 40974 1656 41030
rect 1600 40850 1656 40906
rect 1600 40726 1656 40782
rect 1724 42214 1780 42270
rect 1724 42090 1780 42146
rect 1724 41966 1780 42022
rect 1724 41842 1780 41898
rect 1724 41718 1780 41774
rect 1724 41594 1780 41650
rect 1724 41470 1780 41526
rect 1724 41346 1780 41402
rect 1724 41222 1780 41278
rect 1724 41098 1780 41154
rect 1724 40974 1780 41030
rect 1724 40850 1780 40906
rect 1724 40726 1780 40782
rect 1724 40602 1780 40658
rect 1848 42090 1904 42146
rect 1848 41966 1904 42022
rect 1848 41842 1904 41898
rect 1848 41718 1904 41774
rect 1848 41594 1904 41650
rect 1848 41470 1904 41526
rect 1848 41346 1904 41402
rect 1848 41222 1904 41278
rect 1848 41098 1904 41154
rect 1848 40974 1904 41030
rect 1848 40850 1904 40906
rect 1848 40726 1904 40782
rect 1848 40602 1904 40658
rect 1848 40478 1904 40534
rect 1972 41966 2028 42022
rect 1972 41842 2028 41898
rect 1972 41718 2028 41774
rect 12852 50882 12908 50938
rect 12976 50882 13032 50938
rect 13100 50882 13156 50938
rect 13224 50882 13280 50938
rect 13348 50882 13404 50938
rect 13472 50882 13528 50938
rect 13596 50882 13652 50938
rect 13720 50882 13776 50938
rect 13844 50882 13900 50938
rect 12852 50758 12908 50814
rect 12976 50758 13032 50814
rect 13100 50758 13156 50814
rect 13224 50758 13280 50814
rect 13348 50758 13404 50814
rect 13472 50758 13528 50814
rect 13596 50758 13652 50814
rect 13720 50758 13776 50814
rect 13844 50758 13900 50814
rect 12852 50634 12908 50690
rect 12976 50634 13032 50690
rect 13100 50634 13156 50690
rect 13224 50634 13280 50690
rect 13348 50634 13404 50690
rect 13472 50634 13528 50690
rect 13596 50634 13652 50690
rect 13720 50634 13776 50690
rect 13844 50634 13900 50690
rect 12852 50510 12908 50566
rect 12976 50510 13032 50566
rect 13100 50510 13156 50566
rect 13224 50510 13280 50566
rect 13348 50510 13404 50566
rect 13472 50510 13528 50566
rect 13596 50510 13652 50566
rect 13720 50510 13776 50566
rect 13844 50510 13900 50566
rect 12852 50386 12908 50442
rect 12976 50386 13032 50442
rect 13100 50386 13156 50442
rect 13224 50386 13280 50442
rect 13348 50386 13404 50442
rect 13472 50386 13528 50442
rect 13596 50386 13652 50442
rect 13720 50386 13776 50442
rect 13844 50386 13900 50442
rect 12852 50262 12908 50318
rect 12976 50262 13032 50318
rect 13100 50262 13156 50318
rect 13224 50262 13280 50318
rect 13348 50262 13404 50318
rect 13472 50262 13528 50318
rect 13596 50262 13652 50318
rect 13720 50262 13776 50318
rect 13844 50262 13900 50318
rect 12852 50138 12908 50194
rect 12976 50138 13032 50194
rect 13100 50138 13156 50194
rect 13224 50138 13280 50194
rect 13348 50138 13404 50194
rect 13472 50138 13528 50194
rect 13596 50138 13652 50194
rect 13720 50138 13776 50194
rect 13844 50138 13900 50194
rect 12852 50014 12908 50070
rect 12976 50014 13032 50070
rect 13100 50014 13156 50070
rect 13224 50014 13280 50070
rect 13348 50014 13404 50070
rect 13472 50014 13528 50070
rect 13596 50014 13652 50070
rect 13720 50014 13776 50070
rect 13844 50014 13900 50070
rect 12852 49890 12908 49946
rect 12976 49890 13032 49946
rect 13100 49890 13156 49946
rect 13224 49890 13280 49946
rect 13348 49890 13404 49946
rect 13472 49890 13528 49946
rect 13596 49890 13652 49946
rect 13720 49890 13776 49946
rect 13844 49890 13900 49946
rect 12852 49766 12908 49822
rect 12976 49766 13032 49822
rect 13100 49766 13156 49822
rect 13224 49766 13280 49822
rect 13348 49766 13404 49822
rect 13472 49766 13528 49822
rect 13596 49766 13652 49822
rect 13720 49766 13776 49822
rect 13844 49766 13900 49822
rect 12852 49642 12908 49698
rect 12976 49642 13032 49698
rect 13100 49642 13156 49698
rect 13224 49642 13280 49698
rect 13348 49642 13404 49698
rect 13472 49642 13528 49698
rect 13596 49642 13652 49698
rect 13720 49642 13776 49698
rect 13844 49642 13900 49698
rect 14767 50970 14823 50972
rect 14767 50918 14769 50970
rect 14769 50918 14821 50970
rect 14821 50918 14823 50970
rect 14767 50862 14823 50918
rect 14767 50810 14769 50862
rect 14769 50810 14821 50862
rect 14821 50810 14823 50862
rect 14767 50754 14823 50810
rect 14767 50702 14769 50754
rect 14769 50702 14821 50754
rect 14821 50702 14823 50754
rect 14767 50646 14823 50702
rect 14767 50594 14769 50646
rect 14769 50594 14821 50646
rect 14821 50594 14823 50646
rect 14767 50538 14823 50594
rect 14767 50486 14769 50538
rect 14769 50486 14821 50538
rect 14821 50486 14823 50538
rect 14767 50430 14823 50486
rect 14767 50378 14769 50430
rect 14769 50378 14821 50430
rect 14821 50378 14823 50430
rect 14767 50322 14823 50378
rect 14767 50270 14769 50322
rect 14769 50270 14821 50322
rect 14821 50270 14823 50322
rect 14767 50214 14823 50270
rect 14767 50162 14769 50214
rect 14769 50162 14821 50214
rect 14821 50162 14823 50214
rect 14767 50106 14823 50162
rect 14767 50054 14769 50106
rect 14769 50054 14821 50106
rect 14821 50054 14823 50106
rect 14767 49998 14823 50054
rect 14767 49946 14769 49998
rect 14769 49946 14821 49998
rect 14821 49946 14823 49998
rect 14767 49890 14823 49946
rect 14767 49838 14769 49890
rect 14769 49838 14821 49890
rect 14821 49838 14823 49890
rect 14767 49782 14823 49838
rect 14767 49730 14769 49782
rect 14769 49730 14821 49782
rect 14821 49730 14823 49782
rect 14767 49674 14823 49730
rect 14767 49622 14769 49674
rect 14769 49622 14821 49674
rect 14821 49622 14823 49674
rect 14767 49620 14823 49622
rect 10679 49290 10735 49346
rect 10803 49290 10859 49346
rect 10927 49290 10983 49346
rect 11051 49290 11107 49346
rect 11175 49290 11231 49346
rect 11299 49290 11355 49346
rect 11423 49290 11479 49346
rect 11547 49290 11603 49346
rect 11671 49290 11727 49346
rect 11795 49290 11851 49346
rect 11919 49290 11975 49346
rect 12043 49290 12099 49346
rect 12167 49290 12223 49346
rect 12291 49290 12347 49346
rect 12415 49290 12471 49346
rect 10679 49166 10735 49222
rect 10803 49166 10859 49222
rect 10927 49166 10983 49222
rect 11051 49166 11107 49222
rect 11175 49166 11231 49222
rect 11299 49166 11355 49222
rect 11423 49166 11479 49222
rect 11547 49166 11603 49222
rect 11671 49166 11727 49222
rect 11795 49166 11851 49222
rect 11919 49166 11975 49222
rect 12043 49166 12099 49222
rect 12167 49166 12223 49222
rect 12291 49166 12347 49222
rect 12415 49166 12471 49222
rect 10679 49042 10735 49098
rect 10803 49042 10859 49098
rect 10927 49042 10983 49098
rect 11051 49042 11107 49098
rect 11175 49042 11231 49098
rect 11299 49042 11355 49098
rect 11423 49042 11479 49098
rect 11547 49042 11603 49098
rect 11671 49042 11727 49098
rect 11795 49042 11851 49098
rect 11919 49042 11975 49098
rect 12043 49042 12099 49098
rect 12167 49042 12223 49098
rect 12291 49042 12347 49098
rect 12415 49042 12471 49098
rect 10679 48918 10735 48974
rect 10803 48918 10859 48974
rect 10927 48918 10983 48974
rect 11051 48918 11107 48974
rect 11175 48918 11231 48974
rect 11299 48918 11355 48974
rect 11423 48918 11479 48974
rect 11547 48918 11603 48974
rect 11671 48918 11727 48974
rect 11795 48918 11851 48974
rect 11919 48918 11975 48974
rect 12043 48918 12099 48974
rect 12167 48918 12223 48974
rect 12291 48918 12347 48974
rect 12415 48918 12471 48974
rect 10679 48794 10735 48850
rect 10803 48794 10859 48850
rect 10927 48794 10983 48850
rect 11051 48794 11107 48850
rect 11175 48794 11231 48850
rect 11299 48794 11355 48850
rect 11423 48794 11479 48850
rect 11547 48794 11603 48850
rect 11671 48794 11727 48850
rect 11795 48794 11851 48850
rect 11919 48794 11975 48850
rect 12043 48794 12099 48850
rect 12167 48794 12223 48850
rect 12291 48794 12347 48850
rect 12415 48794 12471 48850
rect 10679 48670 10735 48726
rect 10803 48670 10859 48726
rect 10927 48670 10983 48726
rect 11051 48670 11107 48726
rect 11175 48670 11231 48726
rect 11299 48670 11355 48726
rect 11423 48670 11479 48726
rect 11547 48670 11603 48726
rect 11671 48670 11727 48726
rect 11795 48670 11851 48726
rect 11919 48670 11975 48726
rect 12043 48670 12099 48726
rect 12167 48670 12223 48726
rect 12291 48670 12347 48726
rect 12415 48670 12471 48726
rect 10679 48546 10735 48602
rect 10803 48546 10859 48602
rect 10927 48546 10983 48602
rect 11051 48546 11107 48602
rect 11175 48546 11231 48602
rect 11299 48546 11355 48602
rect 11423 48546 11479 48602
rect 11547 48546 11603 48602
rect 11671 48546 11727 48602
rect 11795 48546 11851 48602
rect 11919 48546 11975 48602
rect 12043 48546 12099 48602
rect 12167 48546 12223 48602
rect 12291 48546 12347 48602
rect 12415 48546 12471 48602
rect 10679 48422 10735 48478
rect 10803 48422 10859 48478
rect 10927 48422 10983 48478
rect 11051 48422 11107 48478
rect 11175 48422 11231 48478
rect 11299 48422 11355 48478
rect 11423 48422 11479 48478
rect 11547 48422 11603 48478
rect 11671 48422 11727 48478
rect 11795 48422 11851 48478
rect 11919 48422 11975 48478
rect 12043 48422 12099 48478
rect 12167 48422 12223 48478
rect 12291 48422 12347 48478
rect 12415 48422 12471 48478
rect 10679 48298 10735 48354
rect 10803 48298 10859 48354
rect 10927 48298 10983 48354
rect 11051 48298 11107 48354
rect 11175 48298 11231 48354
rect 11299 48298 11355 48354
rect 11423 48298 11479 48354
rect 11547 48298 11603 48354
rect 11671 48298 11727 48354
rect 11795 48298 11851 48354
rect 11919 48298 11975 48354
rect 12043 48298 12099 48354
rect 12167 48298 12223 48354
rect 12291 48298 12347 48354
rect 12415 48298 12471 48354
rect 10679 48174 10735 48230
rect 10803 48174 10859 48230
rect 10927 48174 10983 48230
rect 11051 48174 11107 48230
rect 11175 48174 11231 48230
rect 11299 48174 11355 48230
rect 11423 48174 11479 48230
rect 11547 48174 11603 48230
rect 11671 48174 11727 48230
rect 11795 48174 11851 48230
rect 11919 48174 11975 48230
rect 12043 48174 12099 48230
rect 12167 48174 12223 48230
rect 12291 48174 12347 48230
rect 12415 48174 12471 48230
rect 10679 48050 10735 48106
rect 10803 48050 10859 48106
rect 10927 48050 10983 48106
rect 11051 48050 11107 48106
rect 11175 48050 11231 48106
rect 11299 48050 11355 48106
rect 11423 48050 11479 48106
rect 11547 48050 11603 48106
rect 11671 48050 11727 48106
rect 11795 48050 11851 48106
rect 11919 48050 11975 48106
rect 12043 48050 12099 48106
rect 12167 48050 12223 48106
rect 12291 48050 12347 48106
rect 12415 48050 12471 48106
rect 1972 41594 2028 41650
rect 1972 41470 2028 41526
rect 1972 41346 2028 41402
rect 1972 41222 2028 41278
rect 1972 41098 2028 41154
rect 1972 40974 2028 41030
rect 1972 40850 2028 40906
rect 1972 40726 2028 40782
rect 1972 40602 2028 40658
rect 1972 40478 2028 40534
rect 1972 40354 2028 40410
rect 4470 39468 4526 39524
rect 4470 39344 4526 39400
rect 4470 39220 4526 39276
rect 2527 39149 2583 39205
rect 4470 39096 4526 39152
rect 2527 39025 2583 39081
rect 2527 38901 2583 38957
rect 2527 38777 2583 38833
rect 2527 38653 2583 38709
rect 2527 38529 2583 38585
rect 2527 38405 2583 38461
rect 2527 38281 2583 38337
rect 2527 38157 2583 38213
rect 2527 38033 2583 38089
rect 2527 37909 2583 37965
rect 2527 37785 2583 37841
rect 2527 37661 2583 37717
rect 2527 37537 2583 37593
rect 2651 39025 2707 39081
rect 4470 38972 4526 39028
rect 2651 38901 2707 38957
rect 2651 38777 2707 38833
rect 2651 38653 2707 38709
rect 2651 38529 2707 38585
rect 2651 38405 2707 38461
rect 2651 38281 2707 38337
rect 2651 38157 2707 38213
rect 2651 38033 2707 38089
rect 2651 37909 2707 37965
rect 2651 37785 2707 37841
rect 2651 37661 2707 37717
rect 2651 37537 2707 37593
rect 2651 37413 2707 37469
rect 2775 38901 2831 38957
rect 4470 38848 4526 38904
rect 2775 38777 2831 38833
rect 2775 38653 2831 38709
rect 2775 38529 2831 38585
rect 2775 38405 2831 38461
rect 2775 38281 2831 38337
rect 2775 38157 2831 38213
rect 2775 38033 2831 38089
rect 2775 37909 2831 37965
rect 2775 37785 2831 37841
rect 2775 37661 2831 37717
rect 2775 37537 2831 37593
rect 2775 37413 2831 37469
rect 2775 37289 2831 37345
rect 2899 38777 2955 38833
rect 4470 38724 4526 38780
rect 2899 38653 2955 38709
rect 2899 38529 2955 38585
rect 2899 38405 2955 38461
rect 2899 38281 2955 38337
rect 2899 38157 2955 38213
rect 2899 38033 2955 38089
rect 2899 37909 2955 37965
rect 2899 37785 2955 37841
rect 2899 37661 2955 37717
rect 2899 37537 2955 37593
rect 2899 37413 2955 37469
rect 2899 37289 2955 37345
rect 2899 37165 2955 37221
rect 3023 38653 3079 38709
rect 4470 38600 4526 38656
rect 3023 38529 3079 38585
rect 3023 38405 3079 38461
rect 3023 38281 3079 38337
rect 3023 38157 3079 38213
rect 3023 38033 3079 38089
rect 3023 37909 3079 37965
rect 3023 37785 3079 37841
rect 3023 37661 3079 37717
rect 3023 37537 3079 37593
rect 3023 37413 3079 37469
rect 3023 37289 3079 37345
rect 3023 37165 3079 37221
rect 3023 37041 3079 37097
rect 3147 38529 3203 38585
rect 4470 38476 4526 38532
rect 3147 38405 3203 38461
rect 3147 38281 3203 38337
rect 3147 38157 3203 38213
rect 3147 38033 3203 38089
rect 3147 37909 3203 37965
rect 3147 37785 3203 37841
rect 3147 37661 3203 37717
rect 3147 37537 3203 37593
rect 3147 37413 3203 37469
rect 3147 37289 3203 37345
rect 3147 37165 3203 37221
rect 3147 37041 3203 37097
rect 3147 36917 3203 36973
rect 3271 38405 3327 38461
rect 4470 38352 4526 38408
rect 3271 38281 3327 38337
rect 3271 38157 3327 38213
rect 3271 38033 3327 38089
rect 3271 37909 3327 37965
rect 3271 37785 3327 37841
rect 3271 37661 3327 37717
rect 3271 37537 3327 37593
rect 3271 37413 3327 37469
rect 3271 37289 3327 37345
rect 3271 37165 3327 37221
rect 3271 37041 3327 37097
rect 3271 36917 3327 36973
rect 3271 36793 3327 36849
rect 3395 38281 3451 38337
rect 4470 38228 4526 38284
rect 3395 38157 3451 38213
rect 3395 38033 3451 38089
rect 3395 37909 3451 37965
rect 3395 37785 3451 37841
rect 3395 37661 3451 37717
rect 3395 37537 3451 37593
rect 3395 37413 3451 37469
rect 3395 37289 3451 37345
rect 3395 37165 3451 37221
rect 3395 37041 3451 37097
rect 3395 36917 3451 36973
rect 3395 36793 3451 36849
rect 3395 36669 3451 36725
rect 3519 38157 3575 38213
rect 4470 38104 4526 38160
rect 3519 38033 3575 38089
rect 3519 37909 3575 37965
rect 3519 37785 3575 37841
rect 3519 37661 3575 37717
rect 3519 37537 3575 37593
rect 3519 37413 3575 37469
rect 3519 37289 3575 37345
rect 3519 37165 3575 37221
rect 3519 37041 3575 37097
rect 3519 36917 3575 36973
rect 3519 36793 3575 36849
rect 3519 36669 3575 36725
rect 3519 36545 3575 36601
rect 3643 38033 3699 38089
rect 4470 37980 4526 38036
rect 3643 37909 3699 37965
rect 3643 37785 3699 37841
rect 3643 37661 3699 37717
rect 3643 37537 3699 37593
rect 3643 37413 3699 37469
rect 3643 37289 3699 37345
rect 3643 37165 3699 37221
rect 3643 37041 3699 37097
rect 3643 36917 3699 36973
rect 3643 36793 3699 36849
rect 3643 36669 3699 36725
rect 3643 36545 3699 36601
rect 3643 36421 3699 36477
rect 3767 37909 3823 37965
rect 4470 37856 4526 37912
rect 3767 37785 3823 37841
rect 3767 37661 3823 37717
rect 3767 37537 3823 37593
rect 3767 37413 3823 37469
rect 3767 37289 3823 37345
rect 3767 37165 3823 37221
rect 3767 37041 3823 37097
rect 3767 36917 3823 36973
rect 3767 36793 3823 36849
rect 3767 36669 3823 36725
rect 3767 36545 3823 36601
rect 3767 36421 3823 36477
rect 3767 36297 3823 36353
rect 4594 39344 4650 39400
rect 4594 39220 4650 39276
rect 4594 39096 4650 39152
rect 4594 38972 4650 39028
rect 4594 38848 4650 38904
rect 4594 38724 4650 38780
rect 4594 38600 4650 38656
rect 4594 38476 4650 38532
rect 4594 38352 4650 38408
rect 4594 38228 4650 38284
rect 4594 38104 4650 38160
rect 4594 37980 4650 38036
rect 4594 37856 4650 37912
rect 3891 37785 3947 37841
rect 4594 37732 4650 37788
rect 3891 37661 3947 37717
rect 3891 37537 3947 37593
rect 3891 37413 3947 37469
rect 3891 37289 3947 37345
rect 3891 37165 3947 37221
rect 3891 37041 3947 37097
rect 3891 36917 3947 36973
rect 3891 36793 3947 36849
rect 3891 36669 3947 36725
rect 3891 36545 3947 36601
rect 3891 36421 3947 36477
rect 3891 36297 3947 36353
rect 3891 36173 3947 36229
rect 4718 39220 4774 39276
rect 4718 39096 4774 39152
rect 4718 38972 4774 39028
rect 4718 38848 4774 38904
rect 4718 38724 4774 38780
rect 4718 38600 4774 38656
rect 4718 38476 4774 38532
rect 4718 38352 4774 38408
rect 4718 38228 4774 38284
rect 4718 38104 4774 38160
rect 4718 37980 4774 38036
rect 4718 37856 4774 37912
rect 4718 37732 4774 37788
rect 4015 37661 4071 37717
rect 4718 37608 4774 37664
rect 4015 37537 4071 37593
rect 4015 37413 4071 37469
rect 4015 37289 4071 37345
rect 4015 37165 4071 37221
rect 4015 37041 4071 37097
rect 4015 36917 4071 36973
rect 4015 36793 4071 36849
rect 4015 36669 4071 36725
rect 4015 36545 4071 36601
rect 4015 36421 4071 36477
rect 4015 36297 4071 36353
rect 4015 36173 4071 36229
rect 4015 36049 4071 36105
rect 4842 39096 4898 39152
rect 4842 38972 4898 39028
rect 4842 38848 4898 38904
rect 4842 38724 4898 38780
rect 4842 38600 4898 38656
rect 4842 38476 4898 38532
rect 4842 38352 4898 38408
rect 4842 38228 4898 38284
rect 4842 38104 4898 38160
rect 4842 37980 4898 38036
rect 4842 37856 4898 37912
rect 4842 37732 4898 37788
rect 4842 37608 4898 37664
rect 4139 37537 4195 37593
rect 4842 37484 4898 37540
rect 4966 38972 5022 39028
rect 4966 38848 5022 38904
rect 4966 38724 5022 38780
rect 4966 38600 5022 38656
rect 4966 38476 5022 38532
rect 4966 38352 5022 38408
rect 4966 38228 5022 38284
rect 4966 38104 5022 38160
rect 4966 37980 5022 38036
rect 4966 37856 5022 37912
rect 4966 37732 5022 37788
rect 4966 37608 5022 37664
rect 4966 37484 5022 37540
rect 4139 37413 4195 37469
rect 4966 37360 5022 37416
rect 5090 38848 5146 38904
rect 5090 38724 5146 38780
rect 5090 38600 5146 38656
rect 5090 38476 5146 38532
rect 5090 38352 5146 38408
rect 5090 38228 5146 38284
rect 5090 38104 5146 38160
rect 5090 37980 5146 38036
rect 5090 37856 5146 37912
rect 5090 37732 5146 37788
rect 5090 37608 5146 37664
rect 5090 37484 5146 37540
rect 5090 37360 5146 37416
rect 4139 37289 4195 37345
rect 5090 37236 5146 37292
rect 5214 38724 5270 38780
rect 5214 38600 5270 38656
rect 5214 38476 5270 38532
rect 5214 38352 5270 38408
rect 5214 38228 5270 38284
rect 5214 38104 5270 38160
rect 5214 37980 5270 38036
rect 5214 37856 5270 37912
rect 5214 37732 5270 37788
rect 5214 37608 5270 37664
rect 5214 37484 5270 37540
rect 5214 37360 5270 37416
rect 5214 37236 5270 37292
rect 4139 37165 4195 37221
rect 5214 37112 5270 37168
rect 5338 38600 5394 38656
rect 5338 38476 5394 38532
rect 5338 38352 5394 38408
rect 5338 38228 5394 38284
rect 5338 38104 5394 38160
rect 5338 37980 5394 38036
rect 5338 37856 5394 37912
rect 5338 37732 5394 37788
rect 5338 37608 5394 37664
rect 5338 37484 5394 37540
rect 5338 37360 5394 37416
rect 5338 37236 5394 37292
rect 5338 37112 5394 37168
rect 4139 37041 4195 37097
rect 5338 36988 5394 37044
rect 5462 38476 5518 38532
rect 5462 38352 5518 38408
rect 5462 38228 5518 38284
rect 5462 38104 5518 38160
rect 5462 37980 5518 38036
rect 5462 37856 5518 37912
rect 5462 37732 5518 37788
rect 5462 37608 5518 37664
rect 5462 37484 5518 37540
rect 5462 37360 5518 37416
rect 5462 37236 5518 37292
rect 5462 37112 5518 37168
rect 5462 36988 5518 37044
rect 4139 36917 4195 36973
rect 5462 36864 5518 36920
rect 5586 38346 5642 38402
rect 5586 38222 5642 38278
rect 5586 38098 5642 38154
rect 5586 37974 5642 38030
rect 5586 37850 5642 37906
rect 5586 37726 5642 37782
rect 5586 37602 5642 37658
rect 5586 37478 5642 37534
rect 5586 37354 5642 37410
rect 5586 37230 5642 37286
rect 5586 37106 5642 37162
rect 5586 36982 5642 37038
rect 5586 36858 5642 36914
rect 4139 36793 4195 36849
rect 5710 38217 5766 38273
rect 5710 38093 5766 38149
rect 5710 37969 5766 38025
rect 5710 37845 5766 37901
rect 5710 37721 5766 37777
rect 5710 37597 5766 37653
rect 5710 37473 5766 37529
rect 5710 37349 5766 37405
rect 5710 37225 5766 37281
rect 5710 37101 5766 37157
rect 5710 36977 5766 37033
rect 5710 36853 5766 36909
rect 5834 38106 5890 38162
rect 5834 37982 5890 38038
rect 5834 37858 5890 37914
rect 5834 37734 5890 37790
rect 5834 37610 5890 37666
rect 5834 37486 5890 37542
rect 5834 37362 5890 37418
rect 5834 37238 5890 37294
rect 5834 37114 5890 37170
rect 5834 36990 5890 37046
rect 5834 36866 5890 36922
rect 5958 38085 6014 38141
rect 5958 37961 6014 38017
rect 5958 37837 6014 37893
rect 5958 37713 6014 37769
rect 5958 37589 6014 37645
rect 5958 37465 6014 37521
rect 5958 37341 6014 37397
rect 5958 37217 6014 37273
rect 5958 37093 6014 37149
rect 5958 36969 6014 37025
rect 5958 36845 6014 36901
rect 6082 38084 6138 38140
rect 6082 37960 6138 38016
rect 6082 37836 6138 37892
rect 6082 37712 6138 37768
rect 6082 37588 6138 37644
rect 6082 37464 6138 37520
rect 6082 37340 6138 37396
rect 6082 37216 6138 37272
rect 6082 37092 6138 37148
rect 6082 36968 6138 37024
rect 6082 36844 6138 36900
rect 7562 38088 7618 38144
rect 7686 38088 7742 38144
rect 7810 38088 7866 38144
rect 7934 38088 7990 38144
rect 8058 38088 8114 38144
rect 8182 38088 8238 38144
rect 8306 38088 8362 38144
rect 8430 38088 8486 38144
rect 8554 38088 8610 38144
rect 7562 37964 7618 38020
rect 7686 37964 7742 38020
rect 7810 37964 7866 38020
rect 7934 37964 7990 38020
rect 8058 37964 8114 38020
rect 8182 37964 8238 38020
rect 8306 37964 8362 38020
rect 8430 37964 8486 38020
rect 8554 37964 8610 38020
rect 7562 37840 7618 37896
rect 7686 37840 7742 37896
rect 7810 37840 7866 37896
rect 7934 37840 7990 37896
rect 8058 37840 8114 37896
rect 8182 37840 8238 37896
rect 8306 37840 8362 37896
rect 8430 37840 8486 37896
rect 8554 37840 8610 37896
rect 7562 37716 7618 37772
rect 7686 37716 7742 37772
rect 7810 37716 7866 37772
rect 7934 37716 7990 37772
rect 8058 37716 8114 37772
rect 8182 37716 8238 37772
rect 8306 37716 8362 37772
rect 8430 37716 8486 37772
rect 8554 37716 8610 37772
rect 7562 37592 7618 37648
rect 7686 37592 7742 37648
rect 7810 37592 7866 37648
rect 7934 37592 7990 37648
rect 8058 37592 8114 37648
rect 8182 37592 8238 37648
rect 8306 37592 8362 37648
rect 8430 37592 8486 37648
rect 8554 37592 8610 37648
rect 7562 37468 7618 37524
rect 7686 37468 7742 37524
rect 7810 37468 7866 37524
rect 7934 37468 7990 37524
rect 8058 37468 8114 37524
rect 8182 37468 8238 37524
rect 8306 37468 8362 37524
rect 8430 37468 8486 37524
rect 8554 37468 8610 37524
rect 7562 37344 7618 37400
rect 7686 37344 7742 37400
rect 7810 37344 7866 37400
rect 7934 37344 7990 37400
rect 8058 37344 8114 37400
rect 8182 37344 8238 37400
rect 8306 37344 8362 37400
rect 8430 37344 8486 37400
rect 8554 37344 8610 37400
rect 7562 37220 7618 37276
rect 7686 37220 7742 37276
rect 7810 37220 7866 37276
rect 7934 37220 7990 37276
rect 8058 37220 8114 37276
rect 8182 37220 8238 37276
rect 8306 37220 8362 37276
rect 8430 37220 8486 37276
rect 8554 37220 8610 37276
rect 7562 37096 7618 37152
rect 7686 37096 7742 37152
rect 7810 37096 7866 37152
rect 7934 37096 7990 37152
rect 8058 37096 8114 37152
rect 8182 37096 8238 37152
rect 8306 37096 8362 37152
rect 8430 37096 8486 37152
rect 8554 37096 8610 37152
rect 7562 36972 7618 37028
rect 7686 36972 7742 37028
rect 7810 36972 7866 37028
rect 7934 36972 7990 37028
rect 8058 36972 8114 37028
rect 8182 36972 8238 37028
rect 8306 36972 8362 37028
rect 8430 36972 8486 37028
rect 8554 36972 8610 37028
rect 7562 36848 7618 36904
rect 7686 36848 7742 36904
rect 7810 36848 7866 36904
rect 7934 36848 7990 36904
rect 8058 36848 8114 36904
rect 8182 36848 8238 36904
rect 8306 36848 8362 36904
rect 8430 36848 8486 36904
rect 8554 36848 8610 36904
rect 10679 38088 10735 38144
rect 10803 38088 10859 38144
rect 10927 38088 10983 38144
rect 11051 38088 11107 38144
rect 11175 38088 11231 38144
rect 11299 38088 11355 38144
rect 11423 38088 11479 38144
rect 11547 38088 11603 38144
rect 11671 38088 11727 38144
rect 11795 38088 11851 38144
rect 11919 38088 11975 38144
rect 12043 38088 12099 38144
rect 12167 38088 12223 38144
rect 12291 38088 12347 38144
rect 12415 38088 12471 38144
rect 10679 37964 10735 38020
rect 10803 37964 10859 38020
rect 10927 37964 10983 38020
rect 11051 37964 11107 38020
rect 11175 37964 11231 38020
rect 11299 37964 11355 38020
rect 11423 37964 11479 38020
rect 11547 37964 11603 38020
rect 11671 37964 11727 38020
rect 11795 37964 11851 38020
rect 11919 37964 11975 38020
rect 12043 37964 12099 38020
rect 12167 37964 12223 38020
rect 12291 37964 12347 38020
rect 12415 37964 12471 38020
rect 10679 37840 10735 37896
rect 10803 37840 10859 37896
rect 10927 37840 10983 37896
rect 11051 37840 11107 37896
rect 11175 37840 11231 37896
rect 11299 37840 11355 37896
rect 11423 37840 11479 37896
rect 11547 37840 11603 37896
rect 11671 37840 11727 37896
rect 11795 37840 11851 37896
rect 11919 37840 11975 37896
rect 12043 37840 12099 37896
rect 12167 37840 12223 37896
rect 12291 37840 12347 37896
rect 12415 37840 12471 37896
rect 10679 37716 10735 37772
rect 10803 37716 10859 37772
rect 10927 37716 10983 37772
rect 11051 37716 11107 37772
rect 11175 37716 11231 37772
rect 11299 37716 11355 37772
rect 11423 37716 11479 37772
rect 11547 37716 11603 37772
rect 11671 37716 11727 37772
rect 11795 37716 11851 37772
rect 11919 37716 11975 37772
rect 12043 37716 12099 37772
rect 12167 37716 12223 37772
rect 12291 37716 12347 37772
rect 12415 37716 12471 37772
rect 10679 37592 10735 37648
rect 10803 37592 10859 37648
rect 10927 37592 10983 37648
rect 11051 37592 11107 37648
rect 11175 37592 11231 37648
rect 11299 37592 11355 37648
rect 11423 37592 11479 37648
rect 11547 37592 11603 37648
rect 11671 37592 11727 37648
rect 11795 37592 11851 37648
rect 11919 37592 11975 37648
rect 12043 37592 12099 37648
rect 12167 37592 12223 37648
rect 12291 37592 12347 37648
rect 12415 37592 12471 37648
rect 10679 37468 10735 37524
rect 10803 37468 10859 37524
rect 10927 37468 10983 37524
rect 11051 37468 11107 37524
rect 11175 37468 11231 37524
rect 11299 37468 11355 37524
rect 11423 37468 11479 37524
rect 11547 37468 11603 37524
rect 11671 37468 11727 37524
rect 11795 37468 11851 37524
rect 11919 37468 11975 37524
rect 12043 37468 12099 37524
rect 12167 37468 12223 37524
rect 12291 37468 12347 37524
rect 12415 37468 12471 37524
rect 10679 37344 10735 37400
rect 10803 37344 10859 37400
rect 10927 37344 10983 37400
rect 11051 37344 11107 37400
rect 11175 37344 11231 37400
rect 11299 37344 11355 37400
rect 11423 37344 11479 37400
rect 11547 37344 11603 37400
rect 11671 37344 11727 37400
rect 11795 37344 11851 37400
rect 11919 37344 11975 37400
rect 12043 37344 12099 37400
rect 12167 37344 12223 37400
rect 12291 37344 12347 37400
rect 12415 37344 12471 37400
rect 10679 37220 10735 37276
rect 10803 37220 10859 37276
rect 10927 37220 10983 37276
rect 11051 37220 11107 37276
rect 11175 37220 11231 37276
rect 11299 37220 11355 37276
rect 11423 37220 11479 37276
rect 11547 37220 11603 37276
rect 11671 37220 11727 37276
rect 11795 37220 11851 37276
rect 11919 37220 11975 37276
rect 12043 37220 12099 37276
rect 12167 37220 12223 37276
rect 12291 37220 12347 37276
rect 12415 37220 12471 37276
rect 10679 37096 10735 37152
rect 10803 37096 10859 37152
rect 10927 37096 10983 37152
rect 11051 37096 11107 37152
rect 11175 37096 11231 37152
rect 11299 37096 11355 37152
rect 11423 37096 11479 37152
rect 11547 37096 11603 37152
rect 11671 37096 11727 37152
rect 11795 37096 11851 37152
rect 11919 37096 11975 37152
rect 12043 37096 12099 37152
rect 12167 37096 12223 37152
rect 12291 37096 12347 37152
rect 12415 37096 12471 37152
rect 10679 36972 10735 37028
rect 10803 36972 10859 37028
rect 10927 36972 10983 37028
rect 11051 36972 11107 37028
rect 11175 36972 11231 37028
rect 11299 36972 11355 37028
rect 11423 36972 11479 37028
rect 11547 36972 11603 37028
rect 11671 36972 11727 37028
rect 11795 36972 11851 37028
rect 11919 36972 11975 37028
rect 12043 36972 12099 37028
rect 12167 36972 12223 37028
rect 12291 36972 12347 37028
rect 12415 36972 12471 37028
rect 10679 36848 10735 36904
rect 10803 36848 10859 36904
rect 10927 36848 10983 36904
rect 11051 36848 11107 36904
rect 11175 36848 11231 36904
rect 11299 36848 11355 36904
rect 11423 36848 11479 36904
rect 11547 36848 11603 36904
rect 11671 36848 11727 36904
rect 11795 36848 11851 36904
rect 11919 36848 11975 36904
rect 12043 36848 12099 36904
rect 12167 36848 12223 36904
rect 12291 36848 12347 36904
rect 12415 36848 12471 36904
rect 4139 36669 4195 36725
rect 4139 36545 4195 36601
rect 4139 36421 4195 36477
rect 4139 36297 4195 36353
rect 4139 36173 4195 36229
rect 4139 36049 4195 36105
rect 4139 35925 4195 35981
rect 6368 36488 6424 36544
rect 6492 36488 6548 36544
rect 6616 36488 6672 36544
rect 6740 36488 6796 36544
rect 6864 36488 6920 36544
rect 6988 36488 7044 36544
rect 7112 36488 7168 36544
rect 7236 36488 7292 36544
rect 7360 36488 7416 36544
rect 6368 36364 6424 36420
rect 6492 36364 6548 36420
rect 6616 36364 6672 36420
rect 6740 36364 6796 36420
rect 6864 36364 6920 36420
rect 6988 36364 7044 36420
rect 7112 36364 7168 36420
rect 7236 36364 7292 36420
rect 7360 36364 7416 36420
rect 6368 36240 6424 36296
rect 6492 36240 6548 36296
rect 6616 36240 6672 36296
rect 6740 36240 6796 36296
rect 6864 36240 6920 36296
rect 6988 36240 7044 36296
rect 7112 36240 7168 36296
rect 7236 36240 7292 36296
rect 7360 36240 7416 36296
rect 6368 36116 6424 36172
rect 6492 36116 6548 36172
rect 6616 36116 6672 36172
rect 6740 36116 6796 36172
rect 6864 36116 6920 36172
rect 6988 36116 7044 36172
rect 7112 36116 7168 36172
rect 7236 36116 7292 36172
rect 7360 36116 7416 36172
rect 6368 35992 6424 36048
rect 6492 35992 6548 36048
rect 6616 35992 6672 36048
rect 6740 35992 6796 36048
rect 6864 35992 6920 36048
rect 6988 35992 7044 36048
rect 7112 35992 7168 36048
rect 7236 35992 7292 36048
rect 7360 35992 7416 36048
rect 6368 35868 6424 35924
rect 6492 35868 6548 35924
rect 6616 35868 6672 35924
rect 6740 35868 6796 35924
rect 6864 35868 6920 35924
rect 6988 35868 7044 35924
rect 7112 35868 7168 35924
rect 7236 35868 7292 35924
rect 7360 35868 7416 35924
rect 6368 35744 6424 35800
rect 6492 35744 6548 35800
rect 6616 35744 6672 35800
rect 6740 35744 6796 35800
rect 6864 35744 6920 35800
rect 6988 35744 7044 35800
rect 7112 35744 7168 35800
rect 7236 35744 7292 35800
rect 7360 35744 7416 35800
rect 6368 35620 6424 35676
rect 6492 35620 6548 35676
rect 6616 35620 6672 35676
rect 6740 35620 6796 35676
rect 6864 35620 6920 35676
rect 6988 35620 7044 35676
rect 7112 35620 7168 35676
rect 7236 35620 7292 35676
rect 7360 35620 7416 35676
rect 6368 35496 6424 35552
rect 6492 35496 6548 35552
rect 6616 35496 6672 35552
rect 6740 35496 6796 35552
rect 6864 35496 6920 35552
rect 6988 35496 7044 35552
rect 7112 35496 7168 35552
rect 7236 35496 7292 35552
rect 7360 35496 7416 35552
rect 6368 35372 6424 35428
rect 6492 35372 6548 35428
rect 6616 35372 6672 35428
rect 6740 35372 6796 35428
rect 6864 35372 6920 35428
rect 6988 35372 7044 35428
rect 7112 35372 7168 35428
rect 7236 35372 7292 35428
rect 7360 35372 7416 35428
rect 6368 35248 6424 35304
rect 6492 35248 6548 35304
rect 6616 35248 6672 35304
rect 6740 35248 6796 35304
rect 6864 35248 6920 35304
rect 6988 35248 7044 35304
rect 7112 35248 7168 35304
rect 7236 35248 7292 35304
rect 7360 35248 7416 35304
rect 8751 36488 8807 36544
rect 8875 36488 8931 36544
rect 8999 36488 9055 36544
rect 9123 36488 9179 36544
rect 9247 36488 9303 36544
rect 9371 36488 9427 36544
rect 9495 36488 9551 36544
rect 9619 36488 9675 36544
rect 9743 36488 9799 36544
rect 9867 36488 9923 36544
rect 9991 36488 10047 36544
rect 10115 36488 10171 36544
rect 10239 36488 10295 36544
rect 10363 36488 10419 36544
rect 10487 36488 10543 36544
rect 8751 36364 8807 36420
rect 8875 36364 8931 36420
rect 8999 36364 9055 36420
rect 9123 36364 9179 36420
rect 9247 36364 9303 36420
rect 9371 36364 9427 36420
rect 9495 36364 9551 36420
rect 9619 36364 9675 36420
rect 9743 36364 9799 36420
rect 9867 36364 9923 36420
rect 9991 36364 10047 36420
rect 10115 36364 10171 36420
rect 10239 36364 10295 36420
rect 10363 36364 10419 36420
rect 10487 36364 10543 36420
rect 8751 36240 8807 36296
rect 8875 36240 8931 36296
rect 8999 36240 9055 36296
rect 9123 36240 9179 36296
rect 9247 36240 9303 36296
rect 9371 36240 9427 36296
rect 9495 36240 9551 36296
rect 9619 36240 9675 36296
rect 9743 36240 9799 36296
rect 9867 36240 9923 36296
rect 9991 36240 10047 36296
rect 10115 36240 10171 36296
rect 10239 36240 10295 36296
rect 10363 36240 10419 36296
rect 10487 36240 10543 36296
rect 8751 36116 8807 36172
rect 8875 36116 8931 36172
rect 8999 36116 9055 36172
rect 9123 36116 9179 36172
rect 9247 36116 9303 36172
rect 9371 36116 9427 36172
rect 9495 36116 9551 36172
rect 9619 36116 9675 36172
rect 9743 36116 9799 36172
rect 9867 36116 9923 36172
rect 9991 36116 10047 36172
rect 10115 36116 10171 36172
rect 10239 36116 10295 36172
rect 10363 36116 10419 36172
rect 10487 36116 10543 36172
rect 8751 35992 8807 36048
rect 8875 35992 8931 36048
rect 8999 35992 9055 36048
rect 9123 35992 9179 36048
rect 9247 35992 9303 36048
rect 9371 35992 9427 36048
rect 9495 35992 9551 36048
rect 9619 35992 9675 36048
rect 9743 35992 9799 36048
rect 9867 35992 9923 36048
rect 9991 35992 10047 36048
rect 10115 35992 10171 36048
rect 10239 35992 10295 36048
rect 10363 35992 10419 36048
rect 10487 35992 10543 36048
rect 8751 35868 8807 35924
rect 8875 35868 8931 35924
rect 8999 35868 9055 35924
rect 9123 35868 9179 35924
rect 9247 35868 9303 35924
rect 9371 35868 9427 35924
rect 9495 35868 9551 35924
rect 9619 35868 9675 35924
rect 9743 35868 9799 35924
rect 9867 35868 9923 35924
rect 9991 35868 10047 35924
rect 10115 35868 10171 35924
rect 10239 35868 10295 35924
rect 10363 35868 10419 35924
rect 10487 35868 10543 35924
rect 8751 35744 8807 35800
rect 8875 35744 8931 35800
rect 8999 35744 9055 35800
rect 9123 35744 9179 35800
rect 9247 35744 9303 35800
rect 9371 35744 9427 35800
rect 9495 35744 9551 35800
rect 9619 35744 9675 35800
rect 9743 35744 9799 35800
rect 9867 35744 9923 35800
rect 9991 35744 10047 35800
rect 10115 35744 10171 35800
rect 10239 35744 10295 35800
rect 10363 35744 10419 35800
rect 10487 35744 10543 35800
rect 8751 35620 8807 35676
rect 8875 35620 8931 35676
rect 8999 35620 9055 35676
rect 9123 35620 9179 35676
rect 9247 35620 9303 35676
rect 9371 35620 9427 35676
rect 9495 35620 9551 35676
rect 9619 35620 9675 35676
rect 9743 35620 9799 35676
rect 9867 35620 9923 35676
rect 9991 35620 10047 35676
rect 10115 35620 10171 35676
rect 10239 35620 10295 35676
rect 10363 35620 10419 35676
rect 10487 35620 10543 35676
rect 8751 35496 8807 35552
rect 8875 35496 8931 35552
rect 8999 35496 9055 35552
rect 9123 35496 9179 35552
rect 9247 35496 9303 35552
rect 9371 35496 9427 35552
rect 9495 35496 9551 35552
rect 9619 35496 9675 35552
rect 9743 35496 9799 35552
rect 9867 35496 9923 35552
rect 9991 35496 10047 35552
rect 10115 35496 10171 35552
rect 10239 35496 10295 35552
rect 10363 35496 10419 35552
rect 10487 35496 10543 35552
rect 8751 35372 8807 35428
rect 8875 35372 8931 35428
rect 8999 35372 9055 35428
rect 9123 35372 9179 35428
rect 9247 35372 9303 35428
rect 9371 35372 9427 35428
rect 9495 35372 9551 35428
rect 9619 35372 9675 35428
rect 9743 35372 9799 35428
rect 9867 35372 9923 35428
rect 9991 35372 10047 35428
rect 10115 35372 10171 35428
rect 10239 35372 10295 35428
rect 10363 35372 10419 35428
rect 10487 35372 10543 35428
rect 8751 35248 8807 35304
rect 8875 35248 8931 35304
rect 8999 35248 9055 35304
rect 9123 35248 9179 35304
rect 9247 35248 9303 35304
rect 9371 35248 9427 35304
rect 9495 35248 9551 35304
rect 9619 35248 9675 35304
rect 9743 35248 9799 35304
rect 9867 35248 9923 35304
rect 9991 35248 10047 35304
rect 10115 35248 10171 35304
rect 10239 35248 10295 35304
rect 10363 35248 10419 35304
rect 10487 35248 10543 35304
rect 12852 36488 12908 36544
rect 12976 36488 13032 36544
rect 13100 36488 13156 36544
rect 13224 36488 13280 36544
rect 13348 36488 13404 36544
rect 13472 36488 13528 36544
rect 13596 36488 13652 36544
rect 13720 36488 13776 36544
rect 13844 36488 13900 36544
rect 12852 36364 12908 36420
rect 12976 36364 13032 36420
rect 13100 36364 13156 36420
rect 13224 36364 13280 36420
rect 13348 36364 13404 36420
rect 13472 36364 13528 36420
rect 13596 36364 13652 36420
rect 13720 36364 13776 36420
rect 13844 36364 13900 36420
rect 12852 36240 12908 36296
rect 12976 36240 13032 36296
rect 13100 36240 13156 36296
rect 13224 36240 13280 36296
rect 13348 36240 13404 36296
rect 13472 36240 13528 36296
rect 13596 36240 13652 36296
rect 13720 36240 13776 36296
rect 13844 36240 13900 36296
rect 12852 36116 12908 36172
rect 12976 36116 13032 36172
rect 13100 36116 13156 36172
rect 13224 36116 13280 36172
rect 13348 36116 13404 36172
rect 13472 36116 13528 36172
rect 13596 36116 13652 36172
rect 13720 36116 13776 36172
rect 13844 36116 13900 36172
rect 12852 35992 12908 36048
rect 12976 35992 13032 36048
rect 13100 35992 13156 36048
rect 13224 35992 13280 36048
rect 13348 35992 13404 36048
rect 13472 35992 13528 36048
rect 13596 35992 13652 36048
rect 13720 35992 13776 36048
rect 13844 35992 13900 36048
rect 12852 35868 12908 35924
rect 12976 35868 13032 35924
rect 13100 35868 13156 35924
rect 13224 35868 13280 35924
rect 13348 35868 13404 35924
rect 13472 35868 13528 35924
rect 13596 35868 13652 35924
rect 13720 35868 13776 35924
rect 13844 35868 13900 35924
rect 12852 35744 12908 35800
rect 12976 35744 13032 35800
rect 13100 35744 13156 35800
rect 13224 35744 13280 35800
rect 13348 35744 13404 35800
rect 13472 35744 13528 35800
rect 13596 35744 13652 35800
rect 13720 35744 13776 35800
rect 13844 35744 13900 35800
rect 12852 35620 12908 35676
rect 12976 35620 13032 35676
rect 13100 35620 13156 35676
rect 13224 35620 13280 35676
rect 13348 35620 13404 35676
rect 13472 35620 13528 35676
rect 13596 35620 13652 35676
rect 13720 35620 13776 35676
rect 13844 35620 13900 35676
rect 12852 35496 12908 35552
rect 12976 35496 13032 35552
rect 13100 35496 13156 35552
rect 13224 35496 13280 35552
rect 13348 35496 13404 35552
rect 13472 35496 13528 35552
rect 13596 35496 13652 35552
rect 13720 35496 13776 35552
rect 13844 35496 13900 35552
rect 12852 35372 12908 35428
rect 12976 35372 13032 35428
rect 13100 35372 13156 35428
rect 13224 35372 13280 35428
rect 13348 35372 13404 35428
rect 13472 35372 13528 35428
rect 13596 35372 13652 35428
rect 13720 35372 13776 35428
rect 13844 35372 13900 35428
rect 12852 35248 12908 35304
rect 12976 35248 13032 35304
rect 13100 35248 13156 35304
rect 13224 35248 13280 35304
rect 13348 35248 13404 35304
rect 13472 35248 13528 35304
rect 13596 35248 13652 35304
rect 13720 35248 13776 35304
rect 13844 35248 13900 35304
rect 14767 36570 14823 36572
rect 14767 36518 14769 36570
rect 14769 36518 14821 36570
rect 14821 36518 14823 36570
rect 14767 36462 14823 36518
rect 14767 36410 14769 36462
rect 14769 36410 14821 36462
rect 14821 36410 14823 36462
rect 14767 36354 14823 36410
rect 14767 36302 14769 36354
rect 14769 36302 14821 36354
rect 14821 36302 14823 36354
rect 14767 36246 14823 36302
rect 14767 36194 14769 36246
rect 14769 36194 14821 36246
rect 14821 36194 14823 36246
rect 14767 36138 14823 36194
rect 14767 36086 14769 36138
rect 14769 36086 14821 36138
rect 14821 36086 14823 36138
rect 14767 36030 14823 36086
rect 14767 35978 14769 36030
rect 14769 35978 14821 36030
rect 14821 35978 14823 36030
rect 14767 35922 14823 35978
rect 14767 35870 14769 35922
rect 14769 35870 14821 35922
rect 14821 35870 14823 35922
rect 14767 35814 14823 35870
rect 14767 35762 14769 35814
rect 14769 35762 14821 35814
rect 14821 35762 14823 35814
rect 14767 35706 14823 35762
rect 14767 35654 14769 35706
rect 14769 35654 14821 35706
rect 14821 35654 14823 35706
rect 14767 35598 14823 35654
rect 14767 35546 14769 35598
rect 14769 35546 14821 35598
rect 14821 35546 14823 35598
rect 14767 35490 14823 35546
rect 14767 35438 14769 35490
rect 14769 35438 14821 35490
rect 14821 35438 14823 35490
rect 14767 35382 14823 35438
rect 14767 35330 14769 35382
rect 14769 35330 14821 35382
rect 14821 35330 14823 35382
rect 14767 35274 14823 35330
rect 14767 35222 14769 35274
rect 14769 35222 14821 35274
rect 14821 35222 14823 35274
rect 14767 35220 14823 35222
<< metal3 >>
rect 7640 56433 8460 56443
rect 6182 56422 7002 56432
rect 6182 56366 6192 56422
rect 6248 56366 6316 56422
rect 6372 56366 6440 56422
rect 6496 56366 6564 56422
rect 6620 56366 6688 56422
rect 6744 56366 6812 56422
rect 6868 56366 6936 56422
rect 6992 56366 7002 56422
rect 6182 56298 7002 56366
rect 6182 56242 6192 56298
rect 6248 56242 6316 56298
rect 6372 56242 6440 56298
rect 6496 56242 6564 56298
rect 6620 56242 6688 56298
rect 6744 56242 6812 56298
rect 6868 56242 6936 56298
rect 6992 56242 7002 56298
rect 6182 56174 7002 56242
rect 6182 56118 6192 56174
rect 6248 56118 6316 56174
rect 6372 56118 6440 56174
rect 6496 56118 6564 56174
rect 6620 56118 6688 56174
rect 6744 56118 6812 56174
rect 6868 56118 6936 56174
rect 6992 56118 7002 56174
rect 6182 56050 7002 56118
rect 6182 55994 6192 56050
rect 6248 55994 6316 56050
rect 6372 55994 6440 56050
rect 6496 55994 6564 56050
rect 6620 55994 6688 56050
rect 6744 55994 6812 56050
rect 6868 55994 6936 56050
rect 6992 55994 7002 56050
rect 6182 55926 7002 55994
rect 6182 55870 6192 55926
rect 6248 55870 6316 55926
rect 6372 55870 6440 55926
rect 6496 55870 6564 55926
rect 6620 55870 6688 55926
rect 6744 55870 6812 55926
rect 6868 55870 6936 55926
rect 6992 55870 7002 55926
rect 6182 55802 7002 55870
rect 6182 55746 6192 55802
rect 6248 55746 6316 55802
rect 6372 55746 6440 55802
rect 6496 55746 6564 55802
rect 6620 55746 6688 55802
rect 6744 55746 6812 55802
rect 6868 55746 6936 55802
rect 6992 55746 7002 55802
rect 6182 55678 7002 55746
rect 6182 55622 6192 55678
rect 6248 55622 6316 55678
rect 6372 55622 6440 55678
rect 6496 55622 6564 55678
rect 6620 55622 6688 55678
rect 6744 55622 6812 55678
rect 6868 55622 6936 55678
rect 6992 55622 7002 55678
rect 6182 55554 7002 55622
rect 6182 55498 6192 55554
rect 6248 55498 6316 55554
rect 6372 55498 6440 55554
rect 6496 55498 6564 55554
rect 6620 55498 6688 55554
rect 6744 55498 6812 55554
rect 6868 55498 6936 55554
rect 6992 55498 7002 55554
rect 6182 55430 7002 55498
rect 6182 55374 6192 55430
rect 6248 55374 6316 55430
rect 6372 55374 6440 55430
rect 6496 55374 6564 55430
rect 6620 55374 6688 55430
rect 6744 55374 6812 55430
rect 6868 55374 6936 55430
rect 6992 55374 7002 55430
rect 6182 55306 7002 55374
rect 6182 55250 6192 55306
rect 6248 55250 6316 55306
rect 6372 55250 6440 55306
rect 6496 55250 6564 55306
rect 6620 55250 6688 55306
rect 6744 55250 6812 55306
rect 6868 55250 6936 55306
rect 6992 55250 7002 55306
rect 6182 55182 7002 55250
rect 6182 55126 6192 55182
rect 6248 55126 6316 55182
rect 6372 55126 6440 55182
rect 6496 55126 6564 55182
rect 6620 55126 6688 55182
rect 6744 55126 6812 55182
rect 6868 55126 6936 55182
rect 6992 55126 7002 55182
rect 6182 55058 7002 55126
rect 6182 55002 6192 55058
rect 6248 55002 6316 55058
rect 6372 55002 6440 55058
rect 6496 55002 6564 55058
rect 6620 55002 6688 55058
rect 6744 55002 6812 55058
rect 6868 55002 6936 55058
rect 6992 55002 7002 55058
rect 6182 54934 7002 55002
rect 6182 54878 6192 54934
rect 6248 54878 6316 54934
rect 6372 54878 6440 54934
rect 6496 54878 6564 54934
rect 6620 54878 6688 54934
rect 6744 54878 6812 54934
rect 6868 54878 6936 54934
rect 6992 54878 7002 54934
rect 6182 54810 7002 54878
rect 6182 54754 6192 54810
rect 6248 54754 6316 54810
rect 6372 54754 6440 54810
rect 6496 54754 6564 54810
rect 6620 54754 6688 54810
rect 6744 54754 6812 54810
rect 6868 54754 6936 54810
rect 6992 54754 7002 54810
rect 6182 54686 7002 54754
rect 6182 54630 6192 54686
rect 6248 54630 6316 54686
rect 6372 54630 6440 54686
rect 6496 54630 6564 54686
rect 6620 54630 6688 54686
rect 6744 54630 6812 54686
rect 6868 54630 6936 54686
rect 6992 54630 7002 54686
rect 6182 54562 7002 54630
rect 6182 54506 6192 54562
rect 6248 54506 6316 54562
rect 6372 54506 6440 54562
rect 6496 54506 6564 54562
rect 6620 54506 6688 54562
rect 6744 54506 6812 54562
rect 6868 54506 6936 54562
rect 6992 54506 7002 54562
rect 6182 54438 7002 54506
rect 6182 54382 6192 54438
rect 6248 54382 6316 54438
rect 6372 54382 6440 54438
rect 6496 54382 6564 54438
rect 6620 54382 6688 54438
rect 6744 54382 6812 54438
rect 6868 54382 6936 54438
rect 6992 54382 7002 54438
rect 6182 54314 7002 54382
rect 6182 54258 6192 54314
rect 6248 54258 6316 54314
rect 6372 54258 6440 54314
rect 6496 54258 6564 54314
rect 6620 54258 6688 54314
rect 6744 54258 6812 54314
rect 6868 54258 6936 54314
rect 6992 54258 7002 54314
rect 6182 54190 7002 54258
rect 6182 54134 6192 54190
rect 6248 54134 6316 54190
rect 6372 54134 6440 54190
rect 6496 54134 6564 54190
rect 6620 54134 6688 54190
rect 6744 54134 6812 54190
rect 6868 54134 6936 54190
rect 6992 54134 7002 54190
rect 6182 54066 7002 54134
rect 6182 54010 6192 54066
rect 6248 54010 6316 54066
rect 6372 54010 6440 54066
rect 6496 54010 6564 54066
rect 6620 54010 6688 54066
rect 6744 54010 6812 54066
rect 6868 54010 6936 54066
rect 6992 54010 7002 54066
rect 6182 53942 7002 54010
rect 6182 53886 6192 53942
rect 6248 53886 6316 53942
rect 6372 53886 6440 53942
rect 6496 53886 6564 53942
rect 6620 53886 6688 53942
rect 6744 53886 6812 53942
rect 6868 53886 6936 53942
rect 6992 53886 7002 53942
rect 6182 53818 7002 53886
rect 6182 53762 6192 53818
rect 6248 53762 6316 53818
rect 6372 53762 6440 53818
rect 6496 53762 6564 53818
rect 6620 53762 6688 53818
rect 6744 53762 6812 53818
rect 6868 53762 6936 53818
rect 6992 53762 7002 53818
rect 6182 53694 7002 53762
rect 6182 53638 6192 53694
rect 6248 53638 6316 53694
rect 6372 53638 6440 53694
rect 6496 53638 6564 53694
rect 6620 53638 6688 53694
rect 6744 53638 6812 53694
rect 6868 53638 6936 53694
rect 6992 53638 7002 53694
rect 6182 53570 7002 53638
rect 6182 53514 6192 53570
rect 6248 53514 6316 53570
rect 6372 53514 6440 53570
rect 6496 53514 6564 53570
rect 6620 53514 6688 53570
rect 6744 53514 6812 53570
rect 6868 53514 6936 53570
rect 6992 53514 7002 53570
rect 6182 53446 7002 53514
rect 6182 53390 6192 53446
rect 6248 53390 6316 53446
rect 6372 53390 6440 53446
rect 6496 53390 6564 53446
rect 6620 53390 6688 53446
rect 6744 53390 6812 53446
rect 6868 53390 6936 53446
rect 6992 53390 7002 53446
rect 6182 53322 7002 53390
rect 6182 53266 6192 53322
rect 6248 53266 6316 53322
rect 6372 53266 6440 53322
rect 6496 53266 6564 53322
rect 6620 53266 6688 53322
rect 6744 53266 6812 53322
rect 6868 53266 6936 53322
rect 6992 53266 7002 53322
rect 6182 53256 7002 53266
rect 7640 56377 7650 56433
rect 7706 56377 7774 56433
rect 7830 56377 7898 56433
rect 7954 56377 8022 56433
rect 8078 56377 8146 56433
rect 8202 56377 8270 56433
rect 8326 56377 8394 56433
rect 8450 56377 8460 56433
rect 7640 56309 8460 56377
rect 7640 56253 7650 56309
rect 7706 56253 7774 56309
rect 7830 56253 7898 56309
rect 7954 56253 8022 56309
rect 8078 56253 8146 56309
rect 8202 56253 8270 56309
rect 8326 56253 8394 56309
rect 8450 56253 8460 56309
rect 7640 56185 8460 56253
rect 7640 56129 7650 56185
rect 7706 56129 7774 56185
rect 7830 56129 7898 56185
rect 7954 56129 8022 56185
rect 8078 56129 8146 56185
rect 8202 56129 8270 56185
rect 8326 56129 8394 56185
rect 8450 56129 8460 56185
rect 7640 56061 8460 56129
rect 7640 56005 7650 56061
rect 7706 56005 7774 56061
rect 7830 56005 7898 56061
rect 7954 56005 8022 56061
rect 8078 56005 8146 56061
rect 8202 56005 8270 56061
rect 8326 56005 8394 56061
rect 8450 56005 8460 56061
rect 7640 55937 8460 56005
rect 7640 55881 7650 55937
rect 7706 55881 7774 55937
rect 7830 55881 7898 55937
rect 7954 55881 8022 55937
rect 8078 55881 8146 55937
rect 8202 55881 8270 55937
rect 8326 55881 8394 55937
rect 8450 55881 8460 55937
rect 7640 55813 8460 55881
rect 7640 55757 7650 55813
rect 7706 55757 7774 55813
rect 7830 55757 7898 55813
rect 7954 55757 8022 55813
rect 8078 55757 8146 55813
rect 8202 55757 8270 55813
rect 8326 55757 8394 55813
rect 8450 55757 8460 55813
rect 7640 55689 8460 55757
rect 7640 55633 7650 55689
rect 7706 55633 7774 55689
rect 7830 55633 7898 55689
rect 7954 55633 8022 55689
rect 8078 55633 8146 55689
rect 8202 55633 8270 55689
rect 8326 55633 8394 55689
rect 8450 55633 8460 55689
rect 7640 55565 8460 55633
rect 7640 55509 7650 55565
rect 7706 55509 7774 55565
rect 7830 55509 7898 55565
rect 7954 55509 8022 55565
rect 8078 55509 8146 55565
rect 8202 55509 8270 55565
rect 8326 55509 8394 55565
rect 8450 55509 8460 55565
rect 7640 55441 8460 55509
rect 7640 55385 7650 55441
rect 7706 55385 7774 55441
rect 7830 55385 7898 55441
rect 7954 55385 8022 55441
rect 8078 55385 8146 55441
rect 8202 55385 8270 55441
rect 8326 55385 8394 55441
rect 8450 55385 8460 55441
rect 7640 55317 8460 55385
rect 7640 55261 7650 55317
rect 7706 55261 7774 55317
rect 7830 55261 7898 55317
rect 7954 55261 8022 55317
rect 8078 55261 8146 55317
rect 8202 55261 8270 55317
rect 8326 55261 8394 55317
rect 8450 55261 8460 55317
rect 7640 55193 8460 55261
rect 7640 55137 7650 55193
rect 7706 55137 7774 55193
rect 7830 55137 7898 55193
rect 7954 55137 8022 55193
rect 8078 55137 8146 55193
rect 8202 55137 8270 55193
rect 8326 55137 8394 55193
rect 8450 55137 8460 55193
rect 7640 55069 8460 55137
rect 7640 55013 7650 55069
rect 7706 55013 7774 55069
rect 7830 55013 7898 55069
rect 7954 55013 8022 55069
rect 8078 55013 8146 55069
rect 8202 55013 8270 55069
rect 8326 55013 8394 55069
rect 8450 55013 8460 55069
rect 7640 54945 8460 55013
rect 7640 54889 7650 54945
rect 7706 54889 7774 54945
rect 7830 54889 7898 54945
rect 7954 54889 8022 54945
rect 8078 54889 8146 54945
rect 8202 54889 8270 54945
rect 8326 54889 8394 54945
rect 8450 54889 8460 54945
rect 7640 54821 8460 54889
rect 7640 54765 7650 54821
rect 7706 54765 7774 54821
rect 7830 54765 7898 54821
rect 7954 54765 8022 54821
rect 8078 54765 8146 54821
rect 8202 54765 8270 54821
rect 8326 54765 8394 54821
rect 8450 54765 8460 54821
rect 7640 54697 8460 54765
rect 7640 54641 7650 54697
rect 7706 54641 7774 54697
rect 7830 54641 7898 54697
rect 7954 54641 8022 54697
rect 8078 54641 8146 54697
rect 8202 54641 8270 54697
rect 8326 54641 8394 54697
rect 8450 54641 8460 54697
rect 7640 54573 8460 54641
rect 7640 54517 7650 54573
rect 7706 54517 7774 54573
rect 7830 54517 7898 54573
rect 7954 54517 8022 54573
rect 8078 54517 8146 54573
rect 8202 54517 8270 54573
rect 8326 54517 8394 54573
rect 8450 54517 8460 54573
rect 7640 54449 8460 54517
rect 7640 54393 7650 54449
rect 7706 54393 7774 54449
rect 7830 54393 7898 54449
rect 7954 54393 8022 54449
rect 8078 54393 8146 54449
rect 8202 54393 8270 54449
rect 8326 54393 8394 54449
rect 8450 54393 8460 54449
rect 7640 54325 8460 54393
rect 7640 54269 7650 54325
rect 7706 54269 7774 54325
rect 7830 54269 7898 54325
rect 7954 54269 8022 54325
rect 8078 54269 8146 54325
rect 8202 54269 8270 54325
rect 8326 54269 8394 54325
rect 8450 54269 8460 54325
rect 7640 54201 8460 54269
rect 7640 54145 7650 54201
rect 7706 54145 7774 54201
rect 7830 54145 7898 54201
rect 7954 54145 8022 54201
rect 8078 54145 8146 54201
rect 8202 54145 8270 54201
rect 8326 54145 8394 54201
rect 8450 54145 8460 54201
rect 7640 54077 8460 54145
rect 7640 54021 7650 54077
rect 7706 54021 7774 54077
rect 7830 54021 7898 54077
rect 7954 54021 8022 54077
rect 8078 54021 8146 54077
rect 8202 54021 8270 54077
rect 8326 54021 8394 54077
rect 8450 54021 8460 54077
rect 7640 53953 8460 54021
rect 7640 53897 7650 53953
rect 7706 53897 7774 53953
rect 7830 53897 7898 53953
rect 7954 53897 8022 53953
rect 8078 53897 8146 53953
rect 8202 53897 8270 53953
rect 8326 53897 8394 53953
rect 8450 53897 8460 53953
rect 7640 53829 8460 53897
rect 7640 53773 7650 53829
rect 7706 53773 7774 53829
rect 7830 53773 7898 53829
rect 7954 53773 8022 53829
rect 8078 53773 8146 53829
rect 8202 53773 8270 53829
rect 8326 53773 8394 53829
rect 8450 53773 8460 53829
rect 7640 53705 8460 53773
rect 7640 53649 7650 53705
rect 7706 53649 7774 53705
rect 7830 53649 7898 53705
rect 7954 53649 8022 53705
rect 8078 53649 8146 53705
rect 8202 53649 8270 53705
rect 8326 53649 8394 53705
rect 8450 53649 8460 53705
rect 7640 53581 8460 53649
rect 7640 53525 7650 53581
rect 7706 53525 7774 53581
rect 7830 53525 7898 53581
rect 7954 53525 8022 53581
rect 8078 53525 8146 53581
rect 8202 53525 8270 53581
rect 8326 53525 8394 53581
rect 8450 53525 8460 53581
rect 7640 53457 8460 53525
rect 7640 53401 7650 53457
rect 7706 53401 7774 53457
rect 7830 53401 7898 53457
rect 7954 53401 8022 53457
rect 8078 53401 8146 53457
rect 8202 53401 8270 53457
rect 8326 53401 8394 53457
rect 8450 53401 8460 53457
rect 7640 53333 8460 53401
rect 7640 53277 7650 53333
rect 7706 53277 7774 53333
rect 7830 53277 7898 53333
rect 7954 53277 8022 53333
rect 8078 53277 8146 53333
rect 8202 53277 8270 53333
rect 8326 53277 8394 53333
rect 8450 53277 8460 53333
rect 7640 53209 8460 53277
rect 7640 53153 7650 53209
rect 7706 53153 7774 53209
rect 7830 53153 7898 53209
rect 7954 53153 8022 53209
rect 8078 53153 8146 53209
rect 8202 53153 8270 53209
rect 8326 53153 8394 53209
rect 8450 53153 8460 53209
rect 7640 53085 8460 53153
rect 7640 53029 7650 53085
rect 7706 53029 7774 53085
rect 7830 53029 7898 53085
rect 7954 53029 8022 53085
rect 8078 53029 8146 53085
rect 8202 53029 8270 53085
rect 8326 53029 8394 53085
rect 8450 53029 8460 53085
rect 7640 52961 8460 53029
rect 7640 52905 7650 52961
rect 7706 52905 7774 52961
rect 7830 52905 7898 52961
rect 7954 52905 8022 52961
rect 8078 52905 8146 52961
rect 8202 52905 8270 52961
rect 8326 52905 8394 52961
rect 8450 52905 8460 52961
rect 7640 52837 8460 52905
rect 7640 52781 7650 52837
rect 7706 52781 7774 52837
rect 7830 52781 7898 52837
rect 7954 52781 8022 52837
rect 8078 52781 8146 52837
rect 8202 52781 8270 52837
rect 8326 52781 8394 52837
rect 8450 52781 8460 52837
rect 7640 52771 8460 52781
rect 8802 52737 9498 52747
rect 8802 52681 8812 52737
rect 8868 52681 8936 52737
rect 8992 52681 9060 52737
rect 9116 52681 9184 52737
rect 9240 52681 9308 52737
rect 9364 52681 9432 52737
rect 9488 52681 9498 52737
rect 8802 52613 9498 52681
rect 8802 52557 8812 52613
rect 8868 52557 8936 52613
rect 8992 52557 9060 52613
rect 9116 52557 9184 52613
rect 9240 52557 9308 52613
rect 9364 52557 9432 52613
rect 9488 52557 9498 52613
rect 8802 52489 9498 52557
rect 8802 52433 8812 52489
rect 8868 52433 8936 52489
rect 8992 52433 9060 52489
rect 9116 52433 9184 52489
rect 9240 52433 9308 52489
rect 9364 52433 9432 52489
rect 9488 52433 9498 52489
rect 8802 52365 9498 52433
rect 8802 52309 8812 52365
rect 8868 52309 8936 52365
rect 8992 52309 9060 52365
rect 9116 52309 9184 52365
rect 9240 52309 9308 52365
rect 9364 52309 9432 52365
rect 9488 52309 9498 52365
rect 8802 52241 9498 52309
rect 8802 52185 8812 52241
rect 8868 52185 8936 52241
rect 8992 52185 9060 52241
rect 9116 52185 9184 52241
rect 9240 52185 9308 52241
rect 9364 52185 9432 52241
rect 9488 52185 9498 52241
rect 8802 52117 9498 52185
rect 8802 52061 8812 52117
rect 8868 52061 8936 52117
rect 8992 52061 9060 52117
rect 9116 52061 9184 52117
rect 9240 52061 9308 52117
rect 9364 52061 9432 52117
rect 9488 52061 9498 52117
rect 8802 51993 9498 52061
rect 8802 51937 8812 51993
rect 8868 51937 8936 51993
rect 8992 51937 9060 51993
rect 9116 51937 9184 51993
rect 9240 51937 9308 51993
rect 9364 51937 9432 51993
rect 9488 51937 9498 51993
rect 8802 51869 9498 51937
rect 8802 51813 8812 51869
rect 8868 51813 8936 51869
rect 8992 51813 9060 51869
rect 9116 51813 9184 51869
rect 9240 51813 9308 51869
rect 9364 51813 9432 51869
rect 9488 51813 9498 51869
rect 8802 51745 9498 51813
rect 8802 51689 8812 51745
rect 8868 51689 8936 51745
rect 8992 51689 9060 51745
rect 9116 51689 9184 51745
rect 9240 51689 9308 51745
rect 9364 51689 9432 51745
rect 9488 51689 9498 51745
rect 8802 51621 9498 51689
rect 8802 51565 8812 51621
rect 8868 51565 8936 51621
rect 8992 51565 9060 51621
rect 9116 51565 9184 51621
rect 9240 51565 9308 51621
rect 9364 51565 9432 51621
rect 9488 51565 9498 51621
rect 8802 51555 9498 51565
rect 7640 51452 8460 51462
rect 7640 51396 7650 51452
rect 7706 51396 7774 51452
rect 7830 51396 7898 51452
rect 7954 51396 8022 51452
rect 8078 51396 8146 51452
rect 8202 51396 8270 51452
rect 8326 51396 8394 51452
rect 8450 51396 8460 51452
rect 7640 51328 8460 51396
rect 7640 51272 7650 51328
rect 7706 51272 7774 51328
rect 7830 51272 7898 51328
rect 7954 51272 8022 51328
rect 8078 51272 8146 51328
rect 8202 51272 8270 51328
rect 8326 51272 8394 51328
rect 8450 51272 8460 51328
rect 7640 51204 8460 51272
rect 7640 51148 7650 51204
rect 7706 51148 7774 51204
rect 7830 51148 7898 51204
rect 7954 51148 8022 51204
rect 8078 51148 8146 51204
rect 8202 51148 8270 51204
rect 8326 51148 8394 51204
rect 8450 51148 8460 51204
rect 7640 51080 8460 51148
rect 7640 51024 7650 51080
rect 7706 51024 7774 51080
rect 7830 51024 7898 51080
rect 7954 51024 8022 51080
rect 8078 51024 8146 51080
rect 8202 51024 8270 51080
rect 8326 51024 8394 51080
rect 8450 51024 8460 51080
rect 7640 50956 8460 51024
rect 7640 50900 7650 50956
rect 7706 50900 7774 50956
rect 7830 50900 7898 50956
rect 7954 50900 8022 50956
rect 8078 50900 8146 50956
rect 8202 50900 8270 50956
rect 8326 50900 8394 50956
rect 8450 50900 8460 50956
rect 14757 50972 14833 50982
rect 7640 50832 8460 50900
rect 7640 50776 7650 50832
rect 7706 50776 7774 50832
rect 7830 50776 7898 50832
rect 7954 50776 8022 50832
rect 8078 50776 8146 50832
rect 8202 50776 8270 50832
rect 8326 50776 8394 50832
rect 8450 50776 8460 50832
rect 7640 50708 8460 50776
rect 7640 50652 7650 50708
rect 7706 50652 7774 50708
rect 7830 50652 7898 50708
rect 7954 50652 8022 50708
rect 8078 50652 8146 50708
rect 8202 50652 8270 50708
rect 8326 50652 8394 50708
rect 8450 50652 8460 50708
rect 7640 50584 8460 50652
rect 7640 50528 7650 50584
rect 7706 50528 7774 50584
rect 7830 50528 7898 50584
rect 7954 50528 8022 50584
rect 8078 50528 8146 50584
rect 8202 50528 8270 50584
rect 8326 50528 8394 50584
rect 8450 50528 8460 50584
rect 7640 50518 8460 50528
rect 12842 50938 13910 50948
rect 12842 50882 12852 50938
rect 12908 50882 12976 50938
rect 13032 50882 13100 50938
rect 13156 50882 13224 50938
rect 13280 50882 13348 50938
rect 13404 50882 13472 50938
rect 13528 50882 13596 50938
rect 13652 50882 13720 50938
rect 13776 50882 13844 50938
rect 13900 50882 13910 50938
rect 12842 50814 13910 50882
rect 12842 50758 12852 50814
rect 12908 50758 12976 50814
rect 13032 50758 13100 50814
rect 13156 50758 13224 50814
rect 13280 50758 13348 50814
rect 13404 50758 13472 50814
rect 13528 50758 13596 50814
rect 13652 50758 13720 50814
rect 13776 50758 13844 50814
rect 13900 50758 13910 50814
rect 12842 50690 13910 50758
rect 12842 50634 12852 50690
rect 12908 50634 12976 50690
rect 13032 50634 13100 50690
rect 13156 50634 13224 50690
rect 13280 50634 13348 50690
rect 13404 50634 13472 50690
rect 13528 50634 13596 50690
rect 13652 50634 13720 50690
rect 13776 50634 13844 50690
rect 13900 50634 13910 50690
rect 12842 50566 13910 50634
rect 12842 50510 12852 50566
rect 12908 50510 12976 50566
rect 13032 50510 13100 50566
rect 13156 50510 13224 50566
rect 13280 50510 13348 50566
rect 13404 50510 13472 50566
rect 13528 50510 13596 50566
rect 13652 50510 13720 50566
rect 13776 50510 13844 50566
rect 13900 50510 13910 50566
rect 12842 50442 13910 50510
rect 12842 50386 12852 50442
rect 12908 50386 12976 50442
rect 13032 50386 13100 50442
rect 13156 50386 13224 50442
rect 13280 50386 13348 50442
rect 13404 50386 13472 50442
rect 13528 50386 13596 50442
rect 13652 50386 13720 50442
rect 13776 50386 13844 50442
rect 13900 50386 13910 50442
rect 12842 50318 13910 50386
rect 12842 50262 12852 50318
rect 12908 50262 12976 50318
rect 13032 50262 13100 50318
rect 13156 50262 13224 50318
rect 13280 50262 13348 50318
rect 13404 50262 13472 50318
rect 13528 50262 13596 50318
rect 13652 50262 13720 50318
rect 13776 50262 13844 50318
rect 13900 50262 13910 50318
rect 12842 50194 13910 50262
rect 12842 50138 12852 50194
rect 12908 50138 12976 50194
rect 13032 50138 13100 50194
rect 13156 50138 13224 50194
rect 13280 50138 13348 50194
rect 13404 50138 13472 50194
rect 13528 50138 13596 50194
rect 13652 50138 13720 50194
rect 13776 50138 13844 50194
rect 13900 50138 13910 50194
rect 12842 50070 13910 50138
rect 12842 50014 12852 50070
rect 12908 50014 12976 50070
rect 13032 50014 13100 50070
rect 13156 50014 13224 50070
rect 13280 50014 13348 50070
rect 13404 50014 13472 50070
rect 13528 50014 13596 50070
rect 13652 50014 13720 50070
rect 13776 50014 13844 50070
rect 13900 50014 13910 50070
rect 12842 49946 13910 50014
rect 12842 49890 12852 49946
rect 12908 49890 12976 49946
rect 13032 49890 13100 49946
rect 13156 49890 13224 49946
rect 13280 49890 13348 49946
rect 13404 49890 13472 49946
rect 13528 49890 13596 49946
rect 13652 49890 13720 49946
rect 13776 49890 13844 49946
rect 13900 49890 13910 49946
rect 12842 49822 13910 49890
rect 12842 49766 12852 49822
rect 12908 49766 12976 49822
rect 13032 49766 13100 49822
rect 13156 49766 13224 49822
rect 13280 49766 13348 49822
rect 13404 49766 13472 49822
rect 13528 49766 13596 49822
rect 13652 49766 13720 49822
rect 13776 49766 13844 49822
rect 13900 49766 13910 49822
rect 12842 49698 13910 49766
rect 12842 49642 12852 49698
rect 12908 49642 12976 49698
rect 13032 49642 13100 49698
rect 13156 49642 13224 49698
rect 13280 49642 13348 49698
rect 13404 49642 13472 49698
rect 13528 49642 13596 49698
rect 13652 49642 13720 49698
rect 13776 49642 13844 49698
rect 13900 49642 13910 49698
rect 12842 49632 13910 49642
rect 14757 49620 14767 50972
rect 14823 49620 14833 50972
rect 14757 49610 14833 49620
rect 10669 49346 12481 49356
rect 10669 49290 10679 49346
rect 10735 49290 10803 49346
rect 10859 49290 10927 49346
rect 10983 49290 11051 49346
rect 11107 49290 11175 49346
rect 11231 49290 11299 49346
rect 11355 49290 11423 49346
rect 11479 49290 11547 49346
rect 11603 49290 11671 49346
rect 11727 49290 11795 49346
rect 11851 49290 11919 49346
rect 11975 49290 12043 49346
rect 12099 49290 12167 49346
rect 12223 49290 12291 49346
rect 12347 49290 12415 49346
rect 12471 49290 12481 49346
rect 10669 49222 12481 49290
rect 10669 49166 10679 49222
rect 10735 49166 10803 49222
rect 10859 49166 10927 49222
rect 10983 49166 11051 49222
rect 11107 49166 11175 49222
rect 11231 49166 11299 49222
rect 11355 49166 11423 49222
rect 11479 49166 11547 49222
rect 11603 49166 11671 49222
rect 11727 49166 11795 49222
rect 11851 49166 11919 49222
rect 11975 49166 12043 49222
rect 12099 49166 12167 49222
rect 12223 49166 12291 49222
rect 12347 49166 12415 49222
rect 12471 49166 12481 49222
rect 10669 49098 12481 49166
rect 10669 49042 10679 49098
rect 10735 49042 10803 49098
rect 10859 49042 10927 49098
rect 10983 49042 11051 49098
rect 11107 49042 11175 49098
rect 11231 49042 11299 49098
rect 11355 49042 11423 49098
rect 11479 49042 11547 49098
rect 11603 49042 11671 49098
rect 11727 49042 11795 49098
rect 11851 49042 11919 49098
rect 11975 49042 12043 49098
rect 12099 49042 12167 49098
rect 12223 49042 12291 49098
rect 12347 49042 12415 49098
rect 12471 49042 12481 49098
rect 10669 48974 12481 49042
rect 10669 48918 10679 48974
rect 10735 48918 10803 48974
rect 10859 48918 10927 48974
rect 10983 48918 11051 48974
rect 11107 48918 11175 48974
rect 11231 48918 11299 48974
rect 11355 48918 11423 48974
rect 11479 48918 11547 48974
rect 11603 48918 11671 48974
rect 11727 48918 11795 48974
rect 11851 48918 11919 48974
rect 11975 48918 12043 48974
rect 12099 48918 12167 48974
rect 12223 48918 12291 48974
rect 12347 48918 12415 48974
rect 12471 48918 12481 48974
rect 10669 48850 12481 48918
rect 10669 48794 10679 48850
rect 10735 48794 10803 48850
rect 10859 48794 10927 48850
rect 10983 48794 11051 48850
rect 11107 48794 11175 48850
rect 11231 48794 11299 48850
rect 11355 48794 11423 48850
rect 11479 48794 11547 48850
rect 11603 48794 11671 48850
rect 11727 48794 11795 48850
rect 11851 48794 11919 48850
rect 11975 48794 12043 48850
rect 12099 48794 12167 48850
rect 12223 48794 12291 48850
rect 12347 48794 12415 48850
rect 12471 48794 12481 48850
rect 10669 48726 12481 48794
rect 10669 48670 10679 48726
rect 10735 48670 10803 48726
rect 10859 48670 10927 48726
rect 10983 48670 11051 48726
rect 11107 48670 11175 48726
rect 11231 48670 11299 48726
rect 11355 48670 11423 48726
rect 11479 48670 11547 48726
rect 11603 48670 11671 48726
rect 11727 48670 11795 48726
rect 11851 48670 11919 48726
rect 11975 48670 12043 48726
rect 12099 48670 12167 48726
rect 12223 48670 12291 48726
rect 12347 48670 12415 48726
rect 12471 48670 12481 48726
rect 10669 48602 12481 48670
rect 10669 48546 10679 48602
rect 10735 48546 10803 48602
rect 10859 48546 10927 48602
rect 10983 48546 11051 48602
rect 11107 48546 11175 48602
rect 11231 48546 11299 48602
rect 11355 48546 11423 48602
rect 11479 48546 11547 48602
rect 11603 48546 11671 48602
rect 11727 48546 11795 48602
rect 11851 48546 11919 48602
rect 11975 48546 12043 48602
rect 12099 48546 12167 48602
rect 12223 48546 12291 48602
rect 12347 48546 12415 48602
rect 12471 48546 12481 48602
rect 10669 48478 12481 48546
rect 10669 48422 10679 48478
rect 10735 48422 10803 48478
rect 10859 48422 10927 48478
rect 10983 48422 11051 48478
rect 11107 48422 11175 48478
rect 11231 48422 11299 48478
rect 11355 48422 11423 48478
rect 11479 48422 11547 48478
rect 11603 48422 11671 48478
rect 11727 48422 11795 48478
rect 11851 48422 11919 48478
rect 11975 48422 12043 48478
rect 12099 48422 12167 48478
rect 12223 48422 12291 48478
rect 12347 48422 12415 48478
rect 12471 48422 12481 48478
rect 10669 48354 12481 48422
rect 10669 48298 10679 48354
rect 10735 48298 10803 48354
rect 10859 48298 10927 48354
rect 10983 48298 11051 48354
rect 11107 48298 11175 48354
rect 11231 48298 11299 48354
rect 11355 48298 11423 48354
rect 11479 48298 11547 48354
rect 11603 48298 11671 48354
rect 11727 48298 11795 48354
rect 11851 48298 11919 48354
rect 11975 48298 12043 48354
rect 12099 48298 12167 48354
rect 12223 48298 12291 48354
rect 12347 48298 12415 48354
rect 12471 48298 12481 48354
rect 10669 48230 12481 48298
rect 10669 48174 10679 48230
rect 10735 48174 10803 48230
rect 10859 48174 10927 48230
rect 10983 48174 11051 48230
rect 11107 48174 11175 48230
rect 11231 48174 11299 48230
rect 11355 48174 11423 48230
rect 11479 48174 11547 48230
rect 11603 48174 11671 48230
rect 11727 48174 11795 48230
rect 11851 48174 11919 48230
rect 11975 48174 12043 48230
rect 12099 48174 12167 48230
rect 12223 48174 12291 48230
rect 12347 48174 12415 48230
rect 12471 48174 12481 48230
rect 10669 48106 12481 48174
rect 10669 48050 10679 48106
rect 10735 48050 10803 48106
rect 10859 48050 10927 48106
rect 10983 48050 11051 48106
rect 11107 48050 11175 48106
rect 11231 48050 11299 48106
rect 11355 48050 11423 48106
rect 11479 48050 11547 48106
rect 11603 48050 11671 48106
rect 11727 48050 11795 48106
rect 11851 48050 11919 48106
rect 11975 48050 12043 48106
rect 12099 48050 12167 48106
rect 12223 48050 12291 48106
rect 12347 48050 12415 48106
rect 12471 48050 12481 48106
rect 10669 48040 12481 48050
rect 1094 42890 1170 42900
rect 1094 42834 1104 42890
rect 1160 42834 1170 42890
rect 1094 42766 1170 42834
rect 1094 42710 1104 42766
rect 1160 42710 1170 42766
rect 1094 42642 1170 42710
rect 1094 42586 1104 42642
rect 1160 42586 1170 42642
rect 1094 42518 1170 42586
rect 1094 42462 1104 42518
rect 1160 42462 1170 42518
rect 1094 42394 1170 42462
rect 1094 42338 1104 42394
rect 1160 42338 1170 42394
rect 1094 42270 1170 42338
rect 1094 42214 1104 42270
rect 1160 42214 1170 42270
rect 1094 42146 1170 42214
rect 1094 42090 1104 42146
rect 1160 42090 1170 42146
rect 1094 42022 1170 42090
rect 1094 41966 1104 42022
rect 1160 41966 1170 42022
rect 1094 41898 1170 41966
rect 1094 41842 1104 41898
rect 1160 41842 1170 41898
rect 1094 41774 1170 41842
rect 1094 41718 1104 41774
rect 1160 41718 1170 41774
rect 1094 41650 1170 41718
rect 1094 41594 1104 41650
rect 1160 41594 1170 41650
rect 1094 41526 1170 41594
rect 1094 41470 1104 41526
rect 1160 41470 1170 41526
rect 1094 41402 1170 41470
rect 1094 41346 1104 41402
rect 1160 41346 1170 41402
rect 1094 41278 1170 41346
rect 1094 41222 1104 41278
rect 1160 41222 1170 41278
rect 1094 41212 1170 41222
rect 1218 42766 1294 42776
rect 1218 42710 1228 42766
rect 1284 42710 1294 42766
rect 1218 42642 1294 42710
rect 1218 42586 1228 42642
rect 1284 42586 1294 42642
rect 1218 42518 1294 42586
rect 1218 42462 1228 42518
rect 1284 42462 1294 42518
rect 1218 42394 1294 42462
rect 1218 42338 1228 42394
rect 1284 42338 1294 42394
rect 1218 42270 1294 42338
rect 1218 42214 1228 42270
rect 1284 42214 1294 42270
rect 1218 42146 1294 42214
rect 1218 42090 1228 42146
rect 1284 42090 1294 42146
rect 1218 42022 1294 42090
rect 1218 41966 1228 42022
rect 1284 41966 1294 42022
rect 1218 41898 1294 41966
rect 1218 41842 1228 41898
rect 1284 41842 1294 41898
rect 1218 41774 1294 41842
rect 1218 41718 1228 41774
rect 1284 41718 1294 41774
rect 1218 41650 1294 41718
rect 1218 41594 1228 41650
rect 1284 41594 1294 41650
rect 1218 41526 1294 41594
rect 1218 41470 1228 41526
rect 1284 41470 1294 41526
rect 1218 41402 1294 41470
rect 1218 41346 1228 41402
rect 1284 41346 1294 41402
rect 1218 41278 1294 41346
rect 1218 41222 1228 41278
rect 1284 41222 1294 41278
rect 1218 41154 1294 41222
rect 1218 41098 1228 41154
rect 1284 41098 1294 41154
rect 1218 41088 1294 41098
rect 1342 42642 1418 42652
rect 1342 42586 1352 42642
rect 1408 42586 1418 42642
rect 1342 42518 1418 42586
rect 1342 42462 1352 42518
rect 1408 42462 1418 42518
rect 1342 42394 1418 42462
rect 1342 42338 1352 42394
rect 1408 42338 1418 42394
rect 1342 42270 1418 42338
rect 1342 42214 1352 42270
rect 1408 42214 1418 42270
rect 1342 42146 1418 42214
rect 1342 42090 1352 42146
rect 1408 42090 1418 42146
rect 1342 42022 1418 42090
rect 1342 41966 1352 42022
rect 1408 41966 1418 42022
rect 1342 41898 1418 41966
rect 1342 41842 1352 41898
rect 1408 41842 1418 41898
rect 1342 41774 1418 41842
rect 1342 41718 1352 41774
rect 1408 41718 1418 41774
rect 1342 41650 1418 41718
rect 1342 41594 1352 41650
rect 1408 41594 1418 41650
rect 1342 41526 1418 41594
rect 1342 41470 1352 41526
rect 1408 41470 1418 41526
rect 1342 41402 1418 41470
rect 1342 41346 1352 41402
rect 1408 41346 1418 41402
rect 1342 41278 1418 41346
rect 1342 41222 1352 41278
rect 1408 41222 1418 41278
rect 1342 41154 1418 41222
rect 1342 41098 1352 41154
rect 1408 41098 1418 41154
rect 1342 41030 1418 41098
rect 1342 40974 1352 41030
rect 1408 40974 1418 41030
rect 1342 40964 1418 40974
rect 1466 42518 1542 42528
rect 1466 42462 1476 42518
rect 1532 42462 1542 42518
rect 1466 42394 1542 42462
rect 1466 42338 1476 42394
rect 1532 42338 1542 42394
rect 1466 42270 1542 42338
rect 1466 42214 1476 42270
rect 1532 42214 1542 42270
rect 1466 42146 1542 42214
rect 1466 42090 1476 42146
rect 1532 42090 1542 42146
rect 1466 42022 1542 42090
rect 1466 41966 1476 42022
rect 1532 41966 1542 42022
rect 1466 41898 1542 41966
rect 1466 41842 1476 41898
rect 1532 41842 1542 41898
rect 1466 41774 1542 41842
rect 1466 41718 1476 41774
rect 1532 41718 1542 41774
rect 1466 41650 1542 41718
rect 1466 41594 1476 41650
rect 1532 41594 1542 41650
rect 1466 41526 1542 41594
rect 1466 41470 1476 41526
rect 1532 41470 1542 41526
rect 1466 41402 1542 41470
rect 1466 41346 1476 41402
rect 1532 41346 1542 41402
rect 1466 41278 1542 41346
rect 1466 41222 1476 41278
rect 1532 41222 1542 41278
rect 1466 41154 1542 41222
rect 1466 41098 1476 41154
rect 1532 41098 1542 41154
rect 1466 41030 1542 41098
rect 1466 40974 1476 41030
rect 1532 40974 1542 41030
rect 1466 40906 1542 40974
rect 1466 40850 1476 40906
rect 1532 40850 1542 40906
rect 1466 40840 1542 40850
rect 1590 42394 1666 42404
rect 1590 42338 1600 42394
rect 1656 42338 1666 42394
rect 1590 42270 1666 42338
rect 1590 42214 1600 42270
rect 1656 42214 1666 42270
rect 1590 42146 1666 42214
rect 1590 42090 1600 42146
rect 1656 42090 1666 42146
rect 1590 42022 1666 42090
rect 1590 41966 1600 42022
rect 1656 41966 1666 42022
rect 1590 41898 1666 41966
rect 1590 41842 1600 41898
rect 1656 41842 1666 41898
rect 1590 41774 1666 41842
rect 1590 41718 1600 41774
rect 1656 41718 1666 41774
rect 1590 41650 1666 41718
rect 1590 41594 1600 41650
rect 1656 41594 1666 41650
rect 1590 41526 1666 41594
rect 1590 41470 1600 41526
rect 1656 41470 1666 41526
rect 1590 41402 1666 41470
rect 1590 41346 1600 41402
rect 1656 41346 1666 41402
rect 1590 41278 1666 41346
rect 1590 41222 1600 41278
rect 1656 41222 1666 41278
rect 1590 41154 1666 41222
rect 1590 41098 1600 41154
rect 1656 41098 1666 41154
rect 1590 41030 1666 41098
rect 1590 40974 1600 41030
rect 1656 40974 1666 41030
rect 1590 40906 1666 40974
rect 1590 40850 1600 40906
rect 1656 40850 1666 40906
rect 1590 40782 1666 40850
rect 1590 40726 1600 40782
rect 1656 40726 1666 40782
rect 1590 40716 1666 40726
rect 1714 42270 1790 42280
rect 1714 42214 1724 42270
rect 1780 42214 1790 42270
rect 1714 42146 1790 42214
rect 1714 42090 1724 42146
rect 1780 42090 1790 42146
rect 1714 42022 1790 42090
rect 1714 41966 1724 42022
rect 1780 41966 1790 42022
rect 1714 41898 1790 41966
rect 1714 41842 1724 41898
rect 1780 41842 1790 41898
rect 1714 41774 1790 41842
rect 1714 41718 1724 41774
rect 1780 41718 1790 41774
rect 1714 41650 1790 41718
rect 1714 41594 1724 41650
rect 1780 41594 1790 41650
rect 1714 41526 1790 41594
rect 1714 41470 1724 41526
rect 1780 41470 1790 41526
rect 1714 41402 1790 41470
rect 1714 41346 1724 41402
rect 1780 41346 1790 41402
rect 1714 41278 1790 41346
rect 1714 41222 1724 41278
rect 1780 41222 1790 41278
rect 1714 41154 1790 41222
rect 1714 41098 1724 41154
rect 1780 41098 1790 41154
rect 1714 41030 1790 41098
rect 1714 40974 1724 41030
rect 1780 40974 1790 41030
rect 1714 40906 1790 40974
rect 1714 40850 1724 40906
rect 1780 40850 1790 40906
rect 1714 40782 1790 40850
rect 1714 40726 1724 40782
rect 1780 40726 1790 40782
rect 1714 40658 1790 40726
rect 1714 40602 1724 40658
rect 1780 40602 1790 40658
rect 1714 40592 1790 40602
rect 1838 42146 1914 42156
rect 1838 42090 1848 42146
rect 1904 42090 1914 42146
rect 1838 42022 1914 42090
rect 1838 41966 1848 42022
rect 1904 41966 1914 42022
rect 1838 41898 1914 41966
rect 1838 41842 1848 41898
rect 1904 41842 1914 41898
rect 1838 41774 1914 41842
rect 1838 41718 1848 41774
rect 1904 41718 1914 41774
rect 1838 41650 1914 41718
rect 1838 41594 1848 41650
rect 1904 41594 1914 41650
rect 1838 41526 1914 41594
rect 1838 41470 1848 41526
rect 1904 41470 1914 41526
rect 1838 41402 1914 41470
rect 1838 41346 1848 41402
rect 1904 41346 1914 41402
rect 1838 41278 1914 41346
rect 1838 41222 1848 41278
rect 1904 41222 1914 41278
rect 1838 41154 1914 41222
rect 1838 41098 1848 41154
rect 1904 41098 1914 41154
rect 1838 41030 1914 41098
rect 1838 40974 1848 41030
rect 1904 40974 1914 41030
rect 1838 40906 1914 40974
rect 1838 40850 1848 40906
rect 1904 40850 1914 40906
rect 1838 40782 1914 40850
rect 1838 40726 1848 40782
rect 1904 40726 1914 40782
rect 1838 40658 1914 40726
rect 1838 40602 1848 40658
rect 1904 40602 1914 40658
rect 1838 40534 1914 40602
rect 1838 40478 1848 40534
rect 1904 40478 1914 40534
rect 1838 40468 1914 40478
rect 1962 42022 2038 42032
rect 1962 41966 1972 42022
rect 2028 41966 2038 42022
rect 1962 41898 2038 41966
rect 1962 41842 1972 41898
rect 2028 41842 2038 41898
rect 1962 41774 2038 41842
rect 1962 41718 1972 41774
rect 2028 41718 2038 41774
rect 1962 41650 2038 41718
rect 1962 41594 1972 41650
rect 2028 41594 2038 41650
rect 1962 41526 2038 41594
rect 1962 41470 1972 41526
rect 2028 41470 2038 41526
rect 1962 41402 2038 41470
rect 1962 41346 1972 41402
rect 2028 41346 2038 41402
rect 1962 41278 2038 41346
rect 1962 41222 1972 41278
rect 2028 41222 2038 41278
rect 1962 41154 2038 41222
rect 1962 41098 1972 41154
rect 2028 41098 2038 41154
rect 1962 41030 2038 41098
rect 1962 40974 1972 41030
rect 2028 40974 2038 41030
rect 1962 40906 2038 40974
rect 1962 40850 1972 40906
rect 2028 40850 2038 40906
rect 1962 40782 2038 40850
rect 1962 40726 1972 40782
rect 2028 40726 2038 40782
rect 1962 40658 2038 40726
rect 1962 40602 1972 40658
rect 2028 40602 2038 40658
rect 1962 40534 2038 40602
rect 1962 40478 1972 40534
rect 2028 40478 2038 40534
rect 1962 40410 2038 40478
rect 1962 40354 1972 40410
rect 2028 40354 2038 40410
rect 1962 40344 2038 40354
rect 4460 39524 4536 39534
rect 4460 39468 4470 39524
rect 4526 39468 4536 39524
rect 4460 39400 4536 39468
rect 4460 39344 4470 39400
rect 4526 39344 4536 39400
rect 4460 39276 4536 39344
rect 4460 39220 4470 39276
rect 4526 39220 4536 39276
rect 2517 39205 2593 39215
rect 2517 39149 2527 39205
rect 2583 39149 2593 39205
rect 2517 39081 2593 39149
rect 4460 39152 4536 39220
rect 4460 39096 4470 39152
rect 4526 39096 4536 39152
rect 2517 39025 2527 39081
rect 2583 39025 2593 39081
rect 2517 38957 2593 39025
rect 2517 38901 2527 38957
rect 2583 38901 2593 38957
rect 2517 38833 2593 38901
rect 2517 38777 2527 38833
rect 2583 38777 2593 38833
rect 2517 38709 2593 38777
rect 2517 38653 2527 38709
rect 2583 38653 2593 38709
rect 2517 38585 2593 38653
rect 2517 38529 2527 38585
rect 2583 38529 2593 38585
rect 2517 38461 2593 38529
rect 2517 38405 2527 38461
rect 2583 38405 2593 38461
rect 2517 38337 2593 38405
rect 2517 38281 2527 38337
rect 2583 38281 2593 38337
rect 2517 38213 2593 38281
rect 2517 38157 2527 38213
rect 2583 38157 2593 38213
rect 2517 38089 2593 38157
rect 2517 38033 2527 38089
rect 2583 38033 2593 38089
rect 2517 37965 2593 38033
rect 2517 37909 2527 37965
rect 2583 37909 2593 37965
rect 2517 37841 2593 37909
rect 2517 37785 2527 37841
rect 2583 37785 2593 37841
rect 2517 37717 2593 37785
rect 2517 37661 2527 37717
rect 2583 37661 2593 37717
rect 2517 37593 2593 37661
rect 2517 37537 2527 37593
rect 2583 37537 2593 37593
rect 2517 37527 2593 37537
rect 2641 39081 2717 39091
rect 2641 39025 2651 39081
rect 2707 39025 2717 39081
rect 2641 38957 2717 39025
rect 4460 39028 4536 39096
rect 4460 38972 4470 39028
rect 4526 38972 4536 39028
rect 2641 38901 2651 38957
rect 2707 38901 2717 38957
rect 2641 38833 2717 38901
rect 2641 38777 2651 38833
rect 2707 38777 2717 38833
rect 2641 38709 2717 38777
rect 2641 38653 2651 38709
rect 2707 38653 2717 38709
rect 2641 38585 2717 38653
rect 2641 38529 2651 38585
rect 2707 38529 2717 38585
rect 2641 38461 2717 38529
rect 2641 38405 2651 38461
rect 2707 38405 2717 38461
rect 2641 38337 2717 38405
rect 2641 38281 2651 38337
rect 2707 38281 2717 38337
rect 2641 38213 2717 38281
rect 2641 38157 2651 38213
rect 2707 38157 2717 38213
rect 2641 38089 2717 38157
rect 2641 38033 2651 38089
rect 2707 38033 2717 38089
rect 2641 37965 2717 38033
rect 2641 37909 2651 37965
rect 2707 37909 2717 37965
rect 2641 37841 2717 37909
rect 2641 37785 2651 37841
rect 2707 37785 2717 37841
rect 2641 37717 2717 37785
rect 2641 37661 2651 37717
rect 2707 37661 2717 37717
rect 2641 37593 2717 37661
rect 2641 37537 2651 37593
rect 2707 37537 2717 37593
rect 2641 37469 2717 37537
rect 2641 37413 2651 37469
rect 2707 37413 2717 37469
rect 2641 37403 2717 37413
rect 2765 38957 2841 38967
rect 2765 38901 2775 38957
rect 2831 38901 2841 38957
rect 2765 38833 2841 38901
rect 4460 38904 4536 38972
rect 4460 38848 4470 38904
rect 4526 38848 4536 38904
rect 2765 38777 2775 38833
rect 2831 38777 2841 38833
rect 2765 38709 2841 38777
rect 2765 38653 2775 38709
rect 2831 38653 2841 38709
rect 2765 38585 2841 38653
rect 2765 38529 2775 38585
rect 2831 38529 2841 38585
rect 2765 38461 2841 38529
rect 2765 38405 2775 38461
rect 2831 38405 2841 38461
rect 2765 38337 2841 38405
rect 2765 38281 2775 38337
rect 2831 38281 2841 38337
rect 2765 38213 2841 38281
rect 2765 38157 2775 38213
rect 2831 38157 2841 38213
rect 2765 38089 2841 38157
rect 2765 38033 2775 38089
rect 2831 38033 2841 38089
rect 2765 37965 2841 38033
rect 2765 37909 2775 37965
rect 2831 37909 2841 37965
rect 2765 37841 2841 37909
rect 2765 37785 2775 37841
rect 2831 37785 2841 37841
rect 2765 37717 2841 37785
rect 2765 37661 2775 37717
rect 2831 37661 2841 37717
rect 2765 37593 2841 37661
rect 2765 37537 2775 37593
rect 2831 37537 2841 37593
rect 2765 37469 2841 37537
rect 2765 37413 2775 37469
rect 2831 37413 2841 37469
rect 2765 37345 2841 37413
rect 2765 37289 2775 37345
rect 2831 37289 2841 37345
rect 2765 37279 2841 37289
rect 2889 38833 2965 38843
rect 2889 38777 2899 38833
rect 2955 38777 2965 38833
rect 2889 38709 2965 38777
rect 4460 38780 4536 38848
rect 4460 38724 4470 38780
rect 4526 38724 4536 38780
rect 2889 38653 2899 38709
rect 2955 38653 2965 38709
rect 2889 38585 2965 38653
rect 2889 38529 2899 38585
rect 2955 38529 2965 38585
rect 2889 38461 2965 38529
rect 2889 38405 2899 38461
rect 2955 38405 2965 38461
rect 2889 38337 2965 38405
rect 2889 38281 2899 38337
rect 2955 38281 2965 38337
rect 2889 38213 2965 38281
rect 2889 38157 2899 38213
rect 2955 38157 2965 38213
rect 2889 38089 2965 38157
rect 2889 38033 2899 38089
rect 2955 38033 2965 38089
rect 2889 37965 2965 38033
rect 2889 37909 2899 37965
rect 2955 37909 2965 37965
rect 2889 37841 2965 37909
rect 2889 37785 2899 37841
rect 2955 37785 2965 37841
rect 2889 37717 2965 37785
rect 2889 37661 2899 37717
rect 2955 37661 2965 37717
rect 2889 37593 2965 37661
rect 2889 37537 2899 37593
rect 2955 37537 2965 37593
rect 2889 37469 2965 37537
rect 2889 37413 2899 37469
rect 2955 37413 2965 37469
rect 2889 37345 2965 37413
rect 2889 37289 2899 37345
rect 2955 37289 2965 37345
rect 2889 37221 2965 37289
rect 2889 37165 2899 37221
rect 2955 37165 2965 37221
rect 2889 37155 2965 37165
rect 3013 38709 3089 38719
rect 3013 38653 3023 38709
rect 3079 38653 3089 38709
rect 3013 38585 3089 38653
rect 4460 38656 4536 38724
rect 4460 38600 4470 38656
rect 4526 38600 4536 38656
rect 3013 38529 3023 38585
rect 3079 38529 3089 38585
rect 3013 38461 3089 38529
rect 3013 38405 3023 38461
rect 3079 38405 3089 38461
rect 3013 38337 3089 38405
rect 3013 38281 3023 38337
rect 3079 38281 3089 38337
rect 3013 38213 3089 38281
rect 3013 38157 3023 38213
rect 3079 38157 3089 38213
rect 3013 38089 3089 38157
rect 3013 38033 3023 38089
rect 3079 38033 3089 38089
rect 3013 37965 3089 38033
rect 3013 37909 3023 37965
rect 3079 37909 3089 37965
rect 3013 37841 3089 37909
rect 3013 37785 3023 37841
rect 3079 37785 3089 37841
rect 3013 37717 3089 37785
rect 3013 37661 3023 37717
rect 3079 37661 3089 37717
rect 3013 37593 3089 37661
rect 3013 37537 3023 37593
rect 3079 37537 3089 37593
rect 3013 37469 3089 37537
rect 3013 37413 3023 37469
rect 3079 37413 3089 37469
rect 3013 37345 3089 37413
rect 3013 37289 3023 37345
rect 3079 37289 3089 37345
rect 3013 37221 3089 37289
rect 3013 37165 3023 37221
rect 3079 37165 3089 37221
rect 3013 37097 3089 37165
rect 3013 37041 3023 37097
rect 3079 37041 3089 37097
rect 3013 37031 3089 37041
rect 3137 38585 3213 38595
rect 3137 38529 3147 38585
rect 3203 38529 3213 38585
rect 3137 38461 3213 38529
rect 4460 38532 4536 38600
rect 4460 38476 4470 38532
rect 4526 38476 4536 38532
rect 3137 38405 3147 38461
rect 3203 38405 3213 38461
rect 3137 38337 3213 38405
rect 3137 38281 3147 38337
rect 3203 38281 3213 38337
rect 3137 38213 3213 38281
rect 3137 38157 3147 38213
rect 3203 38157 3213 38213
rect 3137 38089 3213 38157
rect 3137 38033 3147 38089
rect 3203 38033 3213 38089
rect 3137 37965 3213 38033
rect 3137 37909 3147 37965
rect 3203 37909 3213 37965
rect 3137 37841 3213 37909
rect 3137 37785 3147 37841
rect 3203 37785 3213 37841
rect 3137 37717 3213 37785
rect 3137 37661 3147 37717
rect 3203 37661 3213 37717
rect 3137 37593 3213 37661
rect 3137 37537 3147 37593
rect 3203 37537 3213 37593
rect 3137 37469 3213 37537
rect 3137 37413 3147 37469
rect 3203 37413 3213 37469
rect 3137 37345 3213 37413
rect 3137 37289 3147 37345
rect 3203 37289 3213 37345
rect 3137 37221 3213 37289
rect 3137 37165 3147 37221
rect 3203 37165 3213 37221
rect 3137 37097 3213 37165
rect 3137 37041 3147 37097
rect 3203 37041 3213 37097
rect 3137 36973 3213 37041
rect 3137 36917 3147 36973
rect 3203 36917 3213 36973
rect 3137 36907 3213 36917
rect 3261 38461 3337 38471
rect 3261 38405 3271 38461
rect 3327 38405 3337 38461
rect 3261 38337 3337 38405
rect 4460 38408 4536 38476
rect 4460 38352 4470 38408
rect 4526 38352 4536 38408
rect 3261 38281 3271 38337
rect 3327 38281 3337 38337
rect 3261 38213 3337 38281
rect 3261 38157 3271 38213
rect 3327 38157 3337 38213
rect 3261 38089 3337 38157
rect 3261 38033 3271 38089
rect 3327 38033 3337 38089
rect 3261 37965 3337 38033
rect 3261 37909 3271 37965
rect 3327 37909 3337 37965
rect 3261 37841 3337 37909
rect 3261 37785 3271 37841
rect 3327 37785 3337 37841
rect 3261 37717 3337 37785
rect 3261 37661 3271 37717
rect 3327 37661 3337 37717
rect 3261 37593 3337 37661
rect 3261 37537 3271 37593
rect 3327 37537 3337 37593
rect 3261 37469 3337 37537
rect 3261 37413 3271 37469
rect 3327 37413 3337 37469
rect 3261 37345 3337 37413
rect 3261 37289 3271 37345
rect 3327 37289 3337 37345
rect 3261 37221 3337 37289
rect 3261 37165 3271 37221
rect 3327 37165 3337 37221
rect 3261 37097 3337 37165
rect 3261 37041 3271 37097
rect 3327 37041 3337 37097
rect 3261 36973 3337 37041
rect 3261 36917 3271 36973
rect 3327 36917 3337 36973
rect 3261 36849 3337 36917
rect 3261 36793 3271 36849
rect 3327 36793 3337 36849
rect 3261 36783 3337 36793
rect 3385 38337 3461 38347
rect 3385 38281 3395 38337
rect 3451 38281 3461 38337
rect 3385 38213 3461 38281
rect 4460 38284 4536 38352
rect 4460 38228 4470 38284
rect 4526 38228 4536 38284
rect 3385 38157 3395 38213
rect 3451 38157 3461 38213
rect 3385 38089 3461 38157
rect 3385 38033 3395 38089
rect 3451 38033 3461 38089
rect 3385 37965 3461 38033
rect 3385 37909 3395 37965
rect 3451 37909 3461 37965
rect 3385 37841 3461 37909
rect 3385 37785 3395 37841
rect 3451 37785 3461 37841
rect 3385 37717 3461 37785
rect 3385 37661 3395 37717
rect 3451 37661 3461 37717
rect 3385 37593 3461 37661
rect 3385 37537 3395 37593
rect 3451 37537 3461 37593
rect 3385 37469 3461 37537
rect 3385 37413 3395 37469
rect 3451 37413 3461 37469
rect 3385 37345 3461 37413
rect 3385 37289 3395 37345
rect 3451 37289 3461 37345
rect 3385 37221 3461 37289
rect 3385 37165 3395 37221
rect 3451 37165 3461 37221
rect 3385 37097 3461 37165
rect 3385 37041 3395 37097
rect 3451 37041 3461 37097
rect 3385 36973 3461 37041
rect 3385 36917 3395 36973
rect 3451 36917 3461 36973
rect 3385 36849 3461 36917
rect 3385 36793 3395 36849
rect 3451 36793 3461 36849
rect 3385 36725 3461 36793
rect 3385 36669 3395 36725
rect 3451 36669 3461 36725
rect 3385 36659 3461 36669
rect 3509 38213 3585 38223
rect 3509 38157 3519 38213
rect 3575 38157 3585 38213
rect 3509 38089 3585 38157
rect 4460 38160 4536 38228
rect 4460 38104 4470 38160
rect 4526 38104 4536 38160
rect 3509 38033 3519 38089
rect 3575 38033 3585 38089
rect 3509 37965 3585 38033
rect 3509 37909 3519 37965
rect 3575 37909 3585 37965
rect 3509 37841 3585 37909
rect 3509 37785 3519 37841
rect 3575 37785 3585 37841
rect 3509 37717 3585 37785
rect 3509 37661 3519 37717
rect 3575 37661 3585 37717
rect 3509 37593 3585 37661
rect 3509 37537 3519 37593
rect 3575 37537 3585 37593
rect 3509 37469 3585 37537
rect 3509 37413 3519 37469
rect 3575 37413 3585 37469
rect 3509 37345 3585 37413
rect 3509 37289 3519 37345
rect 3575 37289 3585 37345
rect 3509 37221 3585 37289
rect 3509 37165 3519 37221
rect 3575 37165 3585 37221
rect 3509 37097 3585 37165
rect 3509 37041 3519 37097
rect 3575 37041 3585 37097
rect 3509 36973 3585 37041
rect 3509 36917 3519 36973
rect 3575 36917 3585 36973
rect 3509 36849 3585 36917
rect 3509 36793 3519 36849
rect 3575 36793 3585 36849
rect 3509 36725 3585 36793
rect 3509 36669 3519 36725
rect 3575 36669 3585 36725
rect 3509 36601 3585 36669
rect 3509 36545 3519 36601
rect 3575 36545 3585 36601
rect 3509 36535 3585 36545
rect 3633 38089 3709 38099
rect 3633 38033 3643 38089
rect 3699 38033 3709 38089
rect 3633 37965 3709 38033
rect 4460 38036 4536 38104
rect 4460 37980 4470 38036
rect 4526 37980 4536 38036
rect 3633 37909 3643 37965
rect 3699 37909 3709 37965
rect 3633 37841 3709 37909
rect 3633 37785 3643 37841
rect 3699 37785 3709 37841
rect 3633 37717 3709 37785
rect 3633 37661 3643 37717
rect 3699 37661 3709 37717
rect 3633 37593 3709 37661
rect 3633 37537 3643 37593
rect 3699 37537 3709 37593
rect 3633 37469 3709 37537
rect 3633 37413 3643 37469
rect 3699 37413 3709 37469
rect 3633 37345 3709 37413
rect 3633 37289 3643 37345
rect 3699 37289 3709 37345
rect 3633 37221 3709 37289
rect 3633 37165 3643 37221
rect 3699 37165 3709 37221
rect 3633 37097 3709 37165
rect 3633 37041 3643 37097
rect 3699 37041 3709 37097
rect 3633 36973 3709 37041
rect 3633 36917 3643 36973
rect 3699 36917 3709 36973
rect 3633 36849 3709 36917
rect 3633 36793 3643 36849
rect 3699 36793 3709 36849
rect 3633 36725 3709 36793
rect 3633 36669 3643 36725
rect 3699 36669 3709 36725
rect 3633 36601 3709 36669
rect 3633 36545 3643 36601
rect 3699 36545 3709 36601
rect 3633 36477 3709 36545
rect 3633 36421 3643 36477
rect 3699 36421 3709 36477
rect 3633 36411 3709 36421
rect 3757 37965 3833 37975
rect 3757 37909 3767 37965
rect 3823 37909 3833 37965
rect 3757 37841 3833 37909
rect 4460 37912 4536 37980
rect 4460 37856 4470 37912
rect 4526 37856 4536 37912
rect 3757 37785 3767 37841
rect 3823 37785 3833 37841
rect 3757 37717 3833 37785
rect 3757 37661 3767 37717
rect 3823 37661 3833 37717
rect 3757 37593 3833 37661
rect 3757 37537 3767 37593
rect 3823 37537 3833 37593
rect 3757 37469 3833 37537
rect 3757 37413 3767 37469
rect 3823 37413 3833 37469
rect 3757 37345 3833 37413
rect 3757 37289 3767 37345
rect 3823 37289 3833 37345
rect 3757 37221 3833 37289
rect 3757 37165 3767 37221
rect 3823 37165 3833 37221
rect 3757 37097 3833 37165
rect 3757 37041 3767 37097
rect 3823 37041 3833 37097
rect 3757 36973 3833 37041
rect 3757 36917 3767 36973
rect 3823 36917 3833 36973
rect 3757 36849 3833 36917
rect 3757 36793 3767 36849
rect 3823 36793 3833 36849
rect 3757 36725 3833 36793
rect 3757 36669 3767 36725
rect 3823 36669 3833 36725
rect 3757 36601 3833 36669
rect 3757 36545 3767 36601
rect 3823 36545 3833 36601
rect 3757 36477 3833 36545
rect 3757 36421 3767 36477
rect 3823 36421 3833 36477
rect 3757 36353 3833 36421
rect 3757 36297 3767 36353
rect 3823 36297 3833 36353
rect 3757 36287 3833 36297
rect 3881 37841 3957 37851
rect 4460 37846 4536 37856
rect 4584 39400 4660 39410
rect 4584 39344 4594 39400
rect 4650 39344 4660 39400
rect 4584 39276 4660 39344
rect 4584 39220 4594 39276
rect 4650 39220 4660 39276
rect 4584 39152 4660 39220
rect 4584 39096 4594 39152
rect 4650 39096 4660 39152
rect 4584 39028 4660 39096
rect 4584 38972 4594 39028
rect 4650 38972 4660 39028
rect 4584 38904 4660 38972
rect 4584 38848 4594 38904
rect 4650 38848 4660 38904
rect 4584 38780 4660 38848
rect 4584 38724 4594 38780
rect 4650 38724 4660 38780
rect 4584 38656 4660 38724
rect 4584 38600 4594 38656
rect 4650 38600 4660 38656
rect 4584 38532 4660 38600
rect 4584 38476 4594 38532
rect 4650 38476 4660 38532
rect 4584 38408 4660 38476
rect 4584 38352 4594 38408
rect 4650 38352 4660 38408
rect 4584 38284 4660 38352
rect 4584 38228 4594 38284
rect 4650 38228 4660 38284
rect 4584 38160 4660 38228
rect 4584 38104 4594 38160
rect 4650 38104 4660 38160
rect 4584 38036 4660 38104
rect 4584 37980 4594 38036
rect 4650 37980 4660 38036
rect 4584 37912 4660 37980
rect 4584 37856 4594 37912
rect 4650 37856 4660 37912
rect 3881 37785 3891 37841
rect 3947 37785 3957 37841
rect 3881 37717 3957 37785
rect 4584 37788 4660 37856
rect 4584 37732 4594 37788
rect 4650 37732 4660 37788
rect 3881 37661 3891 37717
rect 3947 37661 3957 37717
rect 3881 37593 3957 37661
rect 3881 37537 3891 37593
rect 3947 37537 3957 37593
rect 3881 37469 3957 37537
rect 3881 37413 3891 37469
rect 3947 37413 3957 37469
rect 3881 37345 3957 37413
rect 3881 37289 3891 37345
rect 3947 37289 3957 37345
rect 3881 37221 3957 37289
rect 3881 37165 3891 37221
rect 3947 37165 3957 37221
rect 3881 37097 3957 37165
rect 3881 37041 3891 37097
rect 3947 37041 3957 37097
rect 3881 36973 3957 37041
rect 3881 36917 3891 36973
rect 3947 36917 3957 36973
rect 3881 36849 3957 36917
rect 3881 36793 3891 36849
rect 3947 36793 3957 36849
rect 3881 36725 3957 36793
rect 3881 36669 3891 36725
rect 3947 36669 3957 36725
rect 3881 36601 3957 36669
rect 3881 36545 3891 36601
rect 3947 36545 3957 36601
rect 3881 36477 3957 36545
rect 3881 36421 3891 36477
rect 3947 36421 3957 36477
rect 3881 36353 3957 36421
rect 3881 36297 3891 36353
rect 3947 36297 3957 36353
rect 3881 36229 3957 36297
rect 3881 36173 3891 36229
rect 3947 36173 3957 36229
rect 3881 36163 3957 36173
rect 4005 37717 4081 37727
rect 4584 37722 4660 37732
rect 4708 39276 4784 39286
rect 4708 39220 4718 39276
rect 4774 39220 4784 39276
rect 4708 39152 4784 39220
rect 4708 39096 4718 39152
rect 4774 39096 4784 39152
rect 4708 39028 4784 39096
rect 4708 38972 4718 39028
rect 4774 38972 4784 39028
rect 4708 38904 4784 38972
rect 4708 38848 4718 38904
rect 4774 38848 4784 38904
rect 4708 38780 4784 38848
rect 4708 38724 4718 38780
rect 4774 38724 4784 38780
rect 4708 38656 4784 38724
rect 4708 38600 4718 38656
rect 4774 38600 4784 38656
rect 4708 38532 4784 38600
rect 4708 38476 4718 38532
rect 4774 38476 4784 38532
rect 4708 38408 4784 38476
rect 4708 38352 4718 38408
rect 4774 38352 4784 38408
rect 4708 38284 4784 38352
rect 4708 38228 4718 38284
rect 4774 38228 4784 38284
rect 4708 38160 4784 38228
rect 4708 38104 4718 38160
rect 4774 38104 4784 38160
rect 4708 38036 4784 38104
rect 4708 37980 4718 38036
rect 4774 37980 4784 38036
rect 4708 37912 4784 37980
rect 4708 37856 4718 37912
rect 4774 37856 4784 37912
rect 4708 37788 4784 37856
rect 4708 37732 4718 37788
rect 4774 37732 4784 37788
rect 4005 37661 4015 37717
rect 4071 37661 4081 37717
rect 4005 37593 4081 37661
rect 4708 37664 4784 37732
rect 4708 37608 4718 37664
rect 4774 37608 4784 37664
rect 4005 37537 4015 37593
rect 4071 37537 4081 37593
rect 4005 37469 4081 37537
rect 4005 37413 4015 37469
rect 4071 37413 4081 37469
rect 4005 37345 4081 37413
rect 4005 37289 4015 37345
rect 4071 37289 4081 37345
rect 4005 37221 4081 37289
rect 4005 37165 4015 37221
rect 4071 37165 4081 37221
rect 4005 37097 4081 37165
rect 4005 37041 4015 37097
rect 4071 37041 4081 37097
rect 4005 36973 4081 37041
rect 4005 36917 4015 36973
rect 4071 36917 4081 36973
rect 4005 36849 4081 36917
rect 4005 36793 4015 36849
rect 4071 36793 4081 36849
rect 4005 36725 4081 36793
rect 4005 36669 4015 36725
rect 4071 36669 4081 36725
rect 4005 36601 4081 36669
rect 4005 36545 4015 36601
rect 4071 36545 4081 36601
rect 4005 36477 4081 36545
rect 4005 36421 4015 36477
rect 4071 36421 4081 36477
rect 4005 36353 4081 36421
rect 4005 36297 4015 36353
rect 4071 36297 4081 36353
rect 4005 36229 4081 36297
rect 4005 36173 4015 36229
rect 4071 36173 4081 36229
rect 4005 36105 4081 36173
rect 4005 36049 4015 36105
rect 4071 36049 4081 36105
rect 4005 36039 4081 36049
rect 4129 37593 4205 37603
rect 4708 37598 4784 37608
rect 4832 39152 4908 39162
rect 4832 39096 4842 39152
rect 4898 39096 4908 39152
rect 4832 39028 4908 39096
rect 4832 38972 4842 39028
rect 4898 38972 4908 39028
rect 4832 38904 4908 38972
rect 4832 38848 4842 38904
rect 4898 38848 4908 38904
rect 4832 38780 4908 38848
rect 4832 38724 4842 38780
rect 4898 38724 4908 38780
rect 4832 38656 4908 38724
rect 4832 38600 4842 38656
rect 4898 38600 4908 38656
rect 4832 38532 4908 38600
rect 4832 38476 4842 38532
rect 4898 38476 4908 38532
rect 4832 38408 4908 38476
rect 4832 38352 4842 38408
rect 4898 38352 4908 38408
rect 4832 38284 4908 38352
rect 4832 38228 4842 38284
rect 4898 38228 4908 38284
rect 4832 38160 4908 38228
rect 4832 38104 4842 38160
rect 4898 38104 4908 38160
rect 4832 38036 4908 38104
rect 4832 37980 4842 38036
rect 4898 37980 4908 38036
rect 4832 37912 4908 37980
rect 4832 37856 4842 37912
rect 4898 37856 4908 37912
rect 4832 37788 4908 37856
rect 4832 37732 4842 37788
rect 4898 37732 4908 37788
rect 4832 37664 4908 37732
rect 4832 37608 4842 37664
rect 4898 37608 4908 37664
rect 4129 37537 4139 37593
rect 4195 37537 4205 37593
rect 4129 37469 4205 37537
rect 4832 37540 4908 37608
rect 4832 37484 4842 37540
rect 4898 37484 4908 37540
rect 4832 37474 4908 37484
rect 4956 39028 5032 39038
rect 4956 38972 4966 39028
rect 5022 38972 5032 39028
rect 4956 38904 5032 38972
rect 4956 38848 4966 38904
rect 5022 38848 5032 38904
rect 4956 38780 5032 38848
rect 4956 38724 4966 38780
rect 5022 38724 5032 38780
rect 4956 38656 5032 38724
rect 4956 38600 4966 38656
rect 5022 38600 5032 38656
rect 4956 38532 5032 38600
rect 4956 38476 4966 38532
rect 5022 38476 5032 38532
rect 4956 38408 5032 38476
rect 4956 38352 4966 38408
rect 5022 38352 5032 38408
rect 4956 38284 5032 38352
rect 4956 38228 4966 38284
rect 5022 38228 5032 38284
rect 4956 38160 5032 38228
rect 4956 38104 4966 38160
rect 5022 38104 5032 38160
rect 4956 38036 5032 38104
rect 4956 37980 4966 38036
rect 5022 37980 5032 38036
rect 4956 37912 5032 37980
rect 4956 37856 4966 37912
rect 5022 37856 5032 37912
rect 4956 37788 5032 37856
rect 4956 37732 4966 37788
rect 5022 37732 5032 37788
rect 4956 37664 5032 37732
rect 4956 37608 4966 37664
rect 5022 37608 5032 37664
rect 4956 37540 5032 37608
rect 4956 37484 4966 37540
rect 5022 37484 5032 37540
rect 4129 37413 4139 37469
rect 4195 37413 4205 37469
rect 4129 37345 4205 37413
rect 4956 37416 5032 37484
rect 4956 37360 4966 37416
rect 5022 37360 5032 37416
rect 4956 37350 5032 37360
rect 5080 38904 5156 38914
rect 5080 38848 5090 38904
rect 5146 38848 5156 38904
rect 5080 38780 5156 38848
rect 5080 38724 5090 38780
rect 5146 38724 5156 38780
rect 5080 38656 5156 38724
rect 5080 38600 5090 38656
rect 5146 38600 5156 38656
rect 5080 38532 5156 38600
rect 5080 38476 5090 38532
rect 5146 38476 5156 38532
rect 5080 38408 5156 38476
rect 5080 38352 5090 38408
rect 5146 38352 5156 38408
rect 5080 38284 5156 38352
rect 5080 38228 5090 38284
rect 5146 38228 5156 38284
rect 5080 38160 5156 38228
rect 5080 38104 5090 38160
rect 5146 38104 5156 38160
rect 5080 38036 5156 38104
rect 5080 37980 5090 38036
rect 5146 37980 5156 38036
rect 5080 37912 5156 37980
rect 5080 37856 5090 37912
rect 5146 37856 5156 37912
rect 5080 37788 5156 37856
rect 5080 37732 5090 37788
rect 5146 37732 5156 37788
rect 5080 37664 5156 37732
rect 5080 37608 5090 37664
rect 5146 37608 5156 37664
rect 5080 37540 5156 37608
rect 5080 37484 5090 37540
rect 5146 37484 5156 37540
rect 5080 37416 5156 37484
rect 5080 37360 5090 37416
rect 5146 37360 5156 37416
rect 4129 37289 4139 37345
rect 4195 37289 4205 37345
rect 4129 37221 4205 37289
rect 5080 37292 5156 37360
rect 5080 37236 5090 37292
rect 5146 37236 5156 37292
rect 5080 37226 5156 37236
rect 5204 38780 5280 38790
rect 5204 38724 5214 38780
rect 5270 38724 5280 38780
rect 5204 38656 5280 38724
rect 5204 38600 5214 38656
rect 5270 38600 5280 38656
rect 5204 38532 5280 38600
rect 5204 38476 5214 38532
rect 5270 38476 5280 38532
rect 5204 38408 5280 38476
rect 5204 38352 5214 38408
rect 5270 38352 5280 38408
rect 5204 38284 5280 38352
rect 5204 38228 5214 38284
rect 5270 38228 5280 38284
rect 5204 38160 5280 38228
rect 5204 38104 5214 38160
rect 5270 38104 5280 38160
rect 5204 38036 5280 38104
rect 5204 37980 5214 38036
rect 5270 37980 5280 38036
rect 5204 37912 5280 37980
rect 5204 37856 5214 37912
rect 5270 37856 5280 37912
rect 5204 37788 5280 37856
rect 5204 37732 5214 37788
rect 5270 37732 5280 37788
rect 5204 37664 5280 37732
rect 5204 37608 5214 37664
rect 5270 37608 5280 37664
rect 5204 37540 5280 37608
rect 5204 37484 5214 37540
rect 5270 37484 5280 37540
rect 5204 37416 5280 37484
rect 5204 37360 5214 37416
rect 5270 37360 5280 37416
rect 5204 37292 5280 37360
rect 5204 37236 5214 37292
rect 5270 37236 5280 37292
rect 4129 37165 4139 37221
rect 4195 37165 4205 37221
rect 4129 37097 4205 37165
rect 5204 37168 5280 37236
rect 5204 37112 5214 37168
rect 5270 37112 5280 37168
rect 5204 37102 5280 37112
rect 5328 38656 5404 38666
rect 5328 38600 5338 38656
rect 5394 38600 5404 38656
rect 5328 38532 5404 38600
rect 5328 38476 5338 38532
rect 5394 38476 5404 38532
rect 5328 38408 5404 38476
rect 5328 38352 5338 38408
rect 5394 38352 5404 38408
rect 5328 38284 5404 38352
rect 5328 38228 5338 38284
rect 5394 38228 5404 38284
rect 5328 38160 5404 38228
rect 5328 38104 5338 38160
rect 5394 38104 5404 38160
rect 5328 38036 5404 38104
rect 5328 37980 5338 38036
rect 5394 37980 5404 38036
rect 5328 37912 5404 37980
rect 5328 37856 5338 37912
rect 5394 37856 5404 37912
rect 5328 37788 5404 37856
rect 5328 37732 5338 37788
rect 5394 37732 5404 37788
rect 5328 37664 5404 37732
rect 5328 37608 5338 37664
rect 5394 37608 5404 37664
rect 5328 37540 5404 37608
rect 5328 37484 5338 37540
rect 5394 37484 5404 37540
rect 5328 37416 5404 37484
rect 5328 37360 5338 37416
rect 5394 37360 5404 37416
rect 5328 37292 5404 37360
rect 5328 37236 5338 37292
rect 5394 37236 5404 37292
rect 5328 37168 5404 37236
rect 5328 37112 5338 37168
rect 5394 37112 5404 37168
rect 4129 37041 4139 37097
rect 4195 37041 4205 37097
rect 4129 36973 4205 37041
rect 5328 37044 5404 37112
rect 5328 36988 5338 37044
rect 5394 36988 5404 37044
rect 5328 36978 5404 36988
rect 5452 38532 5528 38542
rect 5452 38476 5462 38532
rect 5518 38476 5528 38532
rect 5452 38408 5528 38476
rect 5452 38352 5462 38408
rect 5518 38352 5528 38408
rect 5452 38284 5528 38352
rect 5452 38228 5462 38284
rect 5518 38228 5528 38284
rect 5452 38160 5528 38228
rect 5452 38104 5462 38160
rect 5518 38104 5528 38160
rect 5452 38036 5528 38104
rect 5452 37980 5462 38036
rect 5518 37980 5528 38036
rect 5452 37912 5528 37980
rect 5452 37856 5462 37912
rect 5518 37856 5528 37912
rect 5452 37788 5528 37856
rect 5452 37732 5462 37788
rect 5518 37732 5528 37788
rect 5452 37664 5528 37732
rect 5452 37608 5462 37664
rect 5518 37608 5528 37664
rect 5452 37540 5528 37608
rect 5452 37484 5462 37540
rect 5518 37484 5528 37540
rect 5452 37416 5528 37484
rect 5452 37360 5462 37416
rect 5518 37360 5528 37416
rect 5452 37292 5528 37360
rect 5452 37236 5462 37292
rect 5518 37236 5528 37292
rect 5452 37168 5528 37236
rect 5452 37112 5462 37168
rect 5518 37112 5528 37168
rect 5452 37044 5528 37112
rect 5452 36988 5462 37044
rect 5518 36988 5528 37044
rect 4129 36917 4139 36973
rect 4195 36917 4205 36973
rect 4129 36849 4205 36917
rect 5452 36920 5528 36988
rect 5452 36864 5462 36920
rect 5518 36864 5528 36920
rect 5452 36854 5528 36864
rect 5576 38402 5652 38412
rect 5576 38346 5586 38402
rect 5642 38346 5652 38402
rect 5576 38278 5652 38346
rect 5576 38222 5586 38278
rect 5642 38222 5652 38278
rect 5576 38154 5652 38222
rect 5576 38098 5586 38154
rect 5642 38098 5652 38154
rect 5576 38030 5652 38098
rect 5576 37974 5586 38030
rect 5642 37974 5652 38030
rect 5576 37906 5652 37974
rect 5576 37850 5586 37906
rect 5642 37850 5652 37906
rect 5576 37782 5652 37850
rect 5576 37726 5586 37782
rect 5642 37726 5652 37782
rect 5576 37658 5652 37726
rect 5576 37602 5586 37658
rect 5642 37602 5652 37658
rect 5576 37534 5652 37602
rect 5576 37478 5586 37534
rect 5642 37478 5652 37534
rect 5576 37410 5652 37478
rect 5576 37354 5586 37410
rect 5642 37354 5652 37410
rect 5576 37286 5652 37354
rect 5576 37230 5586 37286
rect 5642 37230 5652 37286
rect 5576 37162 5652 37230
rect 5576 37106 5586 37162
rect 5642 37106 5652 37162
rect 5576 37038 5652 37106
rect 5576 36982 5586 37038
rect 5642 36982 5652 37038
rect 5576 36914 5652 36982
rect 5576 36858 5586 36914
rect 5642 36858 5652 36914
rect 4129 36793 4139 36849
rect 4195 36793 4205 36849
rect 5576 36848 5652 36858
rect 5700 38273 5776 38283
rect 5700 38217 5710 38273
rect 5766 38217 5776 38273
rect 5700 38149 5776 38217
rect 5700 38093 5710 38149
rect 5766 38093 5776 38149
rect 5700 38025 5776 38093
rect 5700 37969 5710 38025
rect 5766 37969 5776 38025
rect 5700 37901 5776 37969
rect 5700 37845 5710 37901
rect 5766 37845 5776 37901
rect 5700 37777 5776 37845
rect 5700 37721 5710 37777
rect 5766 37721 5776 37777
rect 5700 37653 5776 37721
rect 5700 37597 5710 37653
rect 5766 37597 5776 37653
rect 5700 37529 5776 37597
rect 5700 37473 5710 37529
rect 5766 37473 5776 37529
rect 5700 37405 5776 37473
rect 5700 37349 5710 37405
rect 5766 37349 5776 37405
rect 5700 37281 5776 37349
rect 5700 37225 5710 37281
rect 5766 37225 5776 37281
rect 5700 37157 5776 37225
rect 5700 37101 5710 37157
rect 5766 37101 5776 37157
rect 5700 37033 5776 37101
rect 5700 36977 5710 37033
rect 5766 36977 5776 37033
rect 5700 36909 5776 36977
rect 5700 36853 5710 36909
rect 5766 36853 5776 36909
rect 5824 38162 5900 38172
rect 5824 38106 5834 38162
rect 5890 38106 5900 38162
rect 5824 38038 5900 38106
rect 5824 37982 5834 38038
rect 5890 37982 5900 38038
rect 5824 37914 5900 37982
rect 5824 37858 5834 37914
rect 5890 37858 5900 37914
rect 5824 37790 5900 37858
rect 5824 37734 5834 37790
rect 5890 37734 5900 37790
rect 5824 37666 5900 37734
rect 5824 37610 5834 37666
rect 5890 37610 5900 37666
rect 5824 37542 5900 37610
rect 5824 37486 5834 37542
rect 5890 37486 5900 37542
rect 5824 37418 5900 37486
rect 5824 37362 5834 37418
rect 5890 37362 5900 37418
rect 5824 37294 5900 37362
rect 5824 37238 5834 37294
rect 5890 37238 5900 37294
rect 5824 37170 5900 37238
rect 5824 37114 5834 37170
rect 5890 37114 5900 37170
rect 5824 37046 5900 37114
rect 5824 36990 5834 37046
rect 5890 36990 5900 37046
rect 5824 36922 5900 36990
rect 5824 36866 5834 36922
rect 5890 36866 5900 36922
rect 5824 36856 5900 36866
rect 5948 38141 6024 38151
rect 5948 38085 5958 38141
rect 6014 38085 6024 38141
rect 5948 38017 6024 38085
rect 5948 37961 5958 38017
rect 6014 37961 6024 38017
rect 5948 37893 6024 37961
rect 5948 37837 5958 37893
rect 6014 37837 6024 37893
rect 5948 37769 6024 37837
rect 5948 37713 5958 37769
rect 6014 37713 6024 37769
rect 5948 37645 6024 37713
rect 5948 37589 5958 37645
rect 6014 37589 6024 37645
rect 5948 37521 6024 37589
rect 5948 37465 5958 37521
rect 6014 37465 6024 37521
rect 5948 37397 6024 37465
rect 5948 37341 5958 37397
rect 6014 37341 6024 37397
rect 5948 37273 6024 37341
rect 5948 37217 5958 37273
rect 6014 37217 6024 37273
rect 5948 37149 6024 37217
rect 5948 37093 5958 37149
rect 6014 37093 6024 37149
rect 5948 37025 6024 37093
rect 5948 36969 5958 37025
rect 6014 36969 6024 37025
rect 5948 36901 6024 36969
rect 5700 36843 5776 36853
rect 5948 36845 5958 36901
rect 6014 36845 6024 36901
rect 5948 36835 6024 36845
rect 6072 38140 6148 38150
rect 6072 38084 6082 38140
rect 6138 38084 6148 38140
rect 6072 38016 6148 38084
rect 6072 37960 6082 38016
rect 6138 37960 6148 38016
rect 6072 37892 6148 37960
rect 6072 37836 6082 37892
rect 6138 37836 6148 37892
rect 6072 37768 6148 37836
rect 6072 37712 6082 37768
rect 6138 37712 6148 37768
rect 6072 37644 6148 37712
rect 6072 37588 6082 37644
rect 6138 37588 6148 37644
rect 6072 37520 6148 37588
rect 6072 37464 6082 37520
rect 6138 37464 6148 37520
rect 6072 37396 6148 37464
rect 6072 37340 6082 37396
rect 6138 37340 6148 37396
rect 6072 37272 6148 37340
rect 6072 37216 6082 37272
rect 6138 37216 6148 37272
rect 6072 37148 6148 37216
rect 6072 37092 6082 37148
rect 6138 37092 6148 37148
rect 6072 37024 6148 37092
rect 6072 36968 6082 37024
rect 6138 36968 6148 37024
rect 6072 36900 6148 36968
rect 6072 36844 6082 36900
rect 6138 36844 6148 36900
rect 6072 36834 6148 36844
rect 7552 38144 8620 38154
rect 7552 38088 7562 38144
rect 7618 38088 7686 38144
rect 7742 38088 7810 38144
rect 7866 38088 7934 38144
rect 7990 38088 8058 38144
rect 8114 38088 8182 38144
rect 8238 38088 8306 38144
rect 8362 38088 8430 38144
rect 8486 38088 8554 38144
rect 8610 38088 8620 38144
rect 7552 38020 8620 38088
rect 7552 37964 7562 38020
rect 7618 37964 7686 38020
rect 7742 37964 7810 38020
rect 7866 37964 7934 38020
rect 7990 37964 8058 38020
rect 8114 37964 8182 38020
rect 8238 37964 8306 38020
rect 8362 37964 8430 38020
rect 8486 37964 8554 38020
rect 8610 37964 8620 38020
rect 7552 37896 8620 37964
rect 7552 37840 7562 37896
rect 7618 37840 7686 37896
rect 7742 37840 7810 37896
rect 7866 37840 7934 37896
rect 7990 37840 8058 37896
rect 8114 37840 8182 37896
rect 8238 37840 8306 37896
rect 8362 37840 8430 37896
rect 8486 37840 8554 37896
rect 8610 37840 8620 37896
rect 7552 37772 8620 37840
rect 7552 37716 7562 37772
rect 7618 37716 7686 37772
rect 7742 37716 7810 37772
rect 7866 37716 7934 37772
rect 7990 37716 8058 37772
rect 8114 37716 8182 37772
rect 8238 37716 8306 37772
rect 8362 37716 8430 37772
rect 8486 37716 8554 37772
rect 8610 37716 8620 37772
rect 7552 37648 8620 37716
rect 7552 37592 7562 37648
rect 7618 37592 7686 37648
rect 7742 37592 7810 37648
rect 7866 37592 7934 37648
rect 7990 37592 8058 37648
rect 8114 37592 8182 37648
rect 8238 37592 8306 37648
rect 8362 37592 8430 37648
rect 8486 37592 8554 37648
rect 8610 37592 8620 37648
rect 7552 37524 8620 37592
rect 7552 37468 7562 37524
rect 7618 37468 7686 37524
rect 7742 37468 7810 37524
rect 7866 37468 7934 37524
rect 7990 37468 8058 37524
rect 8114 37468 8182 37524
rect 8238 37468 8306 37524
rect 8362 37468 8430 37524
rect 8486 37468 8554 37524
rect 8610 37468 8620 37524
rect 7552 37400 8620 37468
rect 7552 37344 7562 37400
rect 7618 37344 7686 37400
rect 7742 37344 7810 37400
rect 7866 37344 7934 37400
rect 7990 37344 8058 37400
rect 8114 37344 8182 37400
rect 8238 37344 8306 37400
rect 8362 37344 8430 37400
rect 8486 37344 8554 37400
rect 8610 37344 8620 37400
rect 7552 37276 8620 37344
rect 7552 37220 7562 37276
rect 7618 37220 7686 37276
rect 7742 37220 7810 37276
rect 7866 37220 7934 37276
rect 7990 37220 8058 37276
rect 8114 37220 8182 37276
rect 8238 37220 8306 37276
rect 8362 37220 8430 37276
rect 8486 37220 8554 37276
rect 8610 37220 8620 37276
rect 7552 37152 8620 37220
rect 7552 37096 7562 37152
rect 7618 37096 7686 37152
rect 7742 37096 7810 37152
rect 7866 37096 7934 37152
rect 7990 37096 8058 37152
rect 8114 37096 8182 37152
rect 8238 37096 8306 37152
rect 8362 37096 8430 37152
rect 8486 37096 8554 37152
rect 8610 37096 8620 37152
rect 7552 37028 8620 37096
rect 7552 36972 7562 37028
rect 7618 36972 7686 37028
rect 7742 36972 7810 37028
rect 7866 36972 7934 37028
rect 7990 36972 8058 37028
rect 8114 36972 8182 37028
rect 8238 36972 8306 37028
rect 8362 36972 8430 37028
rect 8486 36972 8554 37028
rect 8610 36972 8620 37028
rect 7552 36904 8620 36972
rect 7552 36848 7562 36904
rect 7618 36848 7686 36904
rect 7742 36848 7810 36904
rect 7866 36848 7934 36904
rect 7990 36848 8058 36904
rect 8114 36848 8182 36904
rect 8238 36848 8306 36904
rect 8362 36848 8430 36904
rect 8486 36848 8554 36904
rect 8610 36848 8620 36904
rect 7552 36838 8620 36848
rect 10669 38144 12481 38154
rect 10669 38088 10679 38144
rect 10735 38088 10803 38144
rect 10859 38088 10927 38144
rect 10983 38088 11051 38144
rect 11107 38088 11175 38144
rect 11231 38088 11299 38144
rect 11355 38088 11423 38144
rect 11479 38088 11547 38144
rect 11603 38088 11671 38144
rect 11727 38088 11795 38144
rect 11851 38088 11919 38144
rect 11975 38088 12043 38144
rect 12099 38088 12167 38144
rect 12223 38088 12291 38144
rect 12347 38088 12415 38144
rect 12471 38088 12481 38144
rect 10669 38020 12481 38088
rect 10669 37964 10679 38020
rect 10735 37964 10803 38020
rect 10859 37964 10927 38020
rect 10983 37964 11051 38020
rect 11107 37964 11175 38020
rect 11231 37964 11299 38020
rect 11355 37964 11423 38020
rect 11479 37964 11547 38020
rect 11603 37964 11671 38020
rect 11727 37964 11795 38020
rect 11851 37964 11919 38020
rect 11975 37964 12043 38020
rect 12099 37964 12167 38020
rect 12223 37964 12291 38020
rect 12347 37964 12415 38020
rect 12471 37964 12481 38020
rect 10669 37896 12481 37964
rect 10669 37840 10679 37896
rect 10735 37840 10803 37896
rect 10859 37840 10927 37896
rect 10983 37840 11051 37896
rect 11107 37840 11175 37896
rect 11231 37840 11299 37896
rect 11355 37840 11423 37896
rect 11479 37840 11547 37896
rect 11603 37840 11671 37896
rect 11727 37840 11795 37896
rect 11851 37840 11919 37896
rect 11975 37840 12043 37896
rect 12099 37840 12167 37896
rect 12223 37840 12291 37896
rect 12347 37840 12415 37896
rect 12471 37840 12481 37896
rect 10669 37772 12481 37840
rect 10669 37716 10679 37772
rect 10735 37716 10803 37772
rect 10859 37716 10927 37772
rect 10983 37716 11051 37772
rect 11107 37716 11175 37772
rect 11231 37716 11299 37772
rect 11355 37716 11423 37772
rect 11479 37716 11547 37772
rect 11603 37716 11671 37772
rect 11727 37716 11795 37772
rect 11851 37716 11919 37772
rect 11975 37716 12043 37772
rect 12099 37716 12167 37772
rect 12223 37716 12291 37772
rect 12347 37716 12415 37772
rect 12471 37716 12481 37772
rect 10669 37648 12481 37716
rect 10669 37592 10679 37648
rect 10735 37592 10803 37648
rect 10859 37592 10927 37648
rect 10983 37592 11051 37648
rect 11107 37592 11175 37648
rect 11231 37592 11299 37648
rect 11355 37592 11423 37648
rect 11479 37592 11547 37648
rect 11603 37592 11671 37648
rect 11727 37592 11795 37648
rect 11851 37592 11919 37648
rect 11975 37592 12043 37648
rect 12099 37592 12167 37648
rect 12223 37592 12291 37648
rect 12347 37592 12415 37648
rect 12471 37592 12481 37648
rect 10669 37524 12481 37592
rect 10669 37468 10679 37524
rect 10735 37468 10803 37524
rect 10859 37468 10927 37524
rect 10983 37468 11051 37524
rect 11107 37468 11175 37524
rect 11231 37468 11299 37524
rect 11355 37468 11423 37524
rect 11479 37468 11547 37524
rect 11603 37468 11671 37524
rect 11727 37468 11795 37524
rect 11851 37468 11919 37524
rect 11975 37468 12043 37524
rect 12099 37468 12167 37524
rect 12223 37468 12291 37524
rect 12347 37468 12415 37524
rect 12471 37468 12481 37524
rect 10669 37400 12481 37468
rect 10669 37344 10679 37400
rect 10735 37344 10803 37400
rect 10859 37344 10927 37400
rect 10983 37344 11051 37400
rect 11107 37344 11175 37400
rect 11231 37344 11299 37400
rect 11355 37344 11423 37400
rect 11479 37344 11547 37400
rect 11603 37344 11671 37400
rect 11727 37344 11795 37400
rect 11851 37344 11919 37400
rect 11975 37344 12043 37400
rect 12099 37344 12167 37400
rect 12223 37344 12291 37400
rect 12347 37344 12415 37400
rect 12471 37344 12481 37400
rect 10669 37276 12481 37344
rect 10669 37220 10679 37276
rect 10735 37220 10803 37276
rect 10859 37220 10927 37276
rect 10983 37220 11051 37276
rect 11107 37220 11175 37276
rect 11231 37220 11299 37276
rect 11355 37220 11423 37276
rect 11479 37220 11547 37276
rect 11603 37220 11671 37276
rect 11727 37220 11795 37276
rect 11851 37220 11919 37276
rect 11975 37220 12043 37276
rect 12099 37220 12167 37276
rect 12223 37220 12291 37276
rect 12347 37220 12415 37276
rect 12471 37220 12481 37276
rect 10669 37152 12481 37220
rect 10669 37096 10679 37152
rect 10735 37096 10803 37152
rect 10859 37096 10927 37152
rect 10983 37096 11051 37152
rect 11107 37096 11175 37152
rect 11231 37096 11299 37152
rect 11355 37096 11423 37152
rect 11479 37096 11547 37152
rect 11603 37096 11671 37152
rect 11727 37096 11795 37152
rect 11851 37096 11919 37152
rect 11975 37096 12043 37152
rect 12099 37096 12167 37152
rect 12223 37096 12291 37152
rect 12347 37096 12415 37152
rect 12471 37096 12481 37152
rect 10669 37028 12481 37096
rect 10669 36972 10679 37028
rect 10735 36972 10803 37028
rect 10859 36972 10927 37028
rect 10983 36972 11051 37028
rect 11107 36972 11175 37028
rect 11231 36972 11299 37028
rect 11355 36972 11423 37028
rect 11479 36972 11547 37028
rect 11603 36972 11671 37028
rect 11727 36972 11795 37028
rect 11851 36972 11919 37028
rect 11975 36972 12043 37028
rect 12099 36972 12167 37028
rect 12223 36972 12291 37028
rect 12347 36972 12415 37028
rect 12471 36972 12481 37028
rect 10669 36904 12481 36972
rect 10669 36848 10679 36904
rect 10735 36848 10803 36904
rect 10859 36848 10927 36904
rect 10983 36848 11051 36904
rect 11107 36848 11175 36904
rect 11231 36848 11299 36904
rect 11355 36848 11423 36904
rect 11479 36848 11547 36904
rect 11603 36848 11671 36904
rect 11727 36848 11795 36904
rect 11851 36848 11919 36904
rect 11975 36848 12043 36904
rect 12099 36848 12167 36904
rect 12223 36848 12291 36904
rect 12347 36848 12415 36904
rect 12471 36848 12481 36904
rect 10669 36838 12481 36848
rect 4129 36725 4205 36793
rect 4129 36669 4139 36725
rect 4195 36669 4205 36725
rect 4129 36601 4205 36669
rect 4129 36545 4139 36601
rect 4195 36545 4205 36601
rect 14757 36572 14833 36582
rect 4129 36477 4205 36545
rect 4129 36421 4139 36477
rect 4195 36421 4205 36477
rect 4129 36353 4205 36421
rect 4129 36297 4139 36353
rect 4195 36297 4205 36353
rect 4129 36229 4205 36297
rect 4129 36173 4139 36229
rect 4195 36173 4205 36229
rect 4129 36105 4205 36173
rect 4129 36049 4139 36105
rect 4195 36049 4205 36105
rect 4129 35981 4205 36049
rect 4129 35925 4139 35981
rect 4195 35925 4205 35981
rect 4129 35915 4205 35925
rect 6358 36544 7426 36554
rect 6358 36488 6368 36544
rect 6424 36488 6492 36544
rect 6548 36488 6616 36544
rect 6672 36488 6740 36544
rect 6796 36488 6864 36544
rect 6920 36488 6988 36544
rect 7044 36488 7112 36544
rect 7168 36488 7236 36544
rect 7292 36488 7360 36544
rect 7416 36488 7426 36544
rect 6358 36420 7426 36488
rect 6358 36364 6368 36420
rect 6424 36364 6492 36420
rect 6548 36364 6616 36420
rect 6672 36364 6740 36420
rect 6796 36364 6864 36420
rect 6920 36364 6988 36420
rect 7044 36364 7112 36420
rect 7168 36364 7236 36420
rect 7292 36364 7360 36420
rect 7416 36364 7426 36420
rect 6358 36296 7426 36364
rect 6358 36240 6368 36296
rect 6424 36240 6492 36296
rect 6548 36240 6616 36296
rect 6672 36240 6740 36296
rect 6796 36240 6864 36296
rect 6920 36240 6988 36296
rect 7044 36240 7112 36296
rect 7168 36240 7236 36296
rect 7292 36240 7360 36296
rect 7416 36240 7426 36296
rect 6358 36172 7426 36240
rect 6358 36116 6368 36172
rect 6424 36116 6492 36172
rect 6548 36116 6616 36172
rect 6672 36116 6740 36172
rect 6796 36116 6864 36172
rect 6920 36116 6988 36172
rect 7044 36116 7112 36172
rect 7168 36116 7236 36172
rect 7292 36116 7360 36172
rect 7416 36116 7426 36172
rect 6358 36048 7426 36116
rect 6358 35992 6368 36048
rect 6424 35992 6492 36048
rect 6548 35992 6616 36048
rect 6672 35992 6740 36048
rect 6796 35992 6864 36048
rect 6920 35992 6988 36048
rect 7044 35992 7112 36048
rect 7168 35992 7236 36048
rect 7292 35992 7360 36048
rect 7416 35992 7426 36048
rect 6358 35924 7426 35992
rect 6358 35868 6368 35924
rect 6424 35868 6492 35924
rect 6548 35868 6616 35924
rect 6672 35868 6740 35924
rect 6796 35868 6864 35924
rect 6920 35868 6988 35924
rect 7044 35868 7112 35924
rect 7168 35868 7236 35924
rect 7292 35868 7360 35924
rect 7416 35868 7426 35924
rect 6358 35800 7426 35868
rect 6358 35744 6368 35800
rect 6424 35744 6492 35800
rect 6548 35744 6616 35800
rect 6672 35744 6740 35800
rect 6796 35744 6864 35800
rect 6920 35744 6988 35800
rect 7044 35744 7112 35800
rect 7168 35744 7236 35800
rect 7292 35744 7360 35800
rect 7416 35744 7426 35800
rect 6358 35676 7426 35744
rect 6358 35620 6368 35676
rect 6424 35620 6492 35676
rect 6548 35620 6616 35676
rect 6672 35620 6740 35676
rect 6796 35620 6864 35676
rect 6920 35620 6988 35676
rect 7044 35620 7112 35676
rect 7168 35620 7236 35676
rect 7292 35620 7360 35676
rect 7416 35620 7426 35676
rect 6358 35552 7426 35620
rect 6358 35496 6368 35552
rect 6424 35496 6492 35552
rect 6548 35496 6616 35552
rect 6672 35496 6740 35552
rect 6796 35496 6864 35552
rect 6920 35496 6988 35552
rect 7044 35496 7112 35552
rect 7168 35496 7236 35552
rect 7292 35496 7360 35552
rect 7416 35496 7426 35552
rect 6358 35428 7426 35496
rect 6358 35372 6368 35428
rect 6424 35372 6492 35428
rect 6548 35372 6616 35428
rect 6672 35372 6740 35428
rect 6796 35372 6864 35428
rect 6920 35372 6988 35428
rect 7044 35372 7112 35428
rect 7168 35372 7236 35428
rect 7292 35372 7360 35428
rect 7416 35372 7426 35428
rect 6358 35304 7426 35372
rect 6358 35248 6368 35304
rect 6424 35248 6492 35304
rect 6548 35248 6616 35304
rect 6672 35248 6740 35304
rect 6796 35248 6864 35304
rect 6920 35248 6988 35304
rect 7044 35248 7112 35304
rect 7168 35248 7236 35304
rect 7292 35248 7360 35304
rect 7416 35248 7426 35304
rect 6358 35238 7426 35248
rect 8741 36544 10553 36554
rect 8741 36488 8751 36544
rect 8807 36488 8875 36544
rect 8931 36488 8999 36544
rect 9055 36488 9123 36544
rect 9179 36488 9247 36544
rect 9303 36488 9371 36544
rect 9427 36488 9495 36544
rect 9551 36488 9619 36544
rect 9675 36488 9743 36544
rect 9799 36488 9867 36544
rect 9923 36488 9991 36544
rect 10047 36488 10115 36544
rect 10171 36488 10239 36544
rect 10295 36488 10363 36544
rect 10419 36488 10487 36544
rect 10543 36488 10553 36544
rect 8741 36420 10553 36488
rect 8741 36364 8751 36420
rect 8807 36364 8875 36420
rect 8931 36364 8999 36420
rect 9055 36364 9123 36420
rect 9179 36364 9247 36420
rect 9303 36364 9371 36420
rect 9427 36364 9495 36420
rect 9551 36364 9619 36420
rect 9675 36364 9743 36420
rect 9799 36364 9867 36420
rect 9923 36364 9991 36420
rect 10047 36364 10115 36420
rect 10171 36364 10239 36420
rect 10295 36364 10363 36420
rect 10419 36364 10487 36420
rect 10543 36364 10553 36420
rect 8741 36296 10553 36364
rect 8741 36240 8751 36296
rect 8807 36240 8875 36296
rect 8931 36240 8999 36296
rect 9055 36240 9123 36296
rect 9179 36240 9247 36296
rect 9303 36240 9371 36296
rect 9427 36240 9495 36296
rect 9551 36240 9619 36296
rect 9675 36240 9743 36296
rect 9799 36240 9867 36296
rect 9923 36240 9991 36296
rect 10047 36240 10115 36296
rect 10171 36240 10239 36296
rect 10295 36240 10363 36296
rect 10419 36240 10487 36296
rect 10543 36240 10553 36296
rect 8741 36172 10553 36240
rect 8741 36116 8751 36172
rect 8807 36116 8875 36172
rect 8931 36116 8999 36172
rect 9055 36116 9123 36172
rect 9179 36116 9247 36172
rect 9303 36116 9371 36172
rect 9427 36116 9495 36172
rect 9551 36116 9619 36172
rect 9675 36116 9743 36172
rect 9799 36116 9867 36172
rect 9923 36116 9991 36172
rect 10047 36116 10115 36172
rect 10171 36116 10239 36172
rect 10295 36116 10363 36172
rect 10419 36116 10487 36172
rect 10543 36116 10553 36172
rect 8741 36048 10553 36116
rect 8741 35992 8751 36048
rect 8807 35992 8875 36048
rect 8931 35992 8999 36048
rect 9055 35992 9123 36048
rect 9179 35992 9247 36048
rect 9303 35992 9371 36048
rect 9427 35992 9495 36048
rect 9551 35992 9619 36048
rect 9675 35992 9743 36048
rect 9799 35992 9867 36048
rect 9923 35992 9991 36048
rect 10047 35992 10115 36048
rect 10171 35992 10239 36048
rect 10295 35992 10363 36048
rect 10419 35992 10487 36048
rect 10543 35992 10553 36048
rect 8741 35924 10553 35992
rect 8741 35868 8751 35924
rect 8807 35868 8875 35924
rect 8931 35868 8999 35924
rect 9055 35868 9123 35924
rect 9179 35868 9247 35924
rect 9303 35868 9371 35924
rect 9427 35868 9495 35924
rect 9551 35868 9619 35924
rect 9675 35868 9743 35924
rect 9799 35868 9867 35924
rect 9923 35868 9991 35924
rect 10047 35868 10115 35924
rect 10171 35868 10239 35924
rect 10295 35868 10363 35924
rect 10419 35868 10487 35924
rect 10543 35868 10553 35924
rect 8741 35800 10553 35868
rect 8741 35744 8751 35800
rect 8807 35744 8875 35800
rect 8931 35744 8999 35800
rect 9055 35744 9123 35800
rect 9179 35744 9247 35800
rect 9303 35744 9371 35800
rect 9427 35744 9495 35800
rect 9551 35744 9619 35800
rect 9675 35744 9743 35800
rect 9799 35744 9867 35800
rect 9923 35744 9991 35800
rect 10047 35744 10115 35800
rect 10171 35744 10239 35800
rect 10295 35744 10363 35800
rect 10419 35744 10487 35800
rect 10543 35744 10553 35800
rect 8741 35676 10553 35744
rect 8741 35620 8751 35676
rect 8807 35620 8875 35676
rect 8931 35620 8999 35676
rect 9055 35620 9123 35676
rect 9179 35620 9247 35676
rect 9303 35620 9371 35676
rect 9427 35620 9495 35676
rect 9551 35620 9619 35676
rect 9675 35620 9743 35676
rect 9799 35620 9867 35676
rect 9923 35620 9991 35676
rect 10047 35620 10115 35676
rect 10171 35620 10239 35676
rect 10295 35620 10363 35676
rect 10419 35620 10487 35676
rect 10543 35620 10553 35676
rect 8741 35552 10553 35620
rect 8741 35496 8751 35552
rect 8807 35496 8875 35552
rect 8931 35496 8999 35552
rect 9055 35496 9123 35552
rect 9179 35496 9247 35552
rect 9303 35496 9371 35552
rect 9427 35496 9495 35552
rect 9551 35496 9619 35552
rect 9675 35496 9743 35552
rect 9799 35496 9867 35552
rect 9923 35496 9991 35552
rect 10047 35496 10115 35552
rect 10171 35496 10239 35552
rect 10295 35496 10363 35552
rect 10419 35496 10487 35552
rect 10543 35496 10553 35552
rect 8741 35428 10553 35496
rect 8741 35372 8751 35428
rect 8807 35372 8875 35428
rect 8931 35372 8999 35428
rect 9055 35372 9123 35428
rect 9179 35372 9247 35428
rect 9303 35372 9371 35428
rect 9427 35372 9495 35428
rect 9551 35372 9619 35428
rect 9675 35372 9743 35428
rect 9799 35372 9867 35428
rect 9923 35372 9991 35428
rect 10047 35372 10115 35428
rect 10171 35372 10239 35428
rect 10295 35372 10363 35428
rect 10419 35372 10487 35428
rect 10543 35372 10553 35428
rect 8741 35304 10553 35372
rect 8741 35248 8751 35304
rect 8807 35248 8875 35304
rect 8931 35248 8999 35304
rect 9055 35248 9123 35304
rect 9179 35248 9247 35304
rect 9303 35248 9371 35304
rect 9427 35248 9495 35304
rect 9551 35248 9619 35304
rect 9675 35248 9743 35304
rect 9799 35248 9867 35304
rect 9923 35248 9991 35304
rect 10047 35248 10115 35304
rect 10171 35248 10239 35304
rect 10295 35248 10363 35304
rect 10419 35248 10487 35304
rect 10543 35248 10553 35304
rect 8741 35238 10553 35248
rect 12842 36544 13910 36554
rect 12842 36488 12852 36544
rect 12908 36488 12976 36544
rect 13032 36488 13100 36544
rect 13156 36488 13224 36544
rect 13280 36488 13348 36544
rect 13404 36488 13472 36544
rect 13528 36488 13596 36544
rect 13652 36488 13720 36544
rect 13776 36488 13844 36544
rect 13900 36488 13910 36544
rect 12842 36420 13910 36488
rect 12842 36364 12852 36420
rect 12908 36364 12976 36420
rect 13032 36364 13100 36420
rect 13156 36364 13224 36420
rect 13280 36364 13348 36420
rect 13404 36364 13472 36420
rect 13528 36364 13596 36420
rect 13652 36364 13720 36420
rect 13776 36364 13844 36420
rect 13900 36364 13910 36420
rect 12842 36296 13910 36364
rect 12842 36240 12852 36296
rect 12908 36240 12976 36296
rect 13032 36240 13100 36296
rect 13156 36240 13224 36296
rect 13280 36240 13348 36296
rect 13404 36240 13472 36296
rect 13528 36240 13596 36296
rect 13652 36240 13720 36296
rect 13776 36240 13844 36296
rect 13900 36240 13910 36296
rect 12842 36172 13910 36240
rect 12842 36116 12852 36172
rect 12908 36116 12976 36172
rect 13032 36116 13100 36172
rect 13156 36116 13224 36172
rect 13280 36116 13348 36172
rect 13404 36116 13472 36172
rect 13528 36116 13596 36172
rect 13652 36116 13720 36172
rect 13776 36116 13844 36172
rect 13900 36116 13910 36172
rect 12842 36048 13910 36116
rect 12842 35992 12852 36048
rect 12908 35992 12976 36048
rect 13032 35992 13100 36048
rect 13156 35992 13224 36048
rect 13280 35992 13348 36048
rect 13404 35992 13472 36048
rect 13528 35992 13596 36048
rect 13652 35992 13720 36048
rect 13776 35992 13844 36048
rect 13900 35992 13910 36048
rect 12842 35924 13910 35992
rect 12842 35868 12852 35924
rect 12908 35868 12976 35924
rect 13032 35868 13100 35924
rect 13156 35868 13224 35924
rect 13280 35868 13348 35924
rect 13404 35868 13472 35924
rect 13528 35868 13596 35924
rect 13652 35868 13720 35924
rect 13776 35868 13844 35924
rect 13900 35868 13910 35924
rect 12842 35800 13910 35868
rect 12842 35744 12852 35800
rect 12908 35744 12976 35800
rect 13032 35744 13100 35800
rect 13156 35744 13224 35800
rect 13280 35744 13348 35800
rect 13404 35744 13472 35800
rect 13528 35744 13596 35800
rect 13652 35744 13720 35800
rect 13776 35744 13844 35800
rect 13900 35744 13910 35800
rect 12842 35676 13910 35744
rect 12842 35620 12852 35676
rect 12908 35620 12976 35676
rect 13032 35620 13100 35676
rect 13156 35620 13224 35676
rect 13280 35620 13348 35676
rect 13404 35620 13472 35676
rect 13528 35620 13596 35676
rect 13652 35620 13720 35676
rect 13776 35620 13844 35676
rect 13900 35620 13910 35676
rect 12842 35552 13910 35620
rect 12842 35496 12852 35552
rect 12908 35496 12976 35552
rect 13032 35496 13100 35552
rect 13156 35496 13224 35552
rect 13280 35496 13348 35552
rect 13404 35496 13472 35552
rect 13528 35496 13596 35552
rect 13652 35496 13720 35552
rect 13776 35496 13844 35552
rect 13900 35496 13910 35552
rect 12842 35428 13910 35496
rect 12842 35372 12852 35428
rect 12908 35372 12976 35428
rect 13032 35372 13100 35428
rect 13156 35372 13224 35428
rect 13280 35372 13348 35428
rect 13404 35372 13472 35428
rect 13528 35372 13596 35428
rect 13652 35372 13720 35428
rect 13776 35372 13844 35428
rect 13900 35372 13910 35428
rect 12842 35304 13910 35372
rect 12842 35248 12852 35304
rect 12908 35248 12976 35304
rect 13032 35248 13100 35304
rect 13156 35248 13224 35304
rect 13280 35248 13348 35304
rect 13404 35248 13472 35304
rect 13528 35248 13596 35304
rect 13652 35248 13720 35304
rect 13776 35248 13844 35304
rect 13900 35248 13910 35304
rect 12842 35238 13910 35248
rect 14757 35220 14767 36572
rect 14823 35220 14833 36572
rect 14757 35210 14833 35220
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_0
timestamp 1755005639
transform 1 0 14795 0 1 35896
box 0 0 1 1
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_1
timestamp 1755005639
transform 1 0 14795 0 1 50296
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_0
timestamp 1755005639
transform 1 0 14795 0 1 35896
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_1
timestamp 1755005639
transform 1 0 14795 0 1 50296
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_0
timestamp 1755005639
transform 1 0 9647 0 1 35896
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_1
timestamp 1755005639
transform 1 0 11575 0 1 48698
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_2
timestamp 1755005639
transform 1 0 11575 0 1 37496
box 0 0 1 1
use M3_M2_CDNS_40661953145777  M3_M2_CDNS_40661953145777_0
timestamp 1755005639
transform 1 0 9150 0 1 52151
box 0 0 1 1
use M3_M2_CDNS_40661953145778  M3_M2_CDNS_40661953145778_0
timestamp 1755005639
transform 1 0 8050 0 1 50990
box 0 0 1 1
use M3_M2_CDNS_40661953145779  M3_M2_CDNS_40661953145779_0
timestamp 1755005639
transform 1 0 6592 0 1 54844
box 0 0 1 1
use M3_M2_CDNS_40661953145780  M3_M2_CDNS_40661953145780_0
timestamp 1755005639
transform 1 0 8050 0 1 54607
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_0
timestamp 1755005639
transform 1 0 13376 0 1 35896
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_1
timestamp 1755005639
transform 1 0 13376 0 1 50290
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_2
timestamp 1755005639
transform 1 0 8086 0 1 37496
box 0 0 1 1
use M3_M2_CDNS_40661953145781  M3_M2_CDNS_40661953145781_3
timestamp 1755005639
transform 1 0 6892 0 1 35896
box 0 0 1 1
use M3_M2_CDNS_40661953145782  M3_M2_CDNS_40661953145782_0
timestamp 1755005639
transform 1 0 1132 0 1 42056
box 0 0 1 1
use M3_M2_CDNS_40661953145782  M3_M2_CDNS_40661953145782_1
timestamp 1755005639
transform 1 0 4498 0 1 38690
box 0 0 1 1
use M3_M2_CDNS_40661953145782  M3_M2_CDNS_40661953145782_2
timestamp 1755005639
transform 1 0 2555 0 1 38371
box 0 0 1 1
use M3_M2_CDNS_40661953145783  M3_M2_CDNS_40661953145783_0
timestamp 1755005639
transform 1 0 5862 0 1 37514
box 0 0 1 1
use M3_M2_CDNS_40661953145783  M3_M2_CDNS_40661953145783_1
timestamp 1755005639
transform 1 0 5986 0 1 37493
box 0 0 1 1
use M3_M2_CDNS_40661953145783  M3_M2_CDNS_40661953145783_2
timestamp 1755005639
transform 1 0 6110 0 1 37492
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_0
timestamp 1755005639
transform 1 0 3175 0 1 37751
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_1
timestamp 1755005639
transform 1 0 3299 0 1 37627
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_2
timestamp 1755005639
transform 1 0 4622 0 1 38566
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_3
timestamp 1755005639
transform 1 0 3423 0 1 37503
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_4
timestamp 1755005639
transform 1 0 4167 0 1 36759
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_5
timestamp 1755005639
transform 1 0 4746 0 1 38442
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_6
timestamp 1755005639
transform 1 0 4870 0 1 38318
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_7
timestamp 1755005639
transform 1 0 4994 0 1 38194
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_8
timestamp 1755005639
transform 1 0 5118 0 1 38070
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_9
timestamp 1755005639
transform 1 0 2679 0 1 38247
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_10
timestamp 1755005639
transform 1 0 2803 0 1 38123
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_11
timestamp 1755005639
transform 1 0 2927 0 1 37999
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_12
timestamp 1755005639
transform 1 0 3051 0 1 37875
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_13
timestamp 1755005639
transform 1 0 3547 0 1 37379
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_14
timestamp 1755005639
transform 1 0 4043 0 1 36883
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_15
timestamp 1755005639
transform 1 0 5490 0 1 37698
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_16
timestamp 1755005639
transform 1 0 5366 0 1 37822
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_17
timestamp 1755005639
transform 1 0 5242 0 1 37946
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_18
timestamp 1755005639
transform 1 0 1256 0 1 41932
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_19
timestamp 1755005639
transform 1 0 1380 0 1 41808
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_20
timestamp 1755005639
transform 1 0 1504 0 1 41684
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_21
timestamp 1755005639
transform 1 0 1628 0 1 41560
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_22
timestamp 1755005639
transform 1 0 1752 0 1 41436
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_23
timestamp 1755005639
transform 1 0 1876 0 1 41312
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_24
timestamp 1755005639
transform 1 0 2000 0 1 41188
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_25
timestamp 1755005639
transform 1 0 3671 0 1 37255
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_26
timestamp 1755005639
transform 1 0 3795 0 1 37131
box 0 0 1 1
use M3_M2_CDNS_40661953145784  M3_M2_CDNS_40661953145784_27
timestamp 1755005639
transform 1 0 3919 0 1 37007
box 0 0 1 1
use M3_M2_CDNS_40661953145785  M3_M2_CDNS_40661953145785_0
timestamp 1755005639
transform 1 0 5614 0 1 37630
box 0 0 1 1
use M3_M2_CDNS_40661953145786  M3_M2_CDNS_40661953145786_0
timestamp 1755005639
transform 1 0 5738 0 1 37563
box 0 0 1 1
<< properties >>
string GDS_END 6823174
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 6820442
<< end >>
